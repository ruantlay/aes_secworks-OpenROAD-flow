module aes (clk,
    cs,
    reset_n,
    we,
    address,
    read_data,
    write_data);
 input clk;
 input cs;
 input reset_n;
 input we;
 input [7:0] address;
 output [31:0] read_data;
 input [31:0] write_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire _19089_;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire _19096_;
 wire _19097_;
 wire _19098_;
 wire _19099_;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire _19106_;
 wire _19107_;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire _19112_;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire _19135_;
 wire _19136_;
 wire _19137_;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire _19141_;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire _19168_;
 wire _19169_;
 wire _19170_;
 wire _19171_;
 wire _19172_;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire _19179_;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire _19194_;
 wire _19195_;
 wire _19196_;
 wire _19197_;
 wire _19198_;
 wire _19199_;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire _19216_;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire _19228_;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire _19235_;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire _19241_;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire _19260_;
 wire _19261_;
 wire _19262_;
 wire _19263_;
 wire _19264_;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire _19268_;
 wire _19269_;
 wire _19270_;
 wire _19271_;
 wire _19272_;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire _19395_;
 wire _19396_;
 wire _19397_;
 wire _19398_;
 wire _19399_;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire _19407_;
 wire _19408_;
 wire _19409_;
 wire _19410_;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire _19424_;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire _19461_;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire _19472_;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire _19506_;
 wire _19507_;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire _19512_;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire _19519_;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire _19524_;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire _19530_;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire _19534_;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire _19545_;
 wire _19546_;
 wire _19547_;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire _19557_;
 wire _19558_;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire _19583_;
 wire _19584_;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire _19590_;
 wire _19591_;
 wire _19592_;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire _19605_;
 wire _19606_;
 wire _19607_;
 wire _19608_;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire _19624_;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire _19631_;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire _19635_;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire _19642_;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire _19648_;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire _19653_;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire _19671_;
 wire _19672_;
 wire _19673_;
 wire _19674_;
 wire _19675_;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire _19683_;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire _19692_;
 wire _19693_;
 wire _19694_;
 wire _19695_;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire _19719_;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire _19797_;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire _19839_;
 wire _19840_;
 wire _19841_;
 wire _19842_;
 wire _19843_;
 wire _19844_;
 wire _19845_;
 wire _19846_;
 wire _19847_;
 wire _19848_;
 wire _19849_;
 wire _19850_;
 wire _19851_;
 wire _19852_;
 wire _19853_;
 wire _19854_;
 wire _19855_;
 wire _19856_;
 wire _19857_;
 wire _19858_;
 wire _19859_;
 wire _19860_;
 wire _19861_;
 wire _19862_;
 wire _19863_;
 wire _19864_;
 wire _19865_;
 wire _19866_;
 wire _19867_;
 wire _19868_;
 wire _19869_;
 wire _19870_;
 wire _19871_;
 wire _19872_;
 wire _19873_;
 wire _19874_;
 wire _19875_;
 wire _19876_;
 wire _19877_;
 wire _19878_;
 wire _19879_;
 wire _19880_;
 wire _19881_;
 wire _19882_;
 wire _19883_;
 wire _19884_;
 wire _19885_;
 wire _19886_;
 wire _19887_;
 wire _19888_;
 wire _19889_;
 wire _19890_;
 wire _19891_;
 wire _19892_;
 wire _19893_;
 wire _19894_;
 wire _19895_;
 wire _19896_;
 wire _19897_;
 wire _19898_;
 wire _19899_;
 wire _19900_;
 wire _19901_;
 wire _19902_;
 wire _19903_;
 wire _19904_;
 wire _19905_;
 wire _19906_;
 wire _19907_;
 wire _19908_;
 wire _19909_;
 wire _19910_;
 wire _19911_;
 wire _19912_;
 wire _19913_;
 wire _19914_;
 wire _19915_;
 wire _19916_;
 wire _19917_;
 wire _19918_;
 wire _19919_;
 wire _19920_;
 wire _19921_;
 wire _19922_;
 wire _19923_;
 wire _19924_;
 wire _19925_;
 wire _19926_;
 wire _19927_;
 wire _19928_;
 wire _19929_;
 wire _19930_;
 wire _19931_;
 wire _19932_;
 wire _19933_;
 wire _19934_;
 wire _19935_;
 wire _19936_;
 wire _19937_;
 wire _19938_;
 wire _19939_;
 wire _19940_;
 wire _19941_;
 wire _19942_;
 wire _19943_;
 wire _19944_;
 wire _19945_;
 wire _19946_;
 wire _19947_;
 wire _19948_;
 wire _19949_;
 wire _19950_;
 wire _19951_;
 wire _19952_;
 wire _19953_;
 wire _19954_;
 wire _19955_;
 wire _19956_;
 wire _19957_;
 wire _19958_;
 wire _19959_;
 wire _19960_;
 wire _19961_;
 wire _19962_;
 wire _19963_;
 wire _19964_;
 wire _19965_;
 wire _19966_;
 wire _19967_;
 wire _19968_;
 wire _19969_;
 wire _19970_;
 wire _19971_;
 wire _19972_;
 wire _19973_;
 wire _19974_;
 wire _19975_;
 wire _19976_;
 wire _19977_;
 wire _19978_;
 wire _19979_;
 wire _19980_;
 wire _19981_;
 wire _19982_;
 wire _19983_;
 wire _19984_;
 wire _19985_;
 wire _19986_;
 wire _19987_;
 wire _19988_;
 wire _19989_;
 wire _19990_;
 wire _19991_;
 wire _19992_;
 wire _19993_;
 wire _19994_;
 wire _19995_;
 wire _19996_;
 wire _19997_;
 wire _19998_;
 wire _19999_;
 wire _20000_;
 wire _20001_;
 wire _20002_;
 wire _20003_;
 wire _20004_;
 wire _20005_;
 wire _20006_;
 wire _20007_;
 wire _20008_;
 wire _20009_;
 wire _20010_;
 wire _20011_;
 wire _20012_;
 wire _20013_;
 wire _20014_;
 wire _20015_;
 wire _20016_;
 wire _20017_;
 wire _20018_;
 wire _20019_;
 wire _20020_;
 wire _20021_;
 wire _20022_;
 wire _20023_;
 wire _20024_;
 wire _20025_;
 wire _20026_;
 wire _20027_;
 wire _20028_;
 wire _20029_;
 wire _20030_;
 wire _20031_;
 wire _20032_;
 wire _20033_;
 wire _20034_;
 wire _20035_;
 wire _20036_;
 wire _20037_;
 wire _20038_;
 wire _20039_;
 wire _20040_;
 wire _20041_;
 wire _20042_;
 wire _20043_;
 wire _20044_;
 wire _20045_;
 wire _20046_;
 wire _20047_;
 wire _20048_;
 wire _20049_;
 wire _20050_;
 wire _20051_;
 wire _20052_;
 wire _20053_;
 wire _20054_;
 wire _20055_;
 wire _20056_;
 wire _20057_;
 wire _20058_;
 wire _20059_;
 wire _20060_;
 wire _20061_;
 wire _20062_;
 wire _20063_;
 wire _20064_;
 wire _20065_;
 wire _20066_;
 wire _20067_;
 wire _20068_;
 wire _20069_;
 wire _20070_;
 wire _20071_;
 wire _20072_;
 wire _20073_;
 wire _20074_;
 wire _20075_;
 wire _20076_;
 wire _20077_;
 wire _20078_;
 wire _20079_;
 wire _20080_;
 wire _20081_;
 wire _20082_;
 wire _20083_;
 wire _20084_;
 wire _20085_;
 wire _20086_;
 wire _20087_;
 wire _20088_;
 wire _20089_;
 wire _20090_;
 wire _20091_;
 wire _20092_;
 wire _20093_;
 wire _20094_;
 wire _20095_;
 wire _20096_;
 wire _20097_;
 wire _20098_;
 wire _20099_;
 wire _20100_;
 wire _20101_;
 wire _20102_;
 wire _20103_;
 wire _20104_;
 wire _20105_;
 wire _20106_;
 wire _20107_;
 wire _20108_;
 wire _20109_;
 wire _20110_;
 wire _20111_;
 wire _20112_;
 wire _20113_;
 wire _20114_;
 wire _20115_;
 wire _20116_;
 wire _20117_;
 wire _20118_;
 wire _20119_;
 wire _20120_;
 wire _20121_;
 wire _20122_;
 wire _20123_;
 wire _20124_;
 wire _20125_;
 wire _20126_;
 wire _20127_;
 wire _20128_;
 wire _20129_;
 wire _20130_;
 wire _20131_;
 wire _20132_;
 wire _20133_;
 wire _20134_;
 wire _20135_;
 wire _20136_;
 wire _20137_;
 wire _20138_;
 wire _20139_;
 wire _20140_;
 wire _20141_;
 wire _20142_;
 wire _20143_;
 wire _20144_;
 wire _20145_;
 wire _20146_;
 wire _20147_;
 wire _20148_;
 wire _20149_;
 wire _20150_;
 wire _20151_;
 wire _20152_;
 wire _20153_;
 wire _20154_;
 wire _20155_;
 wire _20156_;
 wire _20157_;
 wire _20158_;
 wire _20159_;
 wire _20160_;
 wire _20161_;
 wire _20162_;
 wire _20163_;
 wire _20164_;
 wire _20165_;
 wire _20166_;
 wire _20167_;
 wire _20168_;
 wire _20169_;
 wire _20170_;
 wire _20171_;
 wire _20172_;
 wire _20173_;
 wire _20174_;
 wire _20175_;
 wire _20176_;
 wire _20177_;
 wire _20178_;
 wire _20179_;
 wire _20180_;
 wire _20181_;
 wire _20182_;
 wire _20183_;
 wire _20184_;
 wire _20185_;
 wire _20186_;
 wire _20187_;
 wire _20188_;
 wire _20189_;
 wire _20190_;
 wire _20191_;
 wire _20192_;
 wire _20193_;
 wire _20194_;
 wire _20195_;
 wire _20196_;
 wire _20197_;
 wire _20198_;
 wire _20199_;
 wire _20200_;
 wire _20201_;
 wire _20202_;
 wire _20203_;
 wire _20204_;
 wire _20205_;
 wire _20206_;
 wire _20207_;
 wire _20208_;
 wire _20209_;
 wire _20210_;
 wire _20211_;
 wire _20212_;
 wire _20213_;
 wire _20214_;
 wire _20215_;
 wire _20216_;
 wire _20217_;
 wire _20218_;
 wire _20219_;
 wire _20220_;
 wire _20221_;
 wire _20222_;
 wire _20223_;
 wire _20224_;
 wire _20225_;
 wire _20226_;
 wire _20227_;
 wire _20228_;
 wire _20229_;
 wire _20230_;
 wire _20231_;
 wire _20232_;
 wire _20233_;
 wire _20234_;
 wire _20235_;
 wire _20236_;
 wire _20237_;
 wire _20238_;
 wire _20239_;
 wire _20240_;
 wire _20241_;
 wire _20242_;
 wire _20243_;
 wire _20244_;
 wire _20245_;
 wire _20246_;
 wire _20247_;
 wire _20248_;
 wire _20249_;
 wire _20250_;
 wire _20251_;
 wire _20252_;
 wire _20253_;
 wire _20254_;
 wire _20255_;
 wire _20256_;
 wire _20257_;
 wire _20258_;
 wire _20259_;
 wire _20260_;
 wire _20261_;
 wire _20262_;
 wire _20263_;
 wire _20264_;
 wire _20265_;
 wire _20266_;
 wire _20267_;
 wire _20268_;
 wire _20269_;
 wire _20270_;
 wire _20271_;
 wire _20272_;
 wire _20273_;
 wire _20274_;
 wire _20275_;
 wire _20276_;
 wire _20277_;
 wire _20278_;
 wire _20279_;
 wire _20280_;
 wire _20281_;
 wire _20282_;
 wire _20283_;
 wire _20284_;
 wire _20285_;
 wire _20286_;
 wire _20287_;
 wire _20288_;
 wire _20289_;
 wire _20290_;
 wire _20291_;
 wire _20292_;
 wire _20293_;
 wire _20294_;
 wire _20295_;
 wire _20296_;
 wire _20297_;
 wire _20298_;
 wire _20299_;
 wire _20300_;
 wire _20301_;
 wire _20302_;
 wire _20303_;
 wire _20304_;
 wire _20305_;
 wire _20306_;
 wire _20307_;
 wire _20308_;
 wire _20309_;
 wire _20310_;
 wire _20311_;
 wire _20312_;
 wire _20313_;
 wire _20314_;
 wire _20315_;
 wire _20316_;
 wire _20317_;
 wire _20318_;
 wire _20319_;
 wire _20320_;
 wire _20321_;
 wire _20322_;
 wire _20323_;
 wire _20324_;
 wire _20325_;
 wire _20326_;
 wire _20327_;
 wire _20328_;
 wire _20329_;
 wire _20330_;
 wire _20331_;
 wire _20332_;
 wire _20333_;
 wire _20334_;
 wire _20335_;
 wire _20336_;
 wire _20337_;
 wire _20338_;
 wire _20339_;
 wire _20340_;
 wire _20341_;
 wire _20342_;
 wire _20343_;
 wire _20344_;
 wire _20345_;
 wire _20346_;
 wire _20347_;
 wire _20348_;
 wire _20349_;
 wire _20350_;
 wire _20351_;
 wire _20352_;
 wire _20353_;
 wire _20354_;
 wire _20355_;
 wire _20356_;
 wire _20357_;
 wire _20358_;
 wire _20359_;
 wire _20360_;
 wire _20361_;
 wire _20362_;
 wire _20363_;
 wire _20364_;
 wire _20365_;
 wire _20366_;
 wire _20367_;
 wire _20368_;
 wire _20369_;
 wire _20370_;
 wire _20371_;
 wire _20372_;
 wire _20373_;
 wire _20374_;
 wire _20375_;
 wire _20376_;
 wire _20377_;
 wire _20378_;
 wire _20379_;
 wire _20380_;
 wire _20381_;
 wire _20382_;
 wire _20383_;
 wire _20384_;
 wire _20385_;
 wire _20386_;
 wire _20387_;
 wire _20388_;
 wire _20389_;
 wire _20390_;
 wire _20391_;
 wire _20392_;
 wire _20393_;
 wire _20394_;
 wire _20395_;
 wire _20396_;
 wire _20397_;
 wire _20398_;
 wire _20399_;
 wire _20400_;
 wire _20401_;
 wire _20402_;
 wire _20403_;
 wire _20404_;
 wire _20405_;
 wire _20406_;
 wire _20407_;
 wire _20408_;
 wire _20409_;
 wire _20410_;
 wire _20411_;
 wire _20412_;
 wire _20413_;
 wire _20414_;
 wire _20415_;
 wire _20416_;
 wire _20417_;
 wire _20418_;
 wire _20419_;
 wire _20420_;
 wire _20421_;
 wire _20422_;
 wire _20423_;
 wire _20424_;
 wire _20425_;
 wire _20426_;
 wire _20427_;
 wire _20428_;
 wire _20429_;
 wire _20430_;
 wire _20431_;
 wire _20432_;
 wire _20433_;
 wire _20434_;
 wire _20435_;
 wire _20436_;
 wire _20437_;
 wire _20438_;
 wire _20439_;
 wire _20440_;
 wire _20441_;
 wire _20442_;
 wire _20443_;
 wire _20444_;
 wire _20445_;
 wire _20446_;
 wire _20447_;
 wire _20448_;
 wire _20449_;
 wire _20450_;
 wire _20451_;
 wire _20452_;
 wire _20453_;
 wire _20454_;
 wire _20455_;
 wire _20456_;
 wire _20457_;
 wire _20458_;
 wire _20459_;
 wire _20460_;
 wire _20461_;
 wire _20462_;
 wire _20463_;
 wire _20464_;
 wire _20465_;
 wire _20466_;
 wire _20467_;
 wire _20468_;
 wire _20469_;
 wire _20470_;
 wire _20471_;
 wire _20472_;
 wire _20473_;
 wire _20474_;
 wire _20475_;
 wire _20476_;
 wire _20477_;
 wire _20478_;
 wire _20479_;
 wire _20480_;
 wire _20481_;
 wire _20482_;
 wire _20483_;
 wire _20484_;
 wire _20485_;
 wire _20486_;
 wire _20487_;
 wire _20488_;
 wire _20489_;
 wire _20490_;
 wire _20491_;
 wire _20492_;
 wire _20493_;
 wire _20494_;
 wire _20495_;
 wire _20496_;
 wire _20497_;
 wire _20498_;
 wire _20499_;
 wire _20500_;
 wire _20501_;
 wire _20502_;
 wire _20503_;
 wire _20504_;
 wire _20505_;
 wire _20506_;
 wire _20507_;
 wire _20508_;
 wire _20509_;
 wire _20510_;
 wire _20511_;
 wire _20512_;
 wire _20513_;
 wire _20514_;
 wire _20515_;
 wire _20516_;
 wire _20517_;
 wire _20518_;
 wire _20519_;
 wire _20520_;
 wire _20521_;
 wire _20522_;
 wire _20523_;
 wire _20524_;
 wire _20525_;
 wire _20526_;
 wire _20527_;
 wire _20528_;
 wire _20529_;
 wire _20530_;
 wire _20531_;
 wire _20532_;
 wire _20533_;
 wire _20534_;
 wire _20535_;
 wire _20536_;
 wire _20537_;
 wire _20538_;
 wire _20539_;
 wire _20540_;
 wire _20541_;
 wire _20542_;
 wire _20543_;
 wire _20544_;
 wire _20545_;
 wire _20546_;
 wire _20547_;
 wire _20548_;
 wire _20549_;
 wire _20550_;
 wire _20551_;
 wire _20552_;
 wire _20553_;
 wire _20554_;
 wire _20555_;
 wire _20556_;
 wire _20557_;
 wire _20558_;
 wire _20559_;
 wire _20560_;
 wire _20561_;
 wire _20562_;
 wire _20563_;
 wire _20564_;
 wire _20565_;
 wire _20566_;
 wire _20567_;
 wire _20568_;
 wire _20569_;
 wire _20570_;
 wire _20571_;
 wire _20572_;
 wire _20573_;
 wire _20574_;
 wire _20575_;
 wire _20576_;
 wire _20577_;
 wire _20578_;
 wire _20579_;
 wire _20580_;
 wire _20581_;
 wire _20582_;
 wire _20583_;
 wire _20584_;
 wire _20585_;
 wire _20586_;
 wire _20587_;
 wire _20588_;
 wire _20589_;
 wire _20590_;
 wire _20591_;
 wire _20592_;
 wire _20593_;
 wire _20594_;
 wire _20595_;
 wire _20596_;
 wire _20597_;
 wire _20598_;
 wire _20599_;
 wire _20600_;
 wire _20601_;
 wire _20602_;
 wire _20603_;
 wire _20604_;
 wire _20605_;
 wire _20606_;
 wire _20607_;
 wire _20608_;
 wire _20609_;
 wire _20610_;
 wire _20611_;
 wire _20612_;
 wire _20613_;
 wire _20614_;
 wire _20615_;
 wire _20616_;
 wire _20617_;
 wire _20618_;
 wire _20619_;
 wire _20620_;
 wire _20621_;
 wire _20622_;
 wire _20623_;
 wire _20624_;
 wire _20625_;
 wire _20626_;
 wire _20627_;
 wire _20628_;
 wire _20629_;
 wire _20630_;
 wire _20631_;
 wire _20632_;
 wire _20633_;
 wire _20634_;
 wire _20635_;
 wire _20636_;
 wire _20637_;
 wire _20638_;
 wire _20639_;
 wire _20640_;
 wire _20641_;
 wire _20642_;
 wire _20643_;
 wire _20644_;
 wire _20645_;
 wire _20646_;
 wire _20647_;
 wire _20648_;
 wire _20649_;
 wire _20650_;
 wire _20651_;
 wire _20652_;
 wire _20653_;
 wire _20654_;
 wire _20655_;
 wire _20656_;
 wire _20657_;
 wire _20658_;
 wire _20659_;
 wire _20660_;
 wire _20661_;
 wire _20662_;
 wire _20663_;
 wire _20664_;
 wire _20665_;
 wire _20666_;
 wire _20667_;
 wire _20668_;
 wire _20669_;
 wire _20670_;
 wire _20671_;
 wire _20672_;
 wire _20673_;
 wire _20674_;
 wire _20675_;
 wire _20676_;
 wire _20677_;
 wire _20678_;
 wire _20679_;
 wire _20680_;
 wire _20681_;
 wire _20682_;
 wire _20683_;
 wire _20684_;
 wire _20685_;
 wire _20686_;
 wire _20687_;
 wire _20688_;
 wire _20689_;
 wire _20690_;
 wire _20691_;
 wire _20692_;
 wire _20693_;
 wire _20694_;
 wire _20695_;
 wire _20696_;
 wire _20697_;
 wire _20698_;
 wire _20699_;
 wire _20700_;
 wire _20701_;
 wire _20702_;
 wire _20703_;
 wire _20704_;
 wire _20705_;
 wire _20706_;
 wire _20707_;
 wire _20708_;
 wire _20709_;
 wire _20710_;
 wire _20711_;
 wire _20712_;
 wire _20713_;
 wire _20714_;
 wire _20715_;
 wire _20716_;
 wire _20717_;
 wire _20718_;
 wire _20719_;
 wire _20720_;
 wire _20721_;
 wire _20722_;
 wire _20723_;
 wire _20724_;
 wire _20725_;
 wire _20726_;
 wire _20727_;
 wire _20728_;
 wire _20729_;
 wire _20730_;
 wire _20731_;
 wire _20732_;
 wire _20733_;
 wire _20734_;
 wire _20735_;
 wire _20736_;
 wire _20737_;
 wire _20738_;
 wire _20739_;
 wire _20740_;
 wire _20741_;
 wire _20742_;
 wire _20743_;
 wire _20744_;
 wire _20745_;
 wire _20746_;
 wire _20747_;
 wire _20748_;
 wire _20749_;
 wire _20750_;
 wire _20751_;
 wire _20752_;
 wire _20753_;
 wire _20754_;
 wire _20755_;
 wire _20756_;
 wire _20757_;
 wire _20758_;
 wire _20759_;
 wire _20760_;
 wire _20761_;
 wire _20762_;
 wire _20763_;
 wire _20764_;
 wire _20765_;
 wire _20766_;
 wire _20767_;
 wire _20768_;
 wire _20769_;
 wire _20770_;
 wire _20771_;
 wire _20772_;
 wire _20773_;
 wire _20774_;
 wire _20775_;
 wire _20776_;
 wire _20777_;
 wire _20778_;
 wire _20779_;
 wire _20780_;
 wire _20781_;
 wire _20782_;
 wire _20783_;
 wire _20784_;
 wire _20785_;
 wire _20786_;
 wire _20787_;
 wire _20788_;
 wire _20789_;
 wire _20790_;
 wire _20791_;
 wire _20792_;
 wire _20793_;
 wire _20794_;
 wire _20795_;
 wire _20796_;
 wire _20797_;
 wire _20798_;
 wire _20799_;
 wire _20800_;
 wire _20801_;
 wire _20802_;
 wire _20803_;
 wire _20804_;
 wire _20805_;
 wire _20806_;
 wire _20807_;
 wire _20808_;
 wire _20809_;
 wire _20810_;
 wire _20811_;
 wire _20812_;
 wire _20813_;
 wire _20814_;
 wire _20815_;
 wire _20816_;
 wire _20817_;
 wire _20818_;
 wire _20819_;
 wire _20820_;
 wire _20821_;
 wire _20822_;
 wire _20823_;
 wire _20824_;
 wire _20825_;
 wire _20826_;
 wire _20827_;
 wire _20828_;
 wire _20829_;
 wire _20830_;
 wire _20831_;
 wire _20832_;
 wire _20833_;
 wire _20834_;
 wire _20835_;
 wire _20836_;
 wire _20837_;
 wire _20838_;
 wire _20839_;
 wire _20840_;
 wire _20841_;
 wire _20842_;
 wire _20843_;
 wire _20844_;
 wire _20845_;
 wire _20846_;
 wire _20847_;
 wire _20848_;
 wire _20849_;
 wire _20850_;
 wire _20851_;
 wire _20852_;
 wire _20853_;
 wire _20854_;
 wire _20855_;
 wire _20856_;
 wire _20857_;
 wire _20858_;
 wire _20859_;
 wire _20860_;
 wire _20861_;
 wire _20862_;
 wire _20863_;
 wire _20864_;
 wire _20865_;
 wire _20866_;
 wire _20867_;
 wire _20868_;
 wire _20869_;
 wire _20870_;
 wire _20871_;
 wire _20872_;
 wire _20873_;
 wire _20874_;
 wire _20875_;
 wire _20876_;
 wire _20877_;
 wire _20878_;
 wire _20879_;
 wire _20880_;
 wire _20881_;
 wire _20882_;
 wire _20883_;
 wire _20884_;
 wire _20885_;
 wire _20886_;
 wire _20887_;
 wire _20888_;
 wire _20889_;
 wire _20890_;
 wire _20891_;
 wire _20892_;
 wire _20893_;
 wire _20894_;
 wire _20895_;
 wire _20896_;
 wire _20897_;
 wire _20898_;
 wire _20899_;
 wire _20900_;
 wire _20901_;
 wire _20902_;
 wire _20903_;
 wire _20904_;
 wire _20905_;
 wire _20906_;
 wire _20907_;
 wire _20908_;
 wire _20909_;
 wire _20910_;
 wire _20911_;
 wire _20912_;
 wire _20913_;
 wire _20914_;
 wire _20915_;
 wire _20916_;
 wire _20917_;
 wire _20918_;
 wire _20919_;
 wire _20920_;
 wire _20921_;
 wire _20922_;
 wire _20923_;
 wire _20924_;
 wire _20925_;
 wire _20926_;
 wire _20927_;
 wire _20928_;
 wire _20929_;
 wire _20930_;
 wire _20931_;
 wire _20932_;
 wire _20933_;
 wire _20934_;
 wire _20935_;
 wire _20936_;
 wire _20937_;
 wire _20938_;
 wire _20939_;
 wire _20940_;
 wire _20941_;
 wire _20942_;
 wire _20943_;
 wire _20944_;
 wire _20945_;
 wire _20946_;
 wire _20947_;
 wire _20948_;
 wire _20949_;
 wire _20950_;
 wire _20951_;
 wire _20952_;
 wire _20953_;
 wire _20954_;
 wire _20955_;
 wire _20956_;
 wire _20957_;
 wire _20958_;
 wire _20959_;
 wire _20960_;
 wire _20961_;
 wire _20962_;
 wire _20963_;
 wire _20964_;
 wire _20965_;
 wire _20966_;
 wire _20967_;
 wire _20968_;
 wire _20969_;
 wire _20970_;
 wire _20971_;
 wire _20972_;
 wire _20973_;
 wire _20974_;
 wire _20975_;
 wire _20976_;
 wire _20977_;
 wire _20978_;
 wire _20979_;
 wire _20980_;
 wire _20981_;
 wire _20982_;
 wire _20983_;
 wire _20984_;
 wire _20985_;
 wire _20986_;
 wire _20987_;
 wire _20988_;
 wire _20989_;
 wire _20990_;
 wire _20991_;
 wire _20992_;
 wire _20993_;
 wire _20994_;
 wire _20995_;
 wire _20996_;
 wire _20997_;
 wire _20998_;
 wire _20999_;
 wire _21000_;
 wire _21001_;
 wire _21002_;
 wire _21003_;
 wire _21004_;
 wire _21005_;
 wire _21006_;
 wire _21007_;
 wire _21008_;
 wire _21009_;
 wire _21010_;
 wire _21011_;
 wire _21012_;
 wire _21013_;
 wire _21014_;
 wire _21015_;
 wire _21016_;
 wire _21017_;
 wire _21018_;
 wire _21019_;
 wire _21020_;
 wire _21021_;
 wire _21022_;
 wire _21023_;
 wire _21024_;
 wire _21025_;
 wire _21026_;
 wire _21027_;
 wire _21028_;
 wire _21029_;
 wire _21030_;
 wire _21031_;
 wire _21032_;
 wire _21033_;
 wire _21034_;
 wire _21035_;
 wire _21036_;
 wire _21037_;
 wire _21038_;
 wire _21039_;
 wire _21040_;
 wire _21041_;
 wire _21042_;
 wire _21043_;
 wire _21044_;
 wire _21045_;
 wire _21046_;
 wire _21047_;
 wire _21048_;
 wire _21049_;
 wire _21050_;
 wire _21051_;
 wire _21052_;
 wire _21053_;
 wire _21054_;
 wire _21055_;
 wire _21056_;
 wire _21057_;
 wire _21058_;
 wire _21059_;
 wire _21060_;
 wire _21061_;
 wire _21062_;
 wire _21063_;
 wire _21064_;
 wire _21065_;
 wire _21066_;
 wire _21067_;
 wire _21068_;
 wire _21069_;
 wire _21070_;
 wire _21071_;
 wire _21072_;
 wire _21073_;
 wire _21074_;
 wire _21075_;
 wire _21076_;
 wire _21077_;
 wire _21078_;
 wire _21079_;
 wire _21080_;
 wire _21081_;
 wire _21082_;
 wire _21083_;
 wire _21084_;
 wire _21085_;
 wire _21086_;
 wire _21087_;
 wire _21088_;
 wire _21089_;
 wire _21090_;
 wire _21091_;
 wire _21092_;
 wire _21093_;
 wire _21094_;
 wire _21095_;
 wire _21096_;
 wire _21097_;
 wire _21098_;
 wire _21099_;
 wire _21100_;
 wire _21101_;
 wire _21102_;
 wire _21103_;
 wire _21104_;
 wire _21105_;
 wire _21106_;
 wire _21107_;
 wire _21108_;
 wire _21109_;
 wire _21110_;
 wire _21111_;
 wire _21112_;
 wire _21113_;
 wire _21114_;
 wire _21115_;
 wire _21116_;
 wire _21117_;
 wire _21118_;
 wire _21119_;
 wire _21120_;
 wire _21121_;
 wire _21122_;
 wire _21123_;
 wire _21124_;
 wire _21125_;
 wire _21126_;
 wire _21127_;
 wire _21128_;
 wire _21129_;
 wire _21130_;
 wire _21131_;
 wire _21132_;
 wire _21133_;
 wire _21134_;
 wire _21135_;
 wire _21136_;
 wire _21137_;
 wire _21138_;
 wire _21139_;
 wire _21140_;
 wire _21141_;
 wire _21142_;
 wire _21143_;
 wire _21144_;
 wire _21145_;
 wire _21146_;
 wire _21147_;
 wire _21148_;
 wire _21149_;
 wire _21150_;
 wire _21151_;
 wire _21152_;
 wire _21153_;
 wire _21154_;
 wire _21155_;
 wire _21156_;
 wire _21157_;
 wire _21158_;
 wire _21159_;
 wire _21160_;
 wire _21161_;
 wire _21162_;
 wire _21163_;
 wire _21164_;
 wire _21165_;
 wire _21166_;
 wire _21167_;
 wire _21168_;
 wire _21169_;
 wire _21170_;
 wire _21171_;
 wire _21172_;
 wire _21173_;
 wire _21174_;
 wire _21175_;
 wire _21176_;
 wire _21177_;
 wire _21178_;
 wire _21179_;
 wire _21180_;
 wire _21181_;
 wire _21182_;
 wire _21183_;
 wire _21184_;
 wire _21185_;
 wire _21186_;
 wire _21187_;
 wire _21188_;
 wire _21189_;
 wire _21190_;
 wire _21191_;
 wire _21192_;
 wire _21193_;
 wire _21194_;
 wire _21195_;
 wire _21196_;
 wire _21197_;
 wire _21198_;
 wire _21199_;
 wire _21200_;
 wire _21201_;
 wire _21202_;
 wire _21203_;
 wire _21204_;
 wire _21205_;
 wire _21206_;
 wire _21207_;
 wire _21208_;
 wire _21209_;
 wire _21210_;
 wire _21211_;
 wire _21212_;
 wire _21213_;
 wire _21214_;
 wire _21215_;
 wire _21216_;
 wire _21217_;
 wire _21218_;
 wire _21219_;
 wire _21220_;
 wire _21221_;
 wire _21222_;
 wire _21223_;
 wire _21224_;
 wire _21225_;
 wire _21226_;
 wire _21227_;
 wire _21228_;
 wire _21229_;
 wire _21230_;
 wire _21231_;
 wire _21232_;
 wire _21233_;
 wire _21234_;
 wire _21235_;
 wire _21236_;
 wire _21237_;
 wire _21238_;
 wire _21239_;
 wire _21240_;
 wire _21241_;
 wire _21242_;
 wire _21243_;
 wire _21244_;
 wire _21245_;
 wire _21246_;
 wire _21247_;
 wire _21248_;
 wire _21249_;
 wire _21250_;
 wire _21251_;
 wire _21252_;
 wire _21253_;
 wire _21254_;
 wire _21255_;
 wire _21256_;
 wire _21257_;
 wire _21258_;
 wire _21259_;
 wire _21260_;
 wire _21261_;
 wire _21262_;
 wire _21263_;
 wire _21264_;
 wire _21265_;
 wire _21266_;
 wire _21267_;
 wire _21268_;
 wire _21269_;
 wire _21270_;
 wire _21271_;
 wire _21272_;
 wire _21273_;
 wire _21274_;
 wire _21275_;
 wire _21276_;
 wire _21277_;
 wire _21278_;
 wire _21279_;
 wire _21280_;
 wire _21281_;
 wire _21282_;
 wire _21283_;
 wire _21284_;
 wire _21285_;
 wire _21286_;
 wire _21287_;
 wire _21288_;
 wire _21289_;
 wire _21290_;
 wire _21291_;
 wire _21292_;
 wire _21293_;
 wire _21294_;
 wire _21295_;
 wire _21296_;
 wire _21297_;
 wire _21298_;
 wire _21299_;
 wire _21300_;
 wire _21301_;
 wire _21302_;
 wire _21303_;
 wire _21304_;
 wire _21305_;
 wire _21306_;
 wire _21307_;
 wire _21308_;
 wire _21309_;
 wire _21310_;
 wire _21311_;
 wire _21312_;
 wire _21313_;
 wire _21314_;
 wire _21315_;
 wire _21316_;
 wire _21317_;
 wire _21318_;
 wire _21319_;
 wire _21320_;
 wire _21321_;
 wire _21322_;
 wire _21323_;
 wire _21324_;
 wire _21325_;
 wire _21326_;
 wire _21327_;
 wire _21328_;
 wire _21329_;
 wire _21330_;
 wire _21331_;
 wire _21332_;
 wire _21333_;
 wire _21334_;
 wire _21335_;
 wire _21336_;
 wire _21337_;
 wire _21338_;
 wire _21339_;
 wire _21340_;
 wire _21341_;
 wire _21342_;
 wire _21343_;
 wire _21344_;
 wire _21345_;
 wire _21346_;
 wire _21347_;
 wire _21348_;
 wire _21349_;
 wire _21350_;
 wire _21351_;
 wire _21352_;
 wire _21353_;
 wire _21354_;
 wire _21355_;
 wire _21356_;
 wire _21357_;
 wire _21358_;
 wire _21359_;
 wire _21360_;
 wire _21361_;
 wire _21362_;
 wire _21363_;
 wire _21364_;
 wire _21365_;
 wire _21366_;
 wire _21367_;
 wire _21368_;
 wire _21369_;
 wire _21370_;
 wire _21371_;
 wire _21372_;
 wire _21373_;
 wire _21374_;
 wire _21375_;
 wire _21376_;
 wire _21377_;
 wire _21378_;
 wire _21379_;
 wire _21380_;
 wire _21381_;
 wire _21382_;
 wire _21383_;
 wire _21384_;
 wire _21385_;
 wire _21386_;
 wire _21387_;
 wire _21388_;
 wire _21389_;
 wire _21390_;
 wire _21391_;
 wire _21392_;
 wire _21393_;
 wire _21394_;
 wire _21395_;
 wire _21396_;
 wire _21397_;
 wire _21398_;
 wire _21399_;
 wire _21400_;
 wire _21401_;
 wire _21402_;
 wire _21403_;
 wire _21404_;
 wire _21405_;
 wire _21406_;
 wire _21407_;
 wire _21408_;
 wire _21409_;
 wire _21410_;
 wire _21411_;
 wire _21412_;
 wire _21413_;
 wire _21414_;
 wire _21415_;
 wire _21416_;
 wire _21417_;
 wire _21418_;
 wire _21419_;
 wire _21420_;
 wire _21421_;
 wire _21422_;
 wire _21423_;
 wire _21424_;
 wire _21425_;
 wire _21426_;
 wire _21427_;
 wire _21428_;
 wire _21429_;
 wire _21430_;
 wire _21431_;
 wire _21432_;
 wire _21433_;
 wire _21434_;
 wire _21435_;
 wire _21436_;
 wire _21437_;
 wire _21438_;
 wire _21439_;
 wire _21440_;
 wire _21441_;
 wire _21442_;
 wire _21443_;
 wire _21444_;
 wire _21445_;
 wire _21446_;
 wire _21447_;
 wire _21448_;
 wire _21449_;
 wire _21450_;
 wire _21451_;
 wire _21452_;
 wire _21453_;
 wire _21454_;
 wire _21455_;
 wire _21456_;
 wire _21457_;
 wire _21458_;
 wire _21459_;
 wire _21460_;
 wire _21461_;
 wire _21462_;
 wire _21463_;
 wire _21464_;
 wire _21465_;
 wire _21466_;
 wire _21467_;
 wire _21468_;
 wire _21469_;
 wire _21470_;
 wire _21471_;
 wire _21472_;
 wire _21473_;
 wire _21474_;
 wire _21475_;
 wire _21476_;
 wire _21477_;
 wire _21478_;
 wire _21479_;
 wire _21480_;
 wire _21481_;
 wire _21482_;
 wire _21483_;
 wire _21484_;
 wire _21485_;
 wire _21486_;
 wire _21487_;
 wire _21488_;
 wire _21489_;
 wire _21490_;
 wire _21491_;
 wire _21492_;
 wire _21493_;
 wire _21494_;
 wire _21495_;
 wire _21496_;
 wire _21497_;
 wire _21498_;
 wire _21499_;
 wire _21500_;
 wire _21501_;
 wire _21502_;
 wire _21503_;
 wire _21504_;
 wire _21505_;
 wire _21506_;
 wire _21507_;
 wire _21508_;
 wire _21509_;
 wire _21510_;
 wire _21511_;
 wire _21512_;
 wire _21513_;
 wire _21514_;
 wire _21515_;
 wire _21516_;
 wire _21517_;
 wire _21518_;
 wire _21519_;
 wire _21520_;
 wire _21521_;
 wire _21522_;
 wire _21523_;
 wire _21524_;
 wire _21525_;
 wire _21526_;
 wire _21527_;
 wire _21528_;
 wire _21529_;
 wire _21530_;
 wire _21531_;
 wire _21532_;
 wire _21533_;
 wire _21534_;
 wire _21535_;
 wire _21536_;
 wire _21537_;
 wire _21538_;
 wire _21539_;
 wire _21540_;
 wire _21541_;
 wire _21542_;
 wire _21543_;
 wire _21544_;
 wire _21545_;
 wire _21546_;
 wire _21547_;
 wire _21548_;
 wire _21549_;
 wire _21550_;
 wire _21551_;
 wire _21552_;
 wire _21553_;
 wire _21554_;
 wire _21555_;
 wire _21556_;
 wire _21557_;
 wire _21558_;
 wire _21559_;
 wire _21560_;
 wire _21561_;
 wire _21562_;
 wire _21563_;
 wire _21564_;
 wire _21565_;
 wire _21566_;
 wire _21567_;
 wire _21568_;
 wire _21569_;
 wire _21570_;
 wire _21571_;
 wire _21572_;
 wire _21573_;
 wire _21574_;
 wire _21575_;
 wire _21576_;
 wire _21577_;
 wire _21578_;
 wire _21579_;
 wire _21580_;
 wire _21581_;
 wire _21582_;
 wire _21583_;
 wire _21584_;
 wire _21585_;
 wire _21586_;
 wire _21587_;
 wire _21588_;
 wire _21589_;
 wire _21590_;
 wire _21591_;
 wire _21592_;
 wire _21593_;
 wire _21594_;
 wire _21595_;
 wire _21596_;
 wire _21597_;
 wire _21598_;
 wire _21599_;
 wire _21600_;
 wire _21601_;
 wire _21602_;
 wire _21603_;
 wire _21604_;
 wire _21605_;
 wire _21606_;
 wire _21607_;
 wire _21608_;
 wire _21609_;
 wire _21610_;
 wire _21611_;
 wire _21612_;
 wire _21613_;
 wire _21614_;
 wire _21615_;
 wire _21616_;
 wire _21617_;
 wire _21618_;
 wire _21619_;
 wire _21620_;
 wire _21621_;
 wire _21622_;
 wire _21623_;
 wire _21624_;
 wire _21625_;
 wire _21626_;
 wire _21627_;
 wire _21628_;
 wire _21629_;
 wire _21630_;
 wire _21631_;
 wire _21632_;
 wire _21633_;
 wire _21634_;
 wire _21635_;
 wire _21636_;
 wire _21637_;
 wire _21638_;
 wire _21639_;
 wire _21640_;
 wire _21641_;
 wire _21642_;
 wire _21643_;
 wire _21644_;
 wire _21645_;
 wire _21646_;
 wire _21647_;
 wire _21648_;
 wire _21649_;
 wire _21650_;
 wire _21651_;
 wire _21652_;
 wire _21653_;
 wire _21654_;
 wire _21655_;
 wire _21656_;
 wire _21657_;
 wire _21658_;
 wire _21659_;
 wire _21660_;
 wire _21661_;
 wire _21662_;
 wire _21663_;
 wire _21664_;
 wire _21665_;
 wire _21666_;
 wire _21667_;
 wire _21668_;
 wire _21669_;
 wire _21670_;
 wire _21671_;
 wire _21672_;
 wire _21673_;
 wire _21674_;
 wire _21675_;
 wire _21676_;
 wire _21677_;
 wire _21678_;
 wire _21679_;
 wire _21680_;
 wire _21681_;
 wire _21682_;
 wire _21683_;
 wire _21684_;
 wire _21685_;
 wire _21686_;
 wire _21687_;
 wire _21688_;
 wire _21689_;
 wire _21690_;
 wire _21691_;
 wire _21692_;
 wire _21693_;
 wire _21694_;
 wire _21695_;
 wire _21696_;
 wire _21697_;
 wire _21698_;
 wire _21699_;
 wire _21700_;
 wire _21701_;
 wire _21702_;
 wire _21703_;
 wire _21704_;
 wire _21705_;
 wire _21706_;
 wire _21707_;
 wire _21708_;
 wire _21709_;
 wire _21710_;
 wire _21711_;
 wire _21712_;
 wire _21713_;
 wire _21714_;
 wire _21715_;
 wire _21716_;
 wire _21717_;
 wire _21718_;
 wire _21719_;
 wire _21720_;
 wire _21721_;
 wire _21722_;
 wire _21723_;
 wire _21724_;
 wire _21725_;
 wire _21726_;
 wire _21727_;
 wire _21728_;
 wire _21729_;
 wire _21730_;
 wire _21731_;
 wire _21732_;
 wire _21733_;
 wire _21734_;
 wire _21735_;
 wire _21736_;
 wire _21737_;
 wire _21738_;
 wire _21739_;
 wire _21740_;
 wire _21741_;
 wire _21742_;
 wire _21743_;
 wire _21744_;
 wire _21745_;
 wire _21746_;
 wire _21747_;
 wire _21748_;
 wire _21749_;
 wire _21750_;
 wire _21751_;
 wire _21752_;
 wire _21753_;
 wire _21754_;
 wire _21755_;
 wire _21756_;
 wire _21757_;
 wire _21758_;
 wire _21759_;
 wire _21760_;
 wire _21761_;
 wire _21762_;
 wire _21763_;
 wire _21764_;
 wire _21765_;
 wire _21766_;
 wire _21767_;
 wire _21768_;
 wire _21769_;
 wire _21770_;
 wire _21771_;
 wire _21772_;
 wire _21773_;
 wire _21774_;
 wire _21775_;
 wire _21776_;
 wire _21777_;
 wire _21778_;
 wire _21779_;
 wire _21780_;
 wire _21781_;
 wire _21782_;
 wire _21783_;
 wire _21784_;
 wire _21785_;
 wire _21786_;
 wire _21787_;
 wire _21788_;
 wire _21789_;
 wire _21790_;
 wire _21791_;
 wire _21792_;
 wire _21793_;
 wire _21794_;
 wire _21795_;
 wire _21796_;
 wire _21797_;
 wire _21798_;
 wire _21799_;
 wire _21800_;
 wire _21801_;
 wire _21802_;
 wire _21803_;
 wire _21804_;
 wire _21805_;
 wire _21806_;
 wire _21807_;
 wire _21808_;
 wire _21809_;
 wire _21810_;
 wire _21811_;
 wire _21812_;
 wire _21813_;
 wire _21814_;
 wire _21815_;
 wire _21816_;
 wire _21817_;
 wire _21818_;
 wire _21819_;
 wire _21820_;
 wire _21821_;
 wire _21822_;
 wire _21823_;
 wire _21824_;
 wire _21825_;
 wire _21826_;
 wire _21827_;
 wire _21828_;
 wire _21829_;
 wire _21830_;
 wire _21831_;
 wire _21832_;
 wire _21833_;
 wire _21834_;
 wire _21835_;
 wire _21836_;
 wire _21837_;
 wire _21838_;
 wire _21839_;
 wire _21840_;
 wire _21841_;
 wire _21842_;
 wire _21843_;
 wire _21844_;
 wire _21845_;
 wire _21846_;
 wire _21847_;
 wire _21848_;
 wire _21849_;
 wire _21850_;
 wire _21851_;
 wire _21852_;
 wire _21853_;
 wire _21854_;
 wire _21855_;
 wire _21856_;
 wire _21857_;
 wire _21858_;
 wire _21859_;
 wire _21860_;
 wire _21861_;
 wire _21862_;
 wire _21863_;
 wire _21864_;
 wire _21865_;
 wire _21866_;
 wire _21867_;
 wire _21868_;
 wire _21869_;
 wire _21870_;
 wire _21871_;
 wire _21872_;
 wire _21873_;
 wire _21874_;
 wire _21875_;
 wire _21876_;
 wire _21877_;
 wire _21878_;
 wire _21879_;
 wire _21880_;
 wire _21881_;
 wire _21882_;
 wire _21883_;
 wire _21884_;
 wire _21885_;
 wire _21886_;
 wire _21887_;
 wire _21888_;
 wire _21889_;
 wire _21890_;
 wire _21891_;
 wire _21892_;
 wire _21893_;
 wire _21894_;
 wire _21895_;
 wire _21896_;
 wire _21897_;
 wire _21898_;
 wire _21899_;
 wire _21900_;
 wire _21901_;
 wire _21902_;
 wire _21903_;
 wire _21904_;
 wire _21905_;
 wire _21906_;
 wire _21907_;
 wire _21908_;
 wire _21909_;
 wire _21910_;
 wire _21911_;
 wire _21912_;
 wire _21913_;
 wire _21914_;
 wire _21915_;
 wire _21916_;
 wire _21917_;
 wire _21918_;
 wire _21919_;
 wire _21920_;
 wire _21921_;
 wire _21922_;
 wire _21923_;
 wire _21924_;
 wire _21925_;
 wire _21926_;
 wire _21927_;
 wire _21928_;
 wire _21929_;
 wire _21930_;
 wire _21931_;
 wire _21932_;
 wire _21933_;
 wire _21934_;
 wire _21935_;
 wire _21936_;
 wire _21937_;
 wire _21938_;
 wire _21939_;
 wire _21940_;
 wire _21941_;
 wire _21942_;
 wire _21943_;
 wire _21944_;
 wire _21945_;
 wire _21946_;
 wire _21947_;
 wire _21948_;
 wire _21949_;
 wire _21950_;
 wire _21951_;
 wire _21952_;
 wire _21953_;
 wire _21954_;
 wire _21955_;
 wire _21956_;
 wire _21957_;
 wire _21958_;
 wire _21959_;
 wire _21960_;
 wire _21961_;
 wire _21962_;
 wire _21963_;
 wire _21964_;
 wire _21965_;
 wire _21966_;
 wire _21967_;
 wire _21968_;
 wire _21969_;
 wire _21970_;
 wire _21971_;
 wire _21972_;
 wire _21973_;
 wire _21974_;
 wire _21975_;
 wire _21976_;
 wire _21977_;
 wire _21978_;
 wire _21979_;
 wire _21980_;
 wire _21981_;
 wire _21982_;
 wire _21983_;
 wire _21984_;
 wire _21985_;
 wire _21986_;
 wire _21987_;
 wire _21988_;
 wire _21989_;
 wire _21990_;
 wire _21991_;
 wire _21992_;
 wire _21993_;
 wire _21994_;
 wire _21995_;
 wire _21996_;
 wire _21997_;
 wire _21998_;
 wire _21999_;
 wire _22000_;
 wire _22001_;
 wire _22002_;
 wire _22003_;
 wire _22004_;
 wire _22005_;
 wire _22006_;
 wire _22007_;
 wire _22008_;
 wire _22009_;
 wire _22010_;
 wire _22011_;
 wire _22012_;
 wire _22013_;
 wire _22014_;
 wire _22015_;
 wire _22016_;
 wire _22017_;
 wire _22018_;
 wire _22019_;
 wire _22020_;
 wire _22021_;
 wire _22022_;
 wire _22023_;
 wire _22024_;
 wire _22025_;
 wire _22026_;
 wire _22027_;
 wire _22028_;
 wire _22029_;
 wire _22030_;
 wire _22031_;
 wire _22032_;
 wire _22033_;
 wire _22034_;
 wire _22035_;
 wire _22036_;
 wire _22037_;
 wire _22038_;
 wire _22039_;
 wire _22040_;
 wire _22041_;
 wire _22042_;
 wire _22043_;
 wire _22044_;
 wire _22045_;
 wire _22046_;
 wire _22047_;
 wire _22048_;
 wire _22049_;
 wire _22050_;
 wire _22051_;
 wire _22052_;
 wire _22053_;
 wire _22054_;
 wire _22055_;
 wire _22056_;
 wire _22057_;
 wire _22058_;
 wire _22059_;
 wire _22060_;
 wire _22061_;
 wire _22062_;
 wire _22063_;
 wire _22064_;
 wire _22065_;
 wire _22066_;
 wire _22067_;
 wire _22068_;
 wire _22069_;
 wire _22070_;
 wire _22071_;
 wire _22072_;
 wire _22073_;
 wire _22074_;
 wire _22075_;
 wire _22076_;
 wire _22077_;
 wire _22078_;
 wire _22079_;
 wire _22080_;
 wire _22081_;
 wire _22082_;
 wire _22083_;
 wire _22084_;
 wire _22085_;
 wire _22086_;
 wire _22087_;
 wire _22088_;
 wire _22089_;
 wire _22090_;
 wire _22091_;
 wire _22092_;
 wire _22093_;
 wire _22094_;
 wire _22095_;
 wire _22096_;
 wire _22097_;
 wire _22098_;
 wire _22099_;
 wire _22100_;
 wire _22101_;
 wire _22102_;
 wire _22103_;
 wire _22104_;
 wire _22105_;
 wire _22106_;
 wire _22107_;
 wire _22108_;
 wire _22109_;
 wire _22110_;
 wire _22111_;
 wire _22112_;
 wire _22113_;
 wire _22114_;
 wire _22115_;
 wire _22116_;
 wire _22117_;
 wire _22118_;
 wire _22119_;
 wire _22120_;
 wire _22121_;
 wire _22122_;
 wire _22123_;
 wire _22124_;
 wire _22125_;
 wire _22126_;
 wire _22127_;
 wire _22128_;
 wire _22129_;
 wire _22130_;
 wire _22131_;
 wire _22132_;
 wire _22133_;
 wire _22134_;
 wire _22135_;
 wire _22136_;
 wire _22137_;
 wire _22138_;
 wire _22139_;
 wire \block_reg[0][0] ;
 wire \block_reg[0][10] ;
 wire \block_reg[0][11] ;
 wire \block_reg[0][12] ;
 wire \block_reg[0][13] ;
 wire \block_reg[0][14] ;
 wire \block_reg[0][15] ;
 wire \block_reg[0][16] ;
 wire \block_reg[0][17] ;
 wire \block_reg[0][18] ;
 wire \block_reg[0][19] ;
 wire \block_reg[0][1] ;
 wire \block_reg[0][20] ;
 wire \block_reg[0][21] ;
 wire \block_reg[0][22] ;
 wire \block_reg[0][23] ;
 wire \block_reg[0][24] ;
 wire \block_reg[0][25] ;
 wire \block_reg[0][26] ;
 wire \block_reg[0][27] ;
 wire \block_reg[0][28] ;
 wire \block_reg[0][29] ;
 wire \block_reg[0][2] ;
 wire \block_reg[0][30] ;
 wire \block_reg[0][31] ;
 wire \block_reg[0][3] ;
 wire \block_reg[0][4] ;
 wire \block_reg[0][5] ;
 wire \block_reg[0][6] ;
 wire \block_reg[0][7] ;
 wire \block_reg[0][8] ;
 wire \block_reg[0][9] ;
 wire \block_reg[1][0] ;
 wire \block_reg[1][10] ;
 wire \block_reg[1][11] ;
 wire \block_reg[1][12] ;
 wire \block_reg[1][13] ;
 wire \block_reg[1][14] ;
 wire \block_reg[1][15] ;
 wire \block_reg[1][16] ;
 wire \block_reg[1][17] ;
 wire \block_reg[1][18] ;
 wire \block_reg[1][19] ;
 wire \block_reg[1][1] ;
 wire \block_reg[1][20] ;
 wire \block_reg[1][21] ;
 wire \block_reg[1][22] ;
 wire \block_reg[1][23] ;
 wire \block_reg[1][24] ;
 wire \block_reg[1][25] ;
 wire \block_reg[1][26] ;
 wire \block_reg[1][27] ;
 wire \block_reg[1][28] ;
 wire \block_reg[1][29] ;
 wire \block_reg[1][2] ;
 wire \block_reg[1][30] ;
 wire \block_reg[1][31] ;
 wire \block_reg[1][3] ;
 wire \block_reg[1][4] ;
 wire \block_reg[1][5] ;
 wire \block_reg[1][6] ;
 wire \block_reg[1][7] ;
 wire \block_reg[1][8] ;
 wire \block_reg[1][9] ;
 wire \block_reg[2][0] ;
 wire \block_reg[2][10] ;
 wire \block_reg[2][11] ;
 wire \block_reg[2][12] ;
 wire \block_reg[2][13] ;
 wire \block_reg[2][14] ;
 wire \block_reg[2][15] ;
 wire \block_reg[2][16] ;
 wire \block_reg[2][17] ;
 wire \block_reg[2][18] ;
 wire \block_reg[2][19] ;
 wire \block_reg[2][1] ;
 wire \block_reg[2][20] ;
 wire \block_reg[2][21] ;
 wire \block_reg[2][22] ;
 wire \block_reg[2][23] ;
 wire \block_reg[2][24] ;
 wire \block_reg[2][25] ;
 wire \block_reg[2][26] ;
 wire \block_reg[2][27] ;
 wire \block_reg[2][28] ;
 wire \block_reg[2][29] ;
 wire \block_reg[2][2] ;
 wire \block_reg[2][30] ;
 wire \block_reg[2][31] ;
 wire \block_reg[2][3] ;
 wire \block_reg[2][4] ;
 wire \block_reg[2][5] ;
 wire \block_reg[2][6] ;
 wire \block_reg[2][7] ;
 wire \block_reg[2][8] ;
 wire \block_reg[2][9] ;
 wire \block_reg[3][0] ;
 wire \block_reg[3][10] ;
 wire \block_reg[3][11] ;
 wire \block_reg[3][12] ;
 wire \block_reg[3][13] ;
 wire \block_reg[3][14] ;
 wire \block_reg[3][15] ;
 wire \block_reg[3][16] ;
 wire \block_reg[3][17] ;
 wire \block_reg[3][18] ;
 wire \block_reg[3][19] ;
 wire \block_reg[3][1] ;
 wire \block_reg[3][20] ;
 wire \block_reg[3][21] ;
 wire \block_reg[3][22] ;
 wire \block_reg[3][23] ;
 wire \block_reg[3][24] ;
 wire \block_reg[3][25] ;
 wire \block_reg[3][26] ;
 wire \block_reg[3][27] ;
 wire \block_reg[3][28] ;
 wire \block_reg[3][29] ;
 wire \block_reg[3][2] ;
 wire \block_reg[3][30] ;
 wire \block_reg[3][31] ;
 wire \block_reg[3][3] ;
 wire \block_reg[3][4] ;
 wire \block_reg[3][5] ;
 wire \block_reg[3][6] ;
 wire \block_reg[3][7] ;
 wire \block_reg[3][8] ;
 wire \block_reg[3][9] ;
 wire \core.aes_core_ctrl_reg[0] ;
 wire \core.aes_core_ctrl_reg[1] ;
 wire \core.aes_core_ctrl_reg[2] ;
 wire \core.dec_block.block_w0_reg[0] ;
 wire \core.dec_block.block_w0_reg[10] ;
 wire \core.dec_block.block_w0_reg[11] ;
 wire \core.dec_block.block_w0_reg[12] ;
 wire \core.dec_block.block_w0_reg[13] ;
 wire \core.dec_block.block_w0_reg[14] ;
 wire \core.dec_block.block_w0_reg[15] ;
 wire \core.dec_block.block_w0_reg[16] ;
 wire \core.dec_block.block_w0_reg[17] ;
 wire \core.dec_block.block_w0_reg[18] ;
 wire \core.dec_block.block_w0_reg[19] ;
 wire \core.dec_block.block_w0_reg[1] ;
 wire \core.dec_block.block_w0_reg[20] ;
 wire \core.dec_block.block_w0_reg[21] ;
 wire \core.dec_block.block_w0_reg[22] ;
 wire \core.dec_block.block_w0_reg[23] ;
 wire \core.dec_block.block_w0_reg[24] ;
 wire \core.dec_block.block_w0_reg[25] ;
 wire \core.dec_block.block_w0_reg[26] ;
 wire \core.dec_block.block_w0_reg[27] ;
 wire \core.dec_block.block_w0_reg[28] ;
 wire \core.dec_block.block_w0_reg[29] ;
 wire \core.dec_block.block_w0_reg[2] ;
 wire \core.dec_block.block_w0_reg[30] ;
 wire \core.dec_block.block_w0_reg[31] ;
 wire \core.dec_block.block_w0_reg[3] ;
 wire \core.dec_block.block_w0_reg[4] ;
 wire \core.dec_block.block_w0_reg[5] ;
 wire \core.dec_block.block_w0_reg[6] ;
 wire \core.dec_block.block_w0_reg[7] ;
 wire \core.dec_block.block_w0_reg[8] ;
 wire \core.dec_block.block_w0_reg[9] ;
 wire \core.dec_block.block_w1_reg[0] ;
 wire \core.dec_block.block_w1_reg[10] ;
 wire \core.dec_block.block_w1_reg[11] ;
 wire \core.dec_block.block_w1_reg[12] ;
 wire \core.dec_block.block_w1_reg[13] ;
 wire \core.dec_block.block_w1_reg[14] ;
 wire \core.dec_block.block_w1_reg[15] ;
 wire \core.dec_block.block_w1_reg[16] ;
 wire \core.dec_block.block_w1_reg[17] ;
 wire \core.dec_block.block_w1_reg[18] ;
 wire \core.dec_block.block_w1_reg[19] ;
 wire \core.dec_block.block_w1_reg[1] ;
 wire \core.dec_block.block_w1_reg[20] ;
 wire \core.dec_block.block_w1_reg[21] ;
 wire \core.dec_block.block_w1_reg[22] ;
 wire \core.dec_block.block_w1_reg[23] ;
 wire \core.dec_block.block_w1_reg[24] ;
 wire \core.dec_block.block_w1_reg[25] ;
 wire \core.dec_block.block_w1_reg[26] ;
 wire \core.dec_block.block_w1_reg[27] ;
 wire \core.dec_block.block_w1_reg[28] ;
 wire \core.dec_block.block_w1_reg[29] ;
 wire \core.dec_block.block_w1_reg[2] ;
 wire \core.dec_block.block_w1_reg[30] ;
 wire \core.dec_block.block_w1_reg[31] ;
 wire \core.dec_block.block_w1_reg[3] ;
 wire \core.dec_block.block_w1_reg[4] ;
 wire \core.dec_block.block_w1_reg[5] ;
 wire \core.dec_block.block_w1_reg[6] ;
 wire \core.dec_block.block_w1_reg[7] ;
 wire \core.dec_block.block_w1_reg[8] ;
 wire \core.dec_block.block_w1_reg[9] ;
 wire \core.dec_block.block_w2_reg[0] ;
 wire \core.dec_block.block_w2_reg[10] ;
 wire \core.dec_block.block_w2_reg[11] ;
 wire \core.dec_block.block_w2_reg[12] ;
 wire \core.dec_block.block_w2_reg[13] ;
 wire \core.dec_block.block_w2_reg[14] ;
 wire \core.dec_block.block_w2_reg[15] ;
 wire \core.dec_block.block_w2_reg[16] ;
 wire \core.dec_block.block_w2_reg[17] ;
 wire \core.dec_block.block_w2_reg[18] ;
 wire \core.dec_block.block_w2_reg[19] ;
 wire \core.dec_block.block_w2_reg[1] ;
 wire \core.dec_block.block_w2_reg[20] ;
 wire \core.dec_block.block_w2_reg[21] ;
 wire \core.dec_block.block_w2_reg[22] ;
 wire \core.dec_block.block_w2_reg[23] ;
 wire \core.dec_block.block_w2_reg[24] ;
 wire \core.dec_block.block_w2_reg[25] ;
 wire \core.dec_block.block_w2_reg[26] ;
 wire \core.dec_block.block_w2_reg[27] ;
 wire \core.dec_block.block_w2_reg[28] ;
 wire \core.dec_block.block_w2_reg[29] ;
 wire \core.dec_block.block_w2_reg[2] ;
 wire \core.dec_block.block_w2_reg[30] ;
 wire \core.dec_block.block_w2_reg[31] ;
 wire \core.dec_block.block_w2_reg[3] ;
 wire \core.dec_block.block_w2_reg[4] ;
 wire \core.dec_block.block_w2_reg[5] ;
 wire \core.dec_block.block_w2_reg[6] ;
 wire \core.dec_block.block_w2_reg[7] ;
 wire \core.dec_block.block_w2_reg[8] ;
 wire \core.dec_block.block_w2_reg[9] ;
 wire \core.dec_block.block_w3_reg[0] ;
 wire \core.dec_block.block_w3_reg[10] ;
 wire \core.dec_block.block_w3_reg[11] ;
 wire \core.dec_block.block_w3_reg[12] ;
 wire \core.dec_block.block_w3_reg[13] ;
 wire \core.dec_block.block_w3_reg[14] ;
 wire \core.dec_block.block_w3_reg[15] ;
 wire \core.dec_block.block_w3_reg[16] ;
 wire \core.dec_block.block_w3_reg[17] ;
 wire \core.dec_block.block_w3_reg[18] ;
 wire \core.dec_block.block_w3_reg[19] ;
 wire \core.dec_block.block_w3_reg[1] ;
 wire \core.dec_block.block_w3_reg[20] ;
 wire \core.dec_block.block_w3_reg[21] ;
 wire \core.dec_block.block_w3_reg[22] ;
 wire \core.dec_block.block_w3_reg[23] ;
 wire \core.dec_block.block_w3_reg[24] ;
 wire \core.dec_block.block_w3_reg[25] ;
 wire \core.dec_block.block_w3_reg[26] ;
 wire \core.dec_block.block_w3_reg[27] ;
 wire \core.dec_block.block_w3_reg[28] ;
 wire \core.dec_block.block_w3_reg[29] ;
 wire \core.dec_block.block_w3_reg[2] ;
 wire \core.dec_block.block_w3_reg[30] ;
 wire \core.dec_block.block_w3_reg[31] ;
 wire \core.dec_block.block_w3_reg[3] ;
 wire \core.dec_block.block_w3_reg[4] ;
 wire \core.dec_block.block_w3_reg[5] ;
 wire \core.dec_block.block_w3_reg[6] ;
 wire \core.dec_block.block_w3_reg[7] ;
 wire \core.dec_block.block_w3_reg[8] ;
 wire \core.dec_block.block_w3_reg[9] ;
 wire \core.dec_block.dec_ctrl_reg[0] ;
 wire \core.dec_block.dec_ctrl_reg[1] ;
 wire \core.dec_block.dec_ctrl_reg[2] ;
 wire \core.dec_block.dec_ctrl_reg[3] ;
 wire \core.dec_block.keylen ;
 wire \core.dec_block.ready ;
 wire \core.dec_block.round[0] ;
 wire \core.dec_block.round[1] ;
 wire \core.dec_block.round[2] ;
 wire \core.dec_block.round[3] ;
 wire \core.dec_block.sword_ctr_reg[0] ;
 wire \core.dec_block.sword_ctr_reg[1] ;
 wire \core.enc_block.block_w0_reg[0] ;
 wire \core.enc_block.block_w0_reg[10] ;
 wire \core.enc_block.block_w0_reg[11] ;
 wire \core.enc_block.block_w0_reg[12] ;
 wire \core.enc_block.block_w0_reg[13] ;
 wire \core.enc_block.block_w0_reg[14] ;
 wire \core.enc_block.block_w0_reg[15] ;
 wire \core.enc_block.block_w0_reg[16] ;
 wire \core.enc_block.block_w0_reg[17] ;
 wire \core.enc_block.block_w0_reg[18] ;
 wire \core.enc_block.block_w0_reg[19] ;
 wire \core.enc_block.block_w0_reg[1] ;
 wire \core.enc_block.block_w0_reg[20] ;
 wire \core.enc_block.block_w0_reg[21] ;
 wire \core.enc_block.block_w0_reg[22] ;
 wire \core.enc_block.block_w0_reg[23] ;
 wire \core.enc_block.block_w0_reg[24] ;
 wire \core.enc_block.block_w0_reg[25] ;
 wire \core.enc_block.block_w0_reg[26] ;
 wire \core.enc_block.block_w0_reg[27] ;
 wire \core.enc_block.block_w0_reg[28] ;
 wire \core.enc_block.block_w0_reg[29] ;
 wire \core.enc_block.block_w0_reg[2] ;
 wire \core.enc_block.block_w0_reg[30] ;
 wire \core.enc_block.block_w0_reg[31] ;
 wire \core.enc_block.block_w0_reg[3] ;
 wire \core.enc_block.block_w0_reg[4] ;
 wire \core.enc_block.block_w0_reg[5] ;
 wire \core.enc_block.block_w0_reg[6] ;
 wire \core.enc_block.block_w0_reg[7] ;
 wire \core.enc_block.block_w0_reg[8] ;
 wire \core.enc_block.block_w0_reg[9] ;
 wire \core.enc_block.block_w1_reg[0] ;
 wire \core.enc_block.block_w1_reg[10] ;
 wire \core.enc_block.block_w1_reg[11] ;
 wire \core.enc_block.block_w1_reg[12] ;
 wire \core.enc_block.block_w1_reg[13] ;
 wire \core.enc_block.block_w1_reg[14] ;
 wire \core.enc_block.block_w1_reg[15] ;
 wire \core.enc_block.block_w1_reg[16] ;
 wire \core.enc_block.block_w1_reg[17] ;
 wire \core.enc_block.block_w1_reg[18] ;
 wire \core.enc_block.block_w1_reg[19] ;
 wire \core.enc_block.block_w1_reg[1] ;
 wire \core.enc_block.block_w1_reg[20] ;
 wire \core.enc_block.block_w1_reg[21] ;
 wire \core.enc_block.block_w1_reg[22] ;
 wire \core.enc_block.block_w1_reg[23] ;
 wire \core.enc_block.block_w1_reg[24] ;
 wire \core.enc_block.block_w1_reg[25] ;
 wire \core.enc_block.block_w1_reg[26] ;
 wire \core.enc_block.block_w1_reg[27] ;
 wire \core.enc_block.block_w1_reg[28] ;
 wire \core.enc_block.block_w1_reg[29] ;
 wire \core.enc_block.block_w1_reg[2] ;
 wire \core.enc_block.block_w1_reg[30] ;
 wire \core.enc_block.block_w1_reg[31] ;
 wire \core.enc_block.block_w1_reg[3] ;
 wire \core.enc_block.block_w1_reg[4] ;
 wire \core.enc_block.block_w1_reg[5] ;
 wire \core.enc_block.block_w1_reg[6] ;
 wire \core.enc_block.block_w1_reg[7] ;
 wire \core.enc_block.block_w1_reg[8] ;
 wire \core.enc_block.block_w1_reg[9] ;
 wire \core.enc_block.block_w2_reg[0] ;
 wire \core.enc_block.block_w2_reg[10] ;
 wire \core.enc_block.block_w2_reg[11] ;
 wire \core.enc_block.block_w2_reg[12] ;
 wire \core.enc_block.block_w2_reg[13] ;
 wire \core.enc_block.block_w2_reg[14] ;
 wire \core.enc_block.block_w2_reg[15] ;
 wire \core.enc_block.block_w2_reg[16] ;
 wire \core.enc_block.block_w2_reg[17] ;
 wire \core.enc_block.block_w2_reg[18] ;
 wire \core.enc_block.block_w2_reg[19] ;
 wire \core.enc_block.block_w2_reg[1] ;
 wire \core.enc_block.block_w2_reg[20] ;
 wire \core.enc_block.block_w2_reg[21] ;
 wire \core.enc_block.block_w2_reg[22] ;
 wire \core.enc_block.block_w2_reg[23] ;
 wire \core.enc_block.block_w2_reg[24] ;
 wire \core.enc_block.block_w2_reg[25] ;
 wire \core.enc_block.block_w2_reg[26] ;
 wire \core.enc_block.block_w2_reg[27] ;
 wire \core.enc_block.block_w2_reg[28] ;
 wire \core.enc_block.block_w2_reg[29] ;
 wire \core.enc_block.block_w2_reg[2] ;
 wire \core.enc_block.block_w2_reg[30] ;
 wire \core.enc_block.block_w2_reg[31] ;
 wire \core.enc_block.block_w2_reg[3] ;
 wire \core.enc_block.block_w2_reg[4] ;
 wire \core.enc_block.block_w2_reg[5] ;
 wire \core.enc_block.block_w2_reg[6] ;
 wire \core.enc_block.block_w2_reg[7] ;
 wire \core.enc_block.block_w2_reg[8] ;
 wire \core.enc_block.block_w2_reg[9] ;
 wire \core.enc_block.block_w3_reg[0] ;
 wire \core.enc_block.block_w3_reg[10] ;
 wire \core.enc_block.block_w3_reg[11] ;
 wire \core.enc_block.block_w3_reg[12] ;
 wire \core.enc_block.block_w3_reg[13] ;
 wire \core.enc_block.block_w3_reg[14] ;
 wire \core.enc_block.block_w3_reg[15] ;
 wire \core.enc_block.block_w3_reg[16] ;
 wire \core.enc_block.block_w3_reg[17] ;
 wire \core.enc_block.block_w3_reg[18] ;
 wire \core.enc_block.block_w3_reg[19] ;
 wire \core.enc_block.block_w3_reg[1] ;
 wire \core.enc_block.block_w3_reg[20] ;
 wire \core.enc_block.block_w3_reg[21] ;
 wire \core.enc_block.block_w3_reg[22] ;
 wire \core.enc_block.block_w3_reg[23] ;
 wire \core.enc_block.block_w3_reg[24] ;
 wire \core.enc_block.block_w3_reg[25] ;
 wire \core.enc_block.block_w3_reg[26] ;
 wire \core.enc_block.block_w3_reg[27] ;
 wire \core.enc_block.block_w3_reg[28] ;
 wire \core.enc_block.block_w3_reg[29] ;
 wire \core.enc_block.block_w3_reg[2] ;
 wire \core.enc_block.block_w3_reg[30] ;
 wire \core.enc_block.block_w3_reg[31] ;
 wire \core.enc_block.block_w3_reg[3] ;
 wire \core.enc_block.block_w3_reg[4] ;
 wire \core.enc_block.block_w3_reg[5] ;
 wire \core.enc_block.block_w3_reg[6] ;
 wire \core.enc_block.block_w3_reg[7] ;
 wire \core.enc_block.block_w3_reg[8] ;
 wire \core.enc_block.block_w3_reg[9] ;
 wire \core.enc_block.enc_ctrl_reg[0] ;
 wire \core.enc_block.enc_ctrl_reg[1] ;
 wire \core.enc_block.enc_ctrl_reg[2] ;
 wire \core.enc_block.enc_ctrl_reg[3] ;
 wire \core.enc_block.ready ;
 wire \core.enc_block.round[0] ;
 wire \core.enc_block.round[1] ;
 wire \core.enc_block.round[2] ;
 wire \core.enc_block.round[3] ;
 wire \core.enc_block.sword_ctr_reg[0] ;
 wire \core.enc_block.sword_ctr_reg[1] ;
 wire \core.encdec ;
 wire \core.init ;
 wire \core.key[0] ;
 wire \core.key[100] ;
 wire \core.key[101] ;
 wire \core.key[102] ;
 wire \core.key[103] ;
 wire \core.key[104] ;
 wire \core.key[105] ;
 wire \core.key[106] ;
 wire \core.key[107] ;
 wire \core.key[108] ;
 wire \core.key[109] ;
 wire \core.key[10] ;
 wire \core.key[110] ;
 wire \core.key[111] ;
 wire \core.key[112] ;
 wire \core.key[113] ;
 wire \core.key[114] ;
 wire \core.key[115] ;
 wire \core.key[116] ;
 wire \core.key[117] ;
 wire \core.key[118] ;
 wire \core.key[119] ;
 wire \core.key[11] ;
 wire \core.key[120] ;
 wire \core.key[121] ;
 wire \core.key[122] ;
 wire \core.key[123] ;
 wire \core.key[124] ;
 wire \core.key[125] ;
 wire \core.key[126] ;
 wire \core.key[127] ;
 wire \core.key[128] ;
 wire \core.key[129] ;
 wire \core.key[12] ;
 wire \core.key[130] ;
 wire \core.key[131] ;
 wire \core.key[132] ;
 wire \core.key[133] ;
 wire \core.key[134] ;
 wire \core.key[135] ;
 wire \core.key[136] ;
 wire \core.key[137] ;
 wire \core.key[138] ;
 wire \core.key[139] ;
 wire \core.key[13] ;
 wire \core.key[140] ;
 wire \core.key[141] ;
 wire \core.key[142] ;
 wire \core.key[143] ;
 wire \core.key[144] ;
 wire \core.key[145] ;
 wire \core.key[146] ;
 wire \core.key[147] ;
 wire \core.key[148] ;
 wire \core.key[149] ;
 wire \core.key[14] ;
 wire \core.key[150] ;
 wire \core.key[151] ;
 wire \core.key[152] ;
 wire \core.key[153] ;
 wire \core.key[154] ;
 wire \core.key[155] ;
 wire \core.key[156] ;
 wire \core.key[157] ;
 wire \core.key[158] ;
 wire \core.key[159] ;
 wire \core.key[15] ;
 wire \core.key[160] ;
 wire \core.key[161] ;
 wire \core.key[162] ;
 wire \core.key[163] ;
 wire \core.key[164] ;
 wire \core.key[165] ;
 wire \core.key[166] ;
 wire \core.key[167] ;
 wire \core.key[168] ;
 wire \core.key[169] ;
 wire \core.key[16] ;
 wire \core.key[170] ;
 wire \core.key[171] ;
 wire \core.key[172] ;
 wire \core.key[173] ;
 wire \core.key[174] ;
 wire \core.key[175] ;
 wire \core.key[176] ;
 wire \core.key[177] ;
 wire \core.key[178] ;
 wire \core.key[179] ;
 wire \core.key[17] ;
 wire \core.key[180] ;
 wire \core.key[181] ;
 wire \core.key[182] ;
 wire \core.key[183] ;
 wire \core.key[184] ;
 wire \core.key[185] ;
 wire \core.key[186] ;
 wire \core.key[187] ;
 wire \core.key[188] ;
 wire \core.key[189] ;
 wire \core.key[18] ;
 wire \core.key[190] ;
 wire \core.key[191] ;
 wire \core.key[192] ;
 wire \core.key[193] ;
 wire \core.key[194] ;
 wire \core.key[195] ;
 wire \core.key[196] ;
 wire \core.key[197] ;
 wire \core.key[198] ;
 wire \core.key[199] ;
 wire \core.key[19] ;
 wire \core.key[1] ;
 wire \core.key[200] ;
 wire \core.key[201] ;
 wire \core.key[202] ;
 wire \core.key[203] ;
 wire \core.key[204] ;
 wire \core.key[205] ;
 wire \core.key[206] ;
 wire \core.key[207] ;
 wire \core.key[208] ;
 wire \core.key[209] ;
 wire \core.key[20] ;
 wire \core.key[210] ;
 wire \core.key[211] ;
 wire \core.key[212] ;
 wire \core.key[213] ;
 wire \core.key[214] ;
 wire \core.key[215] ;
 wire \core.key[216] ;
 wire \core.key[217] ;
 wire \core.key[218] ;
 wire \core.key[219] ;
 wire \core.key[21] ;
 wire \core.key[220] ;
 wire \core.key[221] ;
 wire \core.key[222] ;
 wire \core.key[223] ;
 wire \core.key[224] ;
 wire \core.key[225] ;
 wire \core.key[226] ;
 wire \core.key[227] ;
 wire \core.key[228] ;
 wire \core.key[229] ;
 wire \core.key[22] ;
 wire \core.key[230] ;
 wire \core.key[231] ;
 wire \core.key[232] ;
 wire \core.key[233] ;
 wire \core.key[234] ;
 wire \core.key[235] ;
 wire \core.key[236] ;
 wire \core.key[237] ;
 wire \core.key[238] ;
 wire \core.key[239] ;
 wire \core.key[23] ;
 wire \core.key[240] ;
 wire \core.key[241] ;
 wire \core.key[242] ;
 wire \core.key[243] ;
 wire \core.key[244] ;
 wire \core.key[245] ;
 wire \core.key[246] ;
 wire \core.key[247] ;
 wire \core.key[248] ;
 wire \core.key[249] ;
 wire \core.key[24] ;
 wire \core.key[250] ;
 wire \core.key[251] ;
 wire \core.key[252] ;
 wire \core.key[253] ;
 wire \core.key[254] ;
 wire \core.key[255] ;
 wire \core.key[25] ;
 wire \core.key[26] ;
 wire \core.key[27] ;
 wire \core.key[28] ;
 wire \core.key[29] ;
 wire \core.key[2] ;
 wire \core.key[30] ;
 wire \core.key[31] ;
 wire \core.key[32] ;
 wire \core.key[33] ;
 wire \core.key[34] ;
 wire \core.key[35] ;
 wire \core.key[36] ;
 wire \core.key[37] ;
 wire \core.key[38] ;
 wire \core.key[39] ;
 wire \core.key[3] ;
 wire \core.key[40] ;
 wire \core.key[41] ;
 wire \core.key[42] ;
 wire \core.key[43] ;
 wire \core.key[44] ;
 wire \core.key[45] ;
 wire \core.key[46] ;
 wire \core.key[47] ;
 wire \core.key[48] ;
 wire \core.key[49] ;
 wire \core.key[4] ;
 wire \core.key[50] ;
 wire \core.key[51] ;
 wire \core.key[52] ;
 wire \core.key[53] ;
 wire \core.key[54] ;
 wire \core.key[55] ;
 wire \core.key[56] ;
 wire \core.key[57] ;
 wire \core.key[58] ;
 wire \core.key[59] ;
 wire \core.key[5] ;
 wire \core.key[60] ;
 wire \core.key[61] ;
 wire \core.key[62] ;
 wire \core.key[63] ;
 wire \core.key[64] ;
 wire \core.key[65] ;
 wire \core.key[66] ;
 wire \core.key[67] ;
 wire \core.key[68] ;
 wire \core.key[69] ;
 wire \core.key[6] ;
 wire \core.key[70] ;
 wire \core.key[71] ;
 wire \core.key[72] ;
 wire \core.key[73] ;
 wire \core.key[74] ;
 wire \core.key[75] ;
 wire \core.key[76] ;
 wire \core.key[77] ;
 wire \core.key[78] ;
 wire \core.key[79] ;
 wire \core.key[7] ;
 wire \core.key[80] ;
 wire \core.key[81] ;
 wire \core.key[82] ;
 wire \core.key[83] ;
 wire \core.key[84] ;
 wire \core.key[85] ;
 wire \core.key[86] ;
 wire \core.key[87] ;
 wire \core.key[88] ;
 wire \core.key[89] ;
 wire \core.key[8] ;
 wire \core.key[90] ;
 wire \core.key[91] ;
 wire \core.key[92] ;
 wire \core.key[93] ;
 wire \core.key[94] ;
 wire \core.key[95] ;
 wire \core.key[96] ;
 wire \core.key[97] ;
 wire \core.key[98] ;
 wire \core.key[99] ;
 wire \core.key[9] ;
 wire \core.key_ready ;
 wire \core.keymem.key_mem[0][0] ;
 wire \core.keymem.key_mem[0][100] ;
 wire \core.keymem.key_mem[0][101] ;
 wire \core.keymem.key_mem[0][102] ;
 wire \core.keymem.key_mem[0][103] ;
 wire \core.keymem.key_mem[0][104] ;
 wire \core.keymem.key_mem[0][105] ;
 wire \core.keymem.key_mem[0][106] ;
 wire \core.keymem.key_mem[0][107] ;
 wire \core.keymem.key_mem[0][108] ;
 wire \core.keymem.key_mem[0][109] ;
 wire \core.keymem.key_mem[0][10] ;
 wire \core.keymem.key_mem[0][110] ;
 wire \core.keymem.key_mem[0][111] ;
 wire \core.keymem.key_mem[0][112] ;
 wire \core.keymem.key_mem[0][113] ;
 wire \core.keymem.key_mem[0][114] ;
 wire \core.keymem.key_mem[0][115] ;
 wire \core.keymem.key_mem[0][116] ;
 wire \core.keymem.key_mem[0][117] ;
 wire \core.keymem.key_mem[0][118] ;
 wire \core.keymem.key_mem[0][119] ;
 wire \core.keymem.key_mem[0][11] ;
 wire \core.keymem.key_mem[0][120] ;
 wire \core.keymem.key_mem[0][121] ;
 wire \core.keymem.key_mem[0][122] ;
 wire \core.keymem.key_mem[0][123] ;
 wire \core.keymem.key_mem[0][124] ;
 wire \core.keymem.key_mem[0][125] ;
 wire \core.keymem.key_mem[0][126] ;
 wire \core.keymem.key_mem[0][127] ;
 wire \core.keymem.key_mem[0][12] ;
 wire \core.keymem.key_mem[0][13] ;
 wire \core.keymem.key_mem[0][14] ;
 wire \core.keymem.key_mem[0][15] ;
 wire \core.keymem.key_mem[0][16] ;
 wire \core.keymem.key_mem[0][17] ;
 wire \core.keymem.key_mem[0][18] ;
 wire \core.keymem.key_mem[0][19] ;
 wire \core.keymem.key_mem[0][1] ;
 wire \core.keymem.key_mem[0][20] ;
 wire \core.keymem.key_mem[0][21] ;
 wire \core.keymem.key_mem[0][22] ;
 wire \core.keymem.key_mem[0][23] ;
 wire \core.keymem.key_mem[0][24] ;
 wire \core.keymem.key_mem[0][25] ;
 wire \core.keymem.key_mem[0][26] ;
 wire \core.keymem.key_mem[0][27] ;
 wire \core.keymem.key_mem[0][28] ;
 wire \core.keymem.key_mem[0][29] ;
 wire \core.keymem.key_mem[0][2] ;
 wire \core.keymem.key_mem[0][30] ;
 wire \core.keymem.key_mem[0][31] ;
 wire \core.keymem.key_mem[0][32] ;
 wire \core.keymem.key_mem[0][33] ;
 wire \core.keymem.key_mem[0][34] ;
 wire \core.keymem.key_mem[0][35] ;
 wire \core.keymem.key_mem[0][36] ;
 wire \core.keymem.key_mem[0][37] ;
 wire \core.keymem.key_mem[0][38] ;
 wire \core.keymem.key_mem[0][39] ;
 wire \core.keymem.key_mem[0][3] ;
 wire \core.keymem.key_mem[0][40] ;
 wire \core.keymem.key_mem[0][41] ;
 wire \core.keymem.key_mem[0][42] ;
 wire \core.keymem.key_mem[0][43] ;
 wire \core.keymem.key_mem[0][44] ;
 wire \core.keymem.key_mem[0][45] ;
 wire \core.keymem.key_mem[0][46] ;
 wire \core.keymem.key_mem[0][47] ;
 wire \core.keymem.key_mem[0][48] ;
 wire \core.keymem.key_mem[0][49] ;
 wire \core.keymem.key_mem[0][4] ;
 wire \core.keymem.key_mem[0][50] ;
 wire \core.keymem.key_mem[0][51] ;
 wire \core.keymem.key_mem[0][52] ;
 wire \core.keymem.key_mem[0][53] ;
 wire \core.keymem.key_mem[0][54] ;
 wire \core.keymem.key_mem[0][55] ;
 wire \core.keymem.key_mem[0][56] ;
 wire \core.keymem.key_mem[0][57] ;
 wire \core.keymem.key_mem[0][58] ;
 wire \core.keymem.key_mem[0][59] ;
 wire \core.keymem.key_mem[0][5] ;
 wire \core.keymem.key_mem[0][60] ;
 wire \core.keymem.key_mem[0][61] ;
 wire \core.keymem.key_mem[0][62] ;
 wire \core.keymem.key_mem[0][63] ;
 wire \core.keymem.key_mem[0][64] ;
 wire \core.keymem.key_mem[0][65] ;
 wire \core.keymem.key_mem[0][66] ;
 wire \core.keymem.key_mem[0][67] ;
 wire \core.keymem.key_mem[0][68] ;
 wire \core.keymem.key_mem[0][69] ;
 wire \core.keymem.key_mem[0][6] ;
 wire \core.keymem.key_mem[0][70] ;
 wire \core.keymem.key_mem[0][71] ;
 wire \core.keymem.key_mem[0][72] ;
 wire \core.keymem.key_mem[0][73] ;
 wire \core.keymem.key_mem[0][74] ;
 wire \core.keymem.key_mem[0][75] ;
 wire \core.keymem.key_mem[0][76] ;
 wire \core.keymem.key_mem[0][77] ;
 wire \core.keymem.key_mem[0][78] ;
 wire \core.keymem.key_mem[0][79] ;
 wire \core.keymem.key_mem[0][7] ;
 wire \core.keymem.key_mem[0][80] ;
 wire \core.keymem.key_mem[0][81] ;
 wire \core.keymem.key_mem[0][82] ;
 wire \core.keymem.key_mem[0][83] ;
 wire \core.keymem.key_mem[0][84] ;
 wire \core.keymem.key_mem[0][85] ;
 wire \core.keymem.key_mem[0][86] ;
 wire \core.keymem.key_mem[0][87] ;
 wire \core.keymem.key_mem[0][88] ;
 wire \core.keymem.key_mem[0][89] ;
 wire \core.keymem.key_mem[0][8] ;
 wire \core.keymem.key_mem[0][90] ;
 wire \core.keymem.key_mem[0][91] ;
 wire \core.keymem.key_mem[0][92] ;
 wire \core.keymem.key_mem[0][93] ;
 wire \core.keymem.key_mem[0][94] ;
 wire \core.keymem.key_mem[0][95] ;
 wire \core.keymem.key_mem[0][96] ;
 wire \core.keymem.key_mem[0][97] ;
 wire \core.keymem.key_mem[0][98] ;
 wire \core.keymem.key_mem[0][99] ;
 wire \core.keymem.key_mem[0][9] ;
 wire \core.keymem.key_mem[10][0] ;
 wire \core.keymem.key_mem[10][100] ;
 wire \core.keymem.key_mem[10][101] ;
 wire \core.keymem.key_mem[10][102] ;
 wire \core.keymem.key_mem[10][103] ;
 wire \core.keymem.key_mem[10][104] ;
 wire \core.keymem.key_mem[10][105] ;
 wire \core.keymem.key_mem[10][106] ;
 wire \core.keymem.key_mem[10][107] ;
 wire \core.keymem.key_mem[10][108] ;
 wire \core.keymem.key_mem[10][109] ;
 wire \core.keymem.key_mem[10][10] ;
 wire \core.keymem.key_mem[10][110] ;
 wire \core.keymem.key_mem[10][111] ;
 wire \core.keymem.key_mem[10][112] ;
 wire \core.keymem.key_mem[10][113] ;
 wire \core.keymem.key_mem[10][114] ;
 wire \core.keymem.key_mem[10][115] ;
 wire \core.keymem.key_mem[10][116] ;
 wire \core.keymem.key_mem[10][117] ;
 wire \core.keymem.key_mem[10][118] ;
 wire \core.keymem.key_mem[10][119] ;
 wire \core.keymem.key_mem[10][11] ;
 wire \core.keymem.key_mem[10][120] ;
 wire \core.keymem.key_mem[10][121] ;
 wire \core.keymem.key_mem[10][122] ;
 wire \core.keymem.key_mem[10][123] ;
 wire \core.keymem.key_mem[10][124] ;
 wire \core.keymem.key_mem[10][125] ;
 wire \core.keymem.key_mem[10][126] ;
 wire \core.keymem.key_mem[10][127] ;
 wire \core.keymem.key_mem[10][12] ;
 wire \core.keymem.key_mem[10][13] ;
 wire \core.keymem.key_mem[10][14] ;
 wire \core.keymem.key_mem[10][15] ;
 wire \core.keymem.key_mem[10][16] ;
 wire \core.keymem.key_mem[10][17] ;
 wire \core.keymem.key_mem[10][18] ;
 wire \core.keymem.key_mem[10][19] ;
 wire \core.keymem.key_mem[10][1] ;
 wire \core.keymem.key_mem[10][20] ;
 wire \core.keymem.key_mem[10][21] ;
 wire \core.keymem.key_mem[10][22] ;
 wire \core.keymem.key_mem[10][23] ;
 wire \core.keymem.key_mem[10][24] ;
 wire \core.keymem.key_mem[10][25] ;
 wire \core.keymem.key_mem[10][26] ;
 wire \core.keymem.key_mem[10][27] ;
 wire \core.keymem.key_mem[10][28] ;
 wire \core.keymem.key_mem[10][29] ;
 wire \core.keymem.key_mem[10][2] ;
 wire \core.keymem.key_mem[10][30] ;
 wire \core.keymem.key_mem[10][31] ;
 wire \core.keymem.key_mem[10][32] ;
 wire \core.keymem.key_mem[10][33] ;
 wire \core.keymem.key_mem[10][34] ;
 wire \core.keymem.key_mem[10][35] ;
 wire \core.keymem.key_mem[10][36] ;
 wire \core.keymem.key_mem[10][37] ;
 wire \core.keymem.key_mem[10][38] ;
 wire \core.keymem.key_mem[10][39] ;
 wire \core.keymem.key_mem[10][3] ;
 wire \core.keymem.key_mem[10][40] ;
 wire \core.keymem.key_mem[10][41] ;
 wire \core.keymem.key_mem[10][42] ;
 wire \core.keymem.key_mem[10][43] ;
 wire \core.keymem.key_mem[10][44] ;
 wire \core.keymem.key_mem[10][45] ;
 wire \core.keymem.key_mem[10][46] ;
 wire \core.keymem.key_mem[10][47] ;
 wire \core.keymem.key_mem[10][48] ;
 wire \core.keymem.key_mem[10][49] ;
 wire \core.keymem.key_mem[10][4] ;
 wire \core.keymem.key_mem[10][50] ;
 wire \core.keymem.key_mem[10][51] ;
 wire \core.keymem.key_mem[10][52] ;
 wire \core.keymem.key_mem[10][53] ;
 wire \core.keymem.key_mem[10][54] ;
 wire \core.keymem.key_mem[10][55] ;
 wire \core.keymem.key_mem[10][56] ;
 wire \core.keymem.key_mem[10][57] ;
 wire \core.keymem.key_mem[10][58] ;
 wire \core.keymem.key_mem[10][59] ;
 wire \core.keymem.key_mem[10][5] ;
 wire \core.keymem.key_mem[10][60] ;
 wire \core.keymem.key_mem[10][61] ;
 wire \core.keymem.key_mem[10][62] ;
 wire \core.keymem.key_mem[10][63] ;
 wire \core.keymem.key_mem[10][64] ;
 wire \core.keymem.key_mem[10][65] ;
 wire \core.keymem.key_mem[10][66] ;
 wire \core.keymem.key_mem[10][67] ;
 wire \core.keymem.key_mem[10][68] ;
 wire \core.keymem.key_mem[10][69] ;
 wire \core.keymem.key_mem[10][6] ;
 wire \core.keymem.key_mem[10][70] ;
 wire \core.keymem.key_mem[10][71] ;
 wire \core.keymem.key_mem[10][72] ;
 wire \core.keymem.key_mem[10][73] ;
 wire \core.keymem.key_mem[10][74] ;
 wire \core.keymem.key_mem[10][75] ;
 wire \core.keymem.key_mem[10][76] ;
 wire \core.keymem.key_mem[10][77] ;
 wire \core.keymem.key_mem[10][78] ;
 wire \core.keymem.key_mem[10][79] ;
 wire \core.keymem.key_mem[10][7] ;
 wire \core.keymem.key_mem[10][80] ;
 wire \core.keymem.key_mem[10][81] ;
 wire \core.keymem.key_mem[10][82] ;
 wire \core.keymem.key_mem[10][83] ;
 wire \core.keymem.key_mem[10][84] ;
 wire \core.keymem.key_mem[10][85] ;
 wire \core.keymem.key_mem[10][86] ;
 wire \core.keymem.key_mem[10][87] ;
 wire \core.keymem.key_mem[10][88] ;
 wire \core.keymem.key_mem[10][89] ;
 wire \core.keymem.key_mem[10][8] ;
 wire \core.keymem.key_mem[10][90] ;
 wire \core.keymem.key_mem[10][91] ;
 wire \core.keymem.key_mem[10][92] ;
 wire \core.keymem.key_mem[10][93] ;
 wire \core.keymem.key_mem[10][94] ;
 wire \core.keymem.key_mem[10][95] ;
 wire \core.keymem.key_mem[10][96] ;
 wire \core.keymem.key_mem[10][97] ;
 wire \core.keymem.key_mem[10][98] ;
 wire \core.keymem.key_mem[10][99] ;
 wire \core.keymem.key_mem[10][9] ;
 wire \core.keymem.key_mem[11][0] ;
 wire \core.keymem.key_mem[11][100] ;
 wire \core.keymem.key_mem[11][101] ;
 wire \core.keymem.key_mem[11][102] ;
 wire \core.keymem.key_mem[11][103] ;
 wire \core.keymem.key_mem[11][104] ;
 wire \core.keymem.key_mem[11][105] ;
 wire \core.keymem.key_mem[11][106] ;
 wire \core.keymem.key_mem[11][107] ;
 wire \core.keymem.key_mem[11][108] ;
 wire \core.keymem.key_mem[11][109] ;
 wire \core.keymem.key_mem[11][10] ;
 wire \core.keymem.key_mem[11][110] ;
 wire \core.keymem.key_mem[11][111] ;
 wire \core.keymem.key_mem[11][112] ;
 wire \core.keymem.key_mem[11][113] ;
 wire \core.keymem.key_mem[11][114] ;
 wire \core.keymem.key_mem[11][115] ;
 wire \core.keymem.key_mem[11][116] ;
 wire \core.keymem.key_mem[11][117] ;
 wire \core.keymem.key_mem[11][118] ;
 wire \core.keymem.key_mem[11][119] ;
 wire \core.keymem.key_mem[11][11] ;
 wire \core.keymem.key_mem[11][120] ;
 wire \core.keymem.key_mem[11][121] ;
 wire \core.keymem.key_mem[11][122] ;
 wire \core.keymem.key_mem[11][123] ;
 wire \core.keymem.key_mem[11][124] ;
 wire \core.keymem.key_mem[11][125] ;
 wire \core.keymem.key_mem[11][126] ;
 wire \core.keymem.key_mem[11][127] ;
 wire \core.keymem.key_mem[11][12] ;
 wire \core.keymem.key_mem[11][13] ;
 wire \core.keymem.key_mem[11][14] ;
 wire \core.keymem.key_mem[11][15] ;
 wire \core.keymem.key_mem[11][16] ;
 wire \core.keymem.key_mem[11][17] ;
 wire \core.keymem.key_mem[11][18] ;
 wire \core.keymem.key_mem[11][19] ;
 wire \core.keymem.key_mem[11][1] ;
 wire \core.keymem.key_mem[11][20] ;
 wire \core.keymem.key_mem[11][21] ;
 wire \core.keymem.key_mem[11][22] ;
 wire \core.keymem.key_mem[11][23] ;
 wire \core.keymem.key_mem[11][24] ;
 wire \core.keymem.key_mem[11][25] ;
 wire \core.keymem.key_mem[11][26] ;
 wire \core.keymem.key_mem[11][27] ;
 wire \core.keymem.key_mem[11][28] ;
 wire \core.keymem.key_mem[11][29] ;
 wire \core.keymem.key_mem[11][2] ;
 wire \core.keymem.key_mem[11][30] ;
 wire \core.keymem.key_mem[11][31] ;
 wire \core.keymem.key_mem[11][32] ;
 wire \core.keymem.key_mem[11][33] ;
 wire \core.keymem.key_mem[11][34] ;
 wire \core.keymem.key_mem[11][35] ;
 wire \core.keymem.key_mem[11][36] ;
 wire \core.keymem.key_mem[11][37] ;
 wire \core.keymem.key_mem[11][38] ;
 wire \core.keymem.key_mem[11][39] ;
 wire \core.keymem.key_mem[11][3] ;
 wire \core.keymem.key_mem[11][40] ;
 wire \core.keymem.key_mem[11][41] ;
 wire \core.keymem.key_mem[11][42] ;
 wire \core.keymem.key_mem[11][43] ;
 wire \core.keymem.key_mem[11][44] ;
 wire \core.keymem.key_mem[11][45] ;
 wire \core.keymem.key_mem[11][46] ;
 wire \core.keymem.key_mem[11][47] ;
 wire \core.keymem.key_mem[11][48] ;
 wire \core.keymem.key_mem[11][49] ;
 wire \core.keymem.key_mem[11][4] ;
 wire \core.keymem.key_mem[11][50] ;
 wire \core.keymem.key_mem[11][51] ;
 wire \core.keymem.key_mem[11][52] ;
 wire \core.keymem.key_mem[11][53] ;
 wire \core.keymem.key_mem[11][54] ;
 wire \core.keymem.key_mem[11][55] ;
 wire \core.keymem.key_mem[11][56] ;
 wire \core.keymem.key_mem[11][57] ;
 wire \core.keymem.key_mem[11][58] ;
 wire \core.keymem.key_mem[11][59] ;
 wire \core.keymem.key_mem[11][5] ;
 wire \core.keymem.key_mem[11][60] ;
 wire \core.keymem.key_mem[11][61] ;
 wire \core.keymem.key_mem[11][62] ;
 wire \core.keymem.key_mem[11][63] ;
 wire \core.keymem.key_mem[11][64] ;
 wire \core.keymem.key_mem[11][65] ;
 wire \core.keymem.key_mem[11][66] ;
 wire \core.keymem.key_mem[11][67] ;
 wire \core.keymem.key_mem[11][68] ;
 wire \core.keymem.key_mem[11][69] ;
 wire \core.keymem.key_mem[11][6] ;
 wire \core.keymem.key_mem[11][70] ;
 wire \core.keymem.key_mem[11][71] ;
 wire \core.keymem.key_mem[11][72] ;
 wire \core.keymem.key_mem[11][73] ;
 wire \core.keymem.key_mem[11][74] ;
 wire \core.keymem.key_mem[11][75] ;
 wire \core.keymem.key_mem[11][76] ;
 wire \core.keymem.key_mem[11][77] ;
 wire \core.keymem.key_mem[11][78] ;
 wire \core.keymem.key_mem[11][79] ;
 wire \core.keymem.key_mem[11][7] ;
 wire \core.keymem.key_mem[11][80] ;
 wire \core.keymem.key_mem[11][81] ;
 wire \core.keymem.key_mem[11][82] ;
 wire \core.keymem.key_mem[11][83] ;
 wire \core.keymem.key_mem[11][84] ;
 wire \core.keymem.key_mem[11][85] ;
 wire \core.keymem.key_mem[11][86] ;
 wire \core.keymem.key_mem[11][87] ;
 wire \core.keymem.key_mem[11][88] ;
 wire \core.keymem.key_mem[11][89] ;
 wire \core.keymem.key_mem[11][8] ;
 wire \core.keymem.key_mem[11][90] ;
 wire \core.keymem.key_mem[11][91] ;
 wire \core.keymem.key_mem[11][92] ;
 wire \core.keymem.key_mem[11][93] ;
 wire \core.keymem.key_mem[11][94] ;
 wire \core.keymem.key_mem[11][95] ;
 wire \core.keymem.key_mem[11][96] ;
 wire \core.keymem.key_mem[11][97] ;
 wire \core.keymem.key_mem[11][98] ;
 wire \core.keymem.key_mem[11][99] ;
 wire \core.keymem.key_mem[11][9] ;
 wire \core.keymem.key_mem[12][0] ;
 wire \core.keymem.key_mem[12][100] ;
 wire \core.keymem.key_mem[12][101] ;
 wire \core.keymem.key_mem[12][102] ;
 wire \core.keymem.key_mem[12][103] ;
 wire \core.keymem.key_mem[12][104] ;
 wire \core.keymem.key_mem[12][105] ;
 wire \core.keymem.key_mem[12][106] ;
 wire \core.keymem.key_mem[12][107] ;
 wire \core.keymem.key_mem[12][108] ;
 wire \core.keymem.key_mem[12][109] ;
 wire \core.keymem.key_mem[12][10] ;
 wire \core.keymem.key_mem[12][110] ;
 wire \core.keymem.key_mem[12][111] ;
 wire \core.keymem.key_mem[12][112] ;
 wire \core.keymem.key_mem[12][113] ;
 wire \core.keymem.key_mem[12][114] ;
 wire \core.keymem.key_mem[12][115] ;
 wire \core.keymem.key_mem[12][116] ;
 wire \core.keymem.key_mem[12][117] ;
 wire \core.keymem.key_mem[12][118] ;
 wire \core.keymem.key_mem[12][119] ;
 wire \core.keymem.key_mem[12][11] ;
 wire \core.keymem.key_mem[12][120] ;
 wire \core.keymem.key_mem[12][121] ;
 wire \core.keymem.key_mem[12][122] ;
 wire \core.keymem.key_mem[12][123] ;
 wire \core.keymem.key_mem[12][124] ;
 wire \core.keymem.key_mem[12][125] ;
 wire \core.keymem.key_mem[12][126] ;
 wire \core.keymem.key_mem[12][127] ;
 wire \core.keymem.key_mem[12][12] ;
 wire \core.keymem.key_mem[12][13] ;
 wire \core.keymem.key_mem[12][14] ;
 wire \core.keymem.key_mem[12][15] ;
 wire \core.keymem.key_mem[12][16] ;
 wire \core.keymem.key_mem[12][17] ;
 wire \core.keymem.key_mem[12][18] ;
 wire \core.keymem.key_mem[12][19] ;
 wire \core.keymem.key_mem[12][1] ;
 wire \core.keymem.key_mem[12][20] ;
 wire \core.keymem.key_mem[12][21] ;
 wire \core.keymem.key_mem[12][22] ;
 wire \core.keymem.key_mem[12][23] ;
 wire \core.keymem.key_mem[12][24] ;
 wire \core.keymem.key_mem[12][25] ;
 wire \core.keymem.key_mem[12][26] ;
 wire \core.keymem.key_mem[12][27] ;
 wire \core.keymem.key_mem[12][28] ;
 wire \core.keymem.key_mem[12][29] ;
 wire \core.keymem.key_mem[12][2] ;
 wire \core.keymem.key_mem[12][30] ;
 wire \core.keymem.key_mem[12][31] ;
 wire \core.keymem.key_mem[12][32] ;
 wire \core.keymem.key_mem[12][33] ;
 wire \core.keymem.key_mem[12][34] ;
 wire \core.keymem.key_mem[12][35] ;
 wire \core.keymem.key_mem[12][36] ;
 wire \core.keymem.key_mem[12][37] ;
 wire \core.keymem.key_mem[12][38] ;
 wire \core.keymem.key_mem[12][39] ;
 wire \core.keymem.key_mem[12][3] ;
 wire \core.keymem.key_mem[12][40] ;
 wire \core.keymem.key_mem[12][41] ;
 wire \core.keymem.key_mem[12][42] ;
 wire \core.keymem.key_mem[12][43] ;
 wire \core.keymem.key_mem[12][44] ;
 wire \core.keymem.key_mem[12][45] ;
 wire \core.keymem.key_mem[12][46] ;
 wire \core.keymem.key_mem[12][47] ;
 wire \core.keymem.key_mem[12][48] ;
 wire \core.keymem.key_mem[12][49] ;
 wire \core.keymem.key_mem[12][4] ;
 wire \core.keymem.key_mem[12][50] ;
 wire \core.keymem.key_mem[12][51] ;
 wire \core.keymem.key_mem[12][52] ;
 wire \core.keymem.key_mem[12][53] ;
 wire \core.keymem.key_mem[12][54] ;
 wire \core.keymem.key_mem[12][55] ;
 wire \core.keymem.key_mem[12][56] ;
 wire \core.keymem.key_mem[12][57] ;
 wire \core.keymem.key_mem[12][58] ;
 wire \core.keymem.key_mem[12][59] ;
 wire \core.keymem.key_mem[12][5] ;
 wire \core.keymem.key_mem[12][60] ;
 wire \core.keymem.key_mem[12][61] ;
 wire \core.keymem.key_mem[12][62] ;
 wire \core.keymem.key_mem[12][63] ;
 wire \core.keymem.key_mem[12][64] ;
 wire \core.keymem.key_mem[12][65] ;
 wire \core.keymem.key_mem[12][66] ;
 wire \core.keymem.key_mem[12][67] ;
 wire \core.keymem.key_mem[12][68] ;
 wire \core.keymem.key_mem[12][69] ;
 wire \core.keymem.key_mem[12][6] ;
 wire \core.keymem.key_mem[12][70] ;
 wire \core.keymem.key_mem[12][71] ;
 wire \core.keymem.key_mem[12][72] ;
 wire \core.keymem.key_mem[12][73] ;
 wire \core.keymem.key_mem[12][74] ;
 wire \core.keymem.key_mem[12][75] ;
 wire \core.keymem.key_mem[12][76] ;
 wire \core.keymem.key_mem[12][77] ;
 wire \core.keymem.key_mem[12][78] ;
 wire \core.keymem.key_mem[12][79] ;
 wire \core.keymem.key_mem[12][7] ;
 wire \core.keymem.key_mem[12][80] ;
 wire \core.keymem.key_mem[12][81] ;
 wire \core.keymem.key_mem[12][82] ;
 wire \core.keymem.key_mem[12][83] ;
 wire \core.keymem.key_mem[12][84] ;
 wire \core.keymem.key_mem[12][85] ;
 wire \core.keymem.key_mem[12][86] ;
 wire \core.keymem.key_mem[12][87] ;
 wire \core.keymem.key_mem[12][88] ;
 wire \core.keymem.key_mem[12][89] ;
 wire \core.keymem.key_mem[12][8] ;
 wire \core.keymem.key_mem[12][90] ;
 wire \core.keymem.key_mem[12][91] ;
 wire \core.keymem.key_mem[12][92] ;
 wire \core.keymem.key_mem[12][93] ;
 wire \core.keymem.key_mem[12][94] ;
 wire \core.keymem.key_mem[12][95] ;
 wire \core.keymem.key_mem[12][96] ;
 wire \core.keymem.key_mem[12][97] ;
 wire \core.keymem.key_mem[12][98] ;
 wire \core.keymem.key_mem[12][99] ;
 wire \core.keymem.key_mem[12][9] ;
 wire \core.keymem.key_mem[13][0] ;
 wire \core.keymem.key_mem[13][100] ;
 wire \core.keymem.key_mem[13][101] ;
 wire \core.keymem.key_mem[13][102] ;
 wire \core.keymem.key_mem[13][103] ;
 wire \core.keymem.key_mem[13][104] ;
 wire \core.keymem.key_mem[13][105] ;
 wire \core.keymem.key_mem[13][106] ;
 wire \core.keymem.key_mem[13][107] ;
 wire \core.keymem.key_mem[13][108] ;
 wire \core.keymem.key_mem[13][109] ;
 wire \core.keymem.key_mem[13][10] ;
 wire \core.keymem.key_mem[13][110] ;
 wire \core.keymem.key_mem[13][111] ;
 wire \core.keymem.key_mem[13][112] ;
 wire \core.keymem.key_mem[13][113] ;
 wire \core.keymem.key_mem[13][114] ;
 wire \core.keymem.key_mem[13][115] ;
 wire \core.keymem.key_mem[13][116] ;
 wire \core.keymem.key_mem[13][117] ;
 wire \core.keymem.key_mem[13][118] ;
 wire \core.keymem.key_mem[13][119] ;
 wire \core.keymem.key_mem[13][11] ;
 wire \core.keymem.key_mem[13][120] ;
 wire \core.keymem.key_mem[13][121] ;
 wire \core.keymem.key_mem[13][122] ;
 wire \core.keymem.key_mem[13][123] ;
 wire \core.keymem.key_mem[13][124] ;
 wire \core.keymem.key_mem[13][125] ;
 wire \core.keymem.key_mem[13][126] ;
 wire \core.keymem.key_mem[13][127] ;
 wire \core.keymem.key_mem[13][12] ;
 wire \core.keymem.key_mem[13][13] ;
 wire \core.keymem.key_mem[13][14] ;
 wire \core.keymem.key_mem[13][15] ;
 wire \core.keymem.key_mem[13][16] ;
 wire \core.keymem.key_mem[13][17] ;
 wire \core.keymem.key_mem[13][18] ;
 wire \core.keymem.key_mem[13][19] ;
 wire \core.keymem.key_mem[13][1] ;
 wire \core.keymem.key_mem[13][20] ;
 wire \core.keymem.key_mem[13][21] ;
 wire \core.keymem.key_mem[13][22] ;
 wire \core.keymem.key_mem[13][23] ;
 wire \core.keymem.key_mem[13][24] ;
 wire \core.keymem.key_mem[13][25] ;
 wire \core.keymem.key_mem[13][26] ;
 wire \core.keymem.key_mem[13][27] ;
 wire \core.keymem.key_mem[13][28] ;
 wire \core.keymem.key_mem[13][29] ;
 wire \core.keymem.key_mem[13][2] ;
 wire \core.keymem.key_mem[13][30] ;
 wire \core.keymem.key_mem[13][31] ;
 wire \core.keymem.key_mem[13][32] ;
 wire \core.keymem.key_mem[13][33] ;
 wire \core.keymem.key_mem[13][34] ;
 wire \core.keymem.key_mem[13][35] ;
 wire \core.keymem.key_mem[13][36] ;
 wire \core.keymem.key_mem[13][37] ;
 wire \core.keymem.key_mem[13][38] ;
 wire \core.keymem.key_mem[13][39] ;
 wire \core.keymem.key_mem[13][3] ;
 wire \core.keymem.key_mem[13][40] ;
 wire \core.keymem.key_mem[13][41] ;
 wire \core.keymem.key_mem[13][42] ;
 wire \core.keymem.key_mem[13][43] ;
 wire \core.keymem.key_mem[13][44] ;
 wire \core.keymem.key_mem[13][45] ;
 wire \core.keymem.key_mem[13][46] ;
 wire \core.keymem.key_mem[13][47] ;
 wire \core.keymem.key_mem[13][48] ;
 wire \core.keymem.key_mem[13][49] ;
 wire \core.keymem.key_mem[13][4] ;
 wire \core.keymem.key_mem[13][50] ;
 wire \core.keymem.key_mem[13][51] ;
 wire \core.keymem.key_mem[13][52] ;
 wire \core.keymem.key_mem[13][53] ;
 wire \core.keymem.key_mem[13][54] ;
 wire \core.keymem.key_mem[13][55] ;
 wire \core.keymem.key_mem[13][56] ;
 wire \core.keymem.key_mem[13][57] ;
 wire \core.keymem.key_mem[13][58] ;
 wire \core.keymem.key_mem[13][59] ;
 wire \core.keymem.key_mem[13][5] ;
 wire \core.keymem.key_mem[13][60] ;
 wire \core.keymem.key_mem[13][61] ;
 wire \core.keymem.key_mem[13][62] ;
 wire \core.keymem.key_mem[13][63] ;
 wire \core.keymem.key_mem[13][64] ;
 wire \core.keymem.key_mem[13][65] ;
 wire \core.keymem.key_mem[13][66] ;
 wire \core.keymem.key_mem[13][67] ;
 wire \core.keymem.key_mem[13][68] ;
 wire \core.keymem.key_mem[13][69] ;
 wire \core.keymem.key_mem[13][6] ;
 wire \core.keymem.key_mem[13][70] ;
 wire \core.keymem.key_mem[13][71] ;
 wire \core.keymem.key_mem[13][72] ;
 wire \core.keymem.key_mem[13][73] ;
 wire \core.keymem.key_mem[13][74] ;
 wire \core.keymem.key_mem[13][75] ;
 wire \core.keymem.key_mem[13][76] ;
 wire \core.keymem.key_mem[13][77] ;
 wire \core.keymem.key_mem[13][78] ;
 wire \core.keymem.key_mem[13][79] ;
 wire \core.keymem.key_mem[13][7] ;
 wire \core.keymem.key_mem[13][80] ;
 wire \core.keymem.key_mem[13][81] ;
 wire \core.keymem.key_mem[13][82] ;
 wire \core.keymem.key_mem[13][83] ;
 wire \core.keymem.key_mem[13][84] ;
 wire \core.keymem.key_mem[13][85] ;
 wire \core.keymem.key_mem[13][86] ;
 wire \core.keymem.key_mem[13][87] ;
 wire \core.keymem.key_mem[13][88] ;
 wire \core.keymem.key_mem[13][89] ;
 wire \core.keymem.key_mem[13][8] ;
 wire \core.keymem.key_mem[13][90] ;
 wire \core.keymem.key_mem[13][91] ;
 wire \core.keymem.key_mem[13][92] ;
 wire \core.keymem.key_mem[13][93] ;
 wire \core.keymem.key_mem[13][94] ;
 wire \core.keymem.key_mem[13][95] ;
 wire \core.keymem.key_mem[13][96] ;
 wire \core.keymem.key_mem[13][97] ;
 wire \core.keymem.key_mem[13][98] ;
 wire \core.keymem.key_mem[13][99] ;
 wire \core.keymem.key_mem[13][9] ;
 wire \core.keymem.key_mem[14][0] ;
 wire \core.keymem.key_mem[14][100] ;
 wire \core.keymem.key_mem[14][101] ;
 wire \core.keymem.key_mem[14][102] ;
 wire \core.keymem.key_mem[14][103] ;
 wire \core.keymem.key_mem[14][104] ;
 wire \core.keymem.key_mem[14][105] ;
 wire \core.keymem.key_mem[14][106] ;
 wire \core.keymem.key_mem[14][107] ;
 wire \core.keymem.key_mem[14][108] ;
 wire \core.keymem.key_mem[14][109] ;
 wire \core.keymem.key_mem[14][10] ;
 wire \core.keymem.key_mem[14][110] ;
 wire \core.keymem.key_mem[14][111] ;
 wire \core.keymem.key_mem[14][112] ;
 wire \core.keymem.key_mem[14][113] ;
 wire \core.keymem.key_mem[14][114] ;
 wire \core.keymem.key_mem[14][115] ;
 wire \core.keymem.key_mem[14][116] ;
 wire \core.keymem.key_mem[14][117] ;
 wire \core.keymem.key_mem[14][118] ;
 wire \core.keymem.key_mem[14][119] ;
 wire \core.keymem.key_mem[14][11] ;
 wire \core.keymem.key_mem[14][120] ;
 wire \core.keymem.key_mem[14][121] ;
 wire \core.keymem.key_mem[14][122] ;
 wire \core.keymem.key_mem[14][123] ;
 wire \core.keymem.key_mem[14][124] ;
 wire \core.keymem.key_mem[14][125] ;
 wire \core.keymem.key_mem[14][126] ;
 wire \core.keymem.key_mem[14][127] ;
 wire \core.keymem.key_mem[14][12] ;
 wire \core.keymem.key_mem[14][13] ;
 wire \core.keymem.key_mem[14][14] ;
 wire \core.keymem.key_mem[14][15] ;
 wire \core.keymem.key_mem[14][16] ;
 wire \core.keymem.key_mem[14][17] ;
 wire \core.keymem.key_mem[14][18] ;
 wire \core.keymem.key_mem[14][19] ;
 wire \core.keymem.key_mem[14][1] ;
 wire \core.keymem.key_mem[14][20] ;
 wire \core.keymem.key_mem[14][21] ;
 wire \core.keymem.key_mem[14][22] ;
 wire \core.keymem.key_mem[14][23] ;
 wire \core.keymem.key_mem[14][24] ;
 wire \core.keymem.key_mem[14][25] ;
 wire \core.keymem.key_mem[14][26] ;
 wire \core.keymem.key_mem[14][27] ;
 wire \core.keymem.key_mem[14][28] ;
 wire \core.keymem.key_mem[14][29] ;
 wire \core.keymem.key_mem[14][2] ;
 wire \core.keymem.key_mem[14][30] ;
 wire \core.keymem.key_mem[14][31] ;
 wire \core.keymem.key_mem[14][32] ;
 wire \core.keymem.key_mem[14][33] ;
 wire \core.keymem.key_mem[14][34] ;
 wire \core.keymem.key_mem[14][35] ;
 wire \core.keymem.key_mem[14][36] ;
 wire \core.keymem.key_mem[14][37] ;
 wire \core.keymem.key_mem[14][38] ;
 wire \core.keymem.key_mem[14][39] ;
 wire \core.keymem.key_mem[14][3] ;
 wire \core.keymem.key_mem[14][40] ;
 wire \core.keymem.key_mem[14][41] ;
 wire \core.keymem.key_mem[14][42] ;
 wire \core.keymem.key_mem[14][43] ;
 wire \core.keymem.key_mem[14][44] ;
 wire \core.keymem.key_mem[14][45] ;
 wire \core.keymem.key_mem[14][46] ;
 wire \core.keymem.key_mem[14][47] ;
 wire \core.keymem.key_mem[14][48] ;
 wire \core.keymem.key_mem[14][49] ;
 wire \core.keymem.key_mem[14][4] ;
 wire \core.keymem.key_mem[14][50] ;
 wire \core.keymem.key_mem[14][51] ;
 wire \core.keymem.key_mem[14][52] ;
 wire \core.keymem.key_mem[14][53] ;
 wire \core.keymem.key_mem[14][54] ;
 wire \core.keymem.key_mem[14][55] ;
 wire \core.keymem.key_mem[14][56] ;
 wire \core.keymem.key_mem[14][57] ;
 wire \core.keymem.key_mem[14][58] ;
 wire \core.keymem.key_mem[14][59] ;
 wire \core.keymem.key_mem[14][5] ;
 wire \core.keymem.key_mem[14][60] ;
 wire \core.keymem.key_mem[14][61] ;
 wire \core.keymem.key_mem[14][62] ;
 wire \core.keymem.key_mem[14][63] ;
 wire \core.keymem.key_mem[14][64] ;
 wire \core.keymem.key_mem[14][65] ;
 wire \core.keymem.key_mem[14][66] ;
 wire \core.keymem.key_mem[14][67] ;
 wire \core.keymem.key_mem[14][68] ;
 wire \core.keymem.key_mem[14][69] ;
 wire \core.keymem.key_mem[14][6] ;
 wire \core.keymem.key_mem[14][70] ;
 wire \core.keymem.key_mem[14][71] ;
 wire \core.keymem.key_mem[14][72] ;
 wire \core.keymem.key_mem[14][73] ;
 wire \core.keymem.key_mem[14][74] ;
 wire \core.keymem.key_mem[14][75] ;
 wire \core.keymem.key_mem[14][76] ;
 wire \core.keymem.key_mem[14][77] ;
 wire \core.keymem.key_mem[14][78] ;
 wire \core.keymem.key_mem[14][79] ;
 wire \core.keymem.key_mem[14][7] ;
 wire \core.keymem.key_mem[14][80] ;
 wire \core.keymem.key_mem[14][81] ;
 wire \core.keymem.key_mem[14][82] ;
 wire \core.keymem.key_mem[14][83] ;
 wire \core.keymem.key_mem[14][84] ;
 wire \core.keymem.key_mem[14][85] ;
 wire \core.keymem.key_mem[14][86] ;
 wire \core.keymem.key_mem[14][87] ;
 wire \core.keymem.key_mem[14][88] ;
 wire \core.keymem.key_mem[14][89] ;
 wire \core.keymem.key_mem[14][8] ;
 wire \core.keymem.key_mem[14][90] ;
 wire \core.keymem.key_mem[14][91] ;
 wire \core.keymem.key_mem[14][92] ;
 wire \core.keymem.key_mem[14][93] ;
 wire \core.keymem.key_mem[14][94] ;
 wire \core.keymem.key_mem[14][95] ;
 wire \core.keymem.key_mem[14][96] ;
 wire \core.keymem.key_mem[14][97] ;
 wire \core.keymem.key_mem[14][98] ;
 wire \core.keymem.key_mem[14][99] ;
 wire \core.keymem.key_mem[14][9] ;
 wire \core.keymem.key_mem[1][0] ;
 wire \core.keymem.key_mem[1][100] ;
 wire \core.keymem.key_mem[1][101] ;
 wire \core.keymem.key_mem[1][102] ;
 wire \core.keymem.key_mem[1][103] ;
 wire \core.keymem.key_mem[1][104] ;
 wire \core.keymem.key_mem[1][105] ;
 wire \core.keymem.key_mem[1][106] ;
 wire \core.keymem.key_mem[1][107] ;
 wire \core.keymem.key_mem[1][108] ;
 wire \core.keymem.key_mem[1][109] ;
 wire \core.keymem.key_mem[1][10] ;
 wire \core.keymem.key_mem[1][110] ;
 wire \core.keymem.key_mem[1][111] ;
 wire \core.keymem.key_mem[1][112] ;
 wire \core.keymem.key_mem[1][113] ;
 wire \core.keymem.key_mem[1][114] ;
 wire \core.keymem.key_mem[1][115] ;
 wire \core.keymem.key_mem[1][116] ;
 wire \core.keymem.key_mem[1][117] ;
 wire \core.keymem.key_mem[1][118] ;
 wire \core.keymem.key_mem[1][119] ;
 wire \core.keymem.key_mem[1][11] ;
 wire \core.keymem.key_mem[1][120] ;
 wire \core.keymem.key_mem[1][121] ;
 wire \core.keymem.key_mem[1][122] ;
 wire \core.keymem.key_mem[1][123] ;
 wire \core.keymem.key_mem[1][124] ;
 wire \core.keymem.key_mem[1][125] ;
 wire \core.keymem.key_mem[1][126] ;
 wire \core.keymem.key_mem[1][127] ;
 wire \core.keymem.key_mem[1][12] ;
 wire \core.keymem.key_mem[1][13] ;
 wire \core.keymem.key_mem[1][14] ;
 wire \core.keymem.key_mem[1][15] ;
 wire \core.keymem.key_mem[1][16] ;
 wire \core.keymem.key_mem[1][17] ;
 wire \core.keymem.key_mem[1][18] ;
 wire \core.keymem.key_mem[1][19] ;
 wire \core.keymem.key_mem[1][1] ;
 wire \core.keymem.key_mem[1][20] ;
 wire \core.keymem.key_mem[1][21] ;
 wire \core.keymem.key_mem[1][22] ;
 wire \core.keymem.key_mem[1][23] ;
 wire \core.keymem.key_mem[1][24] ;
 wire \core.keymem.key_mem[1][25] ;
 wire \core.keymem.key_mem[1][26] ;
 wire \core.keymem.key_mem[1][27] ;
 wire \core.keymem.key_mem[1][28] ;
 wire \core.keymem.key_mem[1][29] ;
 wire \core.keymem.key_mem[1][2] ;
 wire \core.keymem.key_mem[1][30] ;
 wire \core.keymem.key_mem[1][31] ;
 wire \core.keymem.key_mem[1][32] ;
 wire \core.keymem.key_mem[1][33] ;
 wire \core.keymem.key_mem[1][34] ;
 wire \core.keymem.key_mem[1][35] ;
 wire \core.keymem.key_mem[1][36] ;
 wire \core.keymem.key_mem[1][37] ;
 wire \core.keymem.key_mem[1][38] ;
 wire \core.keymem.key_mem[1][39] ;
 wire \core.keymem.key_mem[1][3] ;
 wire \core.keymem.key_mem[1][40] ;
 wire \core.keymem.key_mem[1][41] ;
 wire \core.keymem.key_mem[1][42] ;
 wire \core.keymem.key_mem[1][43] ;
 wire \core.keymem.key_mem[1][44] ;
 wire \core.keymem.key_mem[1][45] ;
 wire \core.keymem.key_mem[1][46] ;
 wire \core.keymem.key_mem[1][47] ;
 wire \core.keymem.key_mem[1][48] ;
 wire \core.keymem.key_mem[1][49] ;
 wire \core.keymem.key_mem[1][4] ;
 wire \core.keymem.key_mem[1][50] ;
 wire \core.keymem.key_mem[1][51] ;
 wire \core.keymem.key_mem[1][52] ;
 wire \core.keymem.key_mem[1][53] ;
 wire \core.keymem.key_mem[1][54] ;
 wire \core.keymem.key_mem[1][55] ;
 wire \core.keymem.key_mem[1][56] ;
 wire \core.keymem.key_mem[1][57] ;
 wire \core.keymem.key_mem[1][58] ;
 wire \core.keymem.key_mem[1][59] ;
 wire \core.keymem.key_mem[1][5] ;
 wire \core.keymem.key_mem[1][60] ;
 wire \core.keymem.key_mem[1][61] ;
 wire \core.keymem.key_mem[1][62] ;
 wire \core.keymem.key_mem[1][63] ;
 wire \core.keymem.key_mem[1][64] ;
 wire \core.keymem.key_mem[1][65] ;
 wire \core.keymem.key_mem[1][66] ;
 wire \core.keymem.key_mem[1][67] ;
 wire \core.keymem.key_mem[1][68] ;
 wire \core.keymem.key_mem[1][69] ;
 wire \core.keymem.key_mem[1][6] ;
 wire \core.keymem.key_mem[1][70] ;
 wire \core.keymem.key_mem[1][71] ;
 wire \core.keymem.key_mem[1][72] ;
 wire \core.keymem.key_mem[1][73] ;
 wire \core.keymem.key_mem[1][74] ;
 wire \core.keymem.key_mem[1][75] ;
 wire \core.keymem.key_mem[1][76] ;
 wire \core.keymem.key_mem[1][77] ;
 wire \core.keymem.key_mem[1][78] ;
 wire \core.keymem.key_mem[1][79] ;
 wire \core.keymem.key_mem[1][7] ;
 wire \core.keymem.key_mem[1][80] ;
 wire \core.keymem.key_mem[1][81] ;
 wire \core.keymem.key_mem[1][82] ;
 wire \core.keymem.key_mem[1][83] ;
 wire \core.keymem.key_mem[1][84] ;
 wire \core.keymem.key_mem[1][85] ;
 wire \core.keymem.key_mem[1][86] ;
 wire \core.keymem.key_mem[1][87] ;
 wire \core.keymem.key_mem[1][88] ;
 wire \core.keymem.key_mem[1][89] ;
 wire \core.keymem.key_mem[1][8] ;
 wire \core.keymem.key_mem[1][90] ;
 wire \core.keymem.key_mem[1][91] ;
 wire \core.keymem.key_mem[1][92] ;
 wire \core.keymem.key_mem[1][93] ;
 wire \core.keymem.key_mem[1][94] ;
 wire \core.keymem.key_mem[1][95] ;
 wire \core.keymem.key_mem[1][96] ;
 wire \core.keymem.key_mem[1][97] ;
 wire \core.keymem.key_mem[1][98] ;
 wire \core.keymem.key_mem[1][99] ;
 wire \core.keymem.key_mem[1][9] ;
 wire \core.keymem.key_mem[2][0] ;
 wire \core.keymem.key_mem[2][100] ;
 wire \core.keymem.key_mem[2][101] ;
 wire \core.keymem.key_mem[2][102] ;
 wire \core.keymem.key_mem[2][103] ;
 wire \core.keymem.key_mem[2][104] ;
 wire \core.keymem.key_mem[2][105] ;
 wire \core.keymem.key_mem[2][106] ;
 wire \core.keymem.key_mem[2][107] ;
 wire \core.keymem.key_mem[2][108] ;
 wire \core.keymem.key_mem[2][109] ;
 wire \core.keymem.key_mem[2][10] ;
 wire \core.keymem.key_mem[2][110] ;
 wire \core.keymem.key_mem[2][111] ;
 wire \core.keymem.key_mem[2][112] ;
 wire \core.keymem.key_mem[2][113] ;
 wire \core.keymem.key_mem[2][114] ;
 wire \core.keymem.key_mem[2][115] ;
 wire \core.keymem.key_mem[2][116] ;
 wire \core.keymem.key_mem[2][117] ;
 wire \core.keymem.key_mem[2][118] ;
 wire \core.keymem.key_mem[2][119] ;
 wire \core.keymem.key_mem[2][11] ;
 wire \core.keymem.key_mem[2][120] ;
 wire \core.keymem.key_mem[2][121] ;
 wire \core.keymem.key_mem[2][122] ;
 wire \core.keymem.key_mem[2][123] ;
 wire \core.keymem.key_mem[2][124] ;
 wire \core.keymem.key_mem[2][125] ;
 wire \core.keymem.key_mem[2][126] ;
 wire \core.keymem.key_mem[2][127] ;
 wire \core.keymem.key_mem[2][12] ;
 wire \core.keymem.key_mem[2][13] ;
 wire \core.keymem.key_mem[2][14] ;
 wire \core.keymem.key_mem[2][15] ;
 wire \core.keymem.key_mem[2][16] ;
 wire \core.keymem.key_mem[2][17] ;
 wire \core.keymem.key_mem[2][18] ;
 wire \core.keymem.key_mem[2][19] ;
 wire \core.keymem.key_mem[2][1] ;
 wire \core.keymem.key_mem[2][20] ;
 wire \core.keymem.key_mem[2][21] ;
 wire \core.keymem.key_mem[2][22] ;
 wire \core.keymem.key_mem[2][23] ;
 wire \core.keymem.key_mem[2][24] ;
 wire \core.keymem.key_mem[2][25] ;
 wire \core.keymem.key_mem[2][26] ;
 wire \core.keymem.key_mem[2][27] ;
 wire \core.keymem.key_mem[2][28] ;
 wire \core.keymem.key_mem[2][29] ;
 wire \core.keymem.key_mem[2][2] ;
 wire \core.keymem.key_mem[2][30] ;
 wire \core.keymem.key_mem[2][31] ;
 wire \core.keymem.key_mem[2][32] ;
 wire \core.keymem.key_mem[2][33] ;
 wire \core.keymem.key_mem[2][34] ;
 wire \core.keymem.key_mem[2][35] ;
 wire \core.keymem.key_mem[2][36] ;
 wire \core.keymem.key_mem[2][37] ;
 wire \core.keymem.key_mem[2][38] ;
 wire \core.keymem.key_mem[2][39] ;
 wire \core.keymem.key_mem[2][3] ;
 wire \core.keymem.key_mem[2][40] ;
 wire \core.keymem.key_mem[2][41] ;
 wire \core.keymem.key_mem[2][42] ;
 wire \core.keymem.key_mem[2][43] ;
 wire \core.keymem.key_mem[2][44] ;
 wire \core.keymem.key_mem[2][45] ;
 wire \core.keymem.key_mem[2][46] ;
 wire \core.keymem.key_mem[2][47] ;
 wire \core.keymem.key_mem[2][48] ;
 wire \core.keymem.key_mem[2][49] ;
 wire \core.keymem.key_mem[2][4] ;
 wire \core.keymem.key_mem[2][50] ;
 wire \core.keymem.key_mem[2][51] ;
 wire \core.keymem.key_mem[2][52] ;
 wire \core.keymem.key_mem[2][53] ;
 wire \core.keymem.key_mem[2][54] ;
 wire \core.keymem.key_mem[2][55] ;
 wire \core.keymem.key_mem[2][56] ;
 wire \core.keymem.key_mem[2][57] ;
 wire \core.keymem.key_mem[2][58] ;
 wire \core.keymem.key_mem[2][59] ;
 wire \core.keymem.key_mem[2][5] ;
 wire \core.keymem.key_mem[2][60] ;
 wire \core.keymem.key_mem[2][61] ;
 wire \core.keymem.key_mem[2][62] ;
 wire \core.keymem.key_mem[2][63] ;
 wire \core.keymem.key_mem[2][64] ;
 wire \core.keymem.key_mem[2][65] ;
 wire \core.keymem.key_mem[2][66] ;
 wire \core.keymem.key_mem[2][67] ;
 wire \core.keymem.key_mem[2][68] ;
 wire \core.keymem.key_mem[2][69] ;
 wire \core.keymem.key_mem[2][6] ;
 wire \core.keymem.key_mem[2][70] ;
 wire \core.keymem.key_mem[2][71] ;
 wire \core.keymem.key_mem[2][72] ;
 wire \core.keymem.key_mem[2][73] ;
 wire \core.keymem.key_mem[2][74] ;
 wire \core.keymem.key_mem[2][75] ;
 wire \core.keymem.key_mem[2][76] ;
 wire \core.keymem.key_mem[2][77] ;
 wire \core.keymem.key_mem[2][78] ;
 wire \core.keymem.key_mem[2][79] ;
 wire \core.keymem.key_mem[2][7] ;
 wire \core.keymem.key_mem[2][80] ;
 wire \core.keymem.key_mem[2][81] ;
 wire \core.keymem.key_mem[2][82] ;
 wire \core.keymem.key_mem[2][83] ;
 wire \core.keymem.key_mem[2][84] ;
 wire \core.keymem.key_mem[2][85] ;
 wire \core.keymem.key_mem[2][86] ;
 wire \core.keymem.key_mem[2][87] ;
 wire \core.keymem.key_mem[2][88] ;
 wire \core.keymem.key_mem[2][89] ;
 wire \core.keymem.key_mem[2][8] ;
 wire \core.keymem.key_mem[2][90] ;
 wire \core.keymem.key_mem[2][91] ;
 wire \core.keymem.key_mem[2][92] ;
 wire \core.keymem.key_mem[2][93] ;
 wire \core.keymem.key_mem[2][94] ;
 wire \core.keymem.key_mem[2][95] ;
 wire \core.keymem.key_mem[2][96] ;
 wire \core.keymem.key_mem[2][97] ;
 wire \core.keymem.key_mem[2][98] ;
 wire \core.keymem.key_mem[2][99] ;
 wire \core.keymem.key_mem[2][9] ;
 wire \core.keymem.key_mem[3][0] ;
 wire \core.keymem.key_mem[3][100] ;
 wire \core.keymem.key_mem[3][101] ;
 wire \core.keymem.key_mem[3][102] ;
 wire \core.keymem.key_mem[3][103] ;
 wire \core.keymem.key_mem[3][104] ;
 wire \core.keymem.key_mem[3][105] ;
 wire \core.keymem.key_mem[3][106] ;
 wire \core.keymem.key_mem[3][107] ;
 wire \core.keymem.key_mem[3][108] ;
 wire \core.keymem.key_mem[3][109] ;
 wire \core.keymem.key_mem[3][10] ;
 wire \core.keymem.key_mem[3][110] ;
 wire \core.keymem.key_mem[3][111] ;
 wire \core.keymem.key_mem[3][112] ;
 wire \core.keymem.key_mem[3][113] ;
 wire \core.keymem.key_mem[3][114] ;
 wire \core.keymem.key_mem[3][115] ;
 wire \core.keymem.key_mem[3][116] ;
 wire \core.keymem.key_mem[3][117] ;
 wire \core.keymem.key_mem[3][118] ;
 wire \core.keymem.key_mem[3][119] ;
 wire \core.keymem.key_mem[3][11] ;
 wire \core.keymem.key_mem[3][120] ;
 wire \core.keymem.key_mem[3][121] ;
 wire \core.keymem.key_mem[3][122] ;
 wire \core.keymem.key_mem[3][123] ;
 wire \core.keymem.key_mem[3][124] ;
 wire \core.keymem.key_mem[3][125] ;
 wire \core.keymem.key_mem[3][126] ;
 wire \core.keymem.key_mem[3][127] ;
 wire \core.keymem.key_mem[3][12] ;
 wire \core.keymem.key_mem[3][13] ;
 wire \core.keymem.key_mem[3][14] ;
 wire \core.keymem.key_mem[3][15] ;
 wire \core.keymem.key_mem[3][16] ;
 wire \core.keymem.key_mem[3][17] ;
 wire \core.keymem.key_mem[3][18] ;
 wire \core.keymem.key_mem[3][19] ;
 wire \core.keymem.key_mem[3][1] ;
 wire \core.keymem.key_mem[3][20] ;
 wire \core.keymem.key_mem[3][21] ;
 wire \core.keymem.key_mem[3][22] ;
 wire \core.keymem.key_mem[3][23] ;
 wire \core.keymem.key_mem[3][24] ;
 wire \core.keymem.key_mem[3][25] ;
 wire \core.keymem.key_mem[3][26] ;
 wire \core.keymem.key_mem[3][27] ;
 wire \core.keymem.key_mem[3][28] ;
 wire \core.keymem.key_mem[3][29] ;
 wire \core.keymem.key_mem[3][2] ;
 wire \core.keymem.key_mem[3][30] ;
 wire \core.keymem.key_mem[3][31] ;
 wire \core.keymem.key_mem[3][32] ;
 wire \core.keymem.key_mem[3][33] ;
 wire \core.keymem.key_mem[3][34] ;
 wire \core.keymem.key_mem[3][35] ;
 wire \core.keymem.key_mem[3][36] ;
 wire \core.keymem.key_mem[3][37] ;
 wire \core.keymem.key_mem[3][38] ;
 wire \core.keymem.key_mem[3][39] ;
 wire \core.keymem.key_mem[3][3] ;
 wire \core.keymem.key_mem[3][40] ;
 wire \core.keymem.key_mem[3][41] ;
 wire \core.keymem.key_mem[3][42] ;
 wire \core.keymem.key_mem[3][43] ;
 wire \core.keymem.key_mem[3][44] ;
 wire \core.keymem.key_mem[3][45] ;
 wire \core.keymem.key_mem[3][46] ;
 wire \core.keymem.key_mem[3][47] ;
 wire \core.keymem.key_mem[3][48] ;
 wire \core.keymem.key_mem[3][49] ;
 wire \core.keymem.key_mem[3][4] ;
 wire \core.keymem.key_mem[3][50] ;
 wire \core.keymem.key_mem[3][51] ;
 wire \core.keymem.key_mem[3][52] ;
 wire \core.keymem.key_mem[3][53] ;
 wire \core.keymem.key_mem[3][54] ;
 wire \core.keymem.key_mem[3][55] ;
 wire \core.keymem.key_mem[3][56] ;
 wire \core.keymem.key_mem[3][57] ;
 wire \core.keymem.key_mem[3][58] ;
 wire \core.keymem.key_mem[3][59] ;
 wire \core.keymem.key_mem[3][5] ;
 wire \core.keymem.key_mem[3][60] ;
 wire \core.keymem.key_mem[3][61] ;
 wire \core.keymem.key_mem[3][62] ;
 wire \core.keymem.key_mem[3][63] ;
 wire \core.keymem.key_mem[3][64] ;
 wire \core.keymem.key_mem[3][65] ;
 wire \core.keymem.key_mem[3][66] ;
 wire \core.keymem.key_mem[3][67] ;
 wire \core.keymem.key_mem[3][68] ;
 wire \core.keymem.key_mem[3][69] ;
 wire \core.keymem.key_mem[3][6] ;
 wire \core.keymem.key_mem[3][70] ;
 wire \core.keymem.key_mem[3][71] ;
 wire \core.keymem.key_mem[3][72] ;
 wire \core.keymem.key_mem[3][73] ;
 wire \core.keymem.key_mem[3][74] ;
 wire \core.keymem.key_mem[3][75] ;
 wire \core.keymem.key_mem[3][76] ;
 wire \core.keymem.key_mem[3][77] ;
 wire \core.keymem.key_mem[3][78] ;
 wire \core.keymem.key_mem[3][79] ;
 wire \core.keymem.key_mem[3][7] ;
 wire \core.keymem.key_mem[3][80] ;
 wire \core.keymem.key_mem[3][81] ;
 wire \core.keymem.key_mem[3][82] ;
 wire \core.keymem.key_mem[3][83] ;
 wire \core.keymem.key_mem[3][84] ;
 wire \core.keymem.key_mem[3][85] ;
 wire \core.keymem.key_mem[3][86] ;
 wire \core.keymem.key_mem[3][87] ;
 wire \core.keymem.key_mem[3][88] ;
 wire \core.keymem.key_mem[3][89] ;
 wire \core.keymem.key_mem[3][8] ;
 wire \core.keymem.key_mem[3][90] ;
 wire \core.keymem.key_mem[3][91] ;
 wire \core.keymem.key_mem[3][92] ;
 wire \core.keymem.key_mem[3][93] ;
 wire \core.keymem.key_mem[3][94] ;
 wire \core.keymem.key_mem[3][95] ;
 wire \core.keymem.key_mem[3][96] ;
 wire \core.keymem.key_mem[3][97] ;
 wire \core.keymem.key_mem[3][98] ;
 wire \core.keymem.key_mem[3][99] ;
 wire \core.keymem.key_mem[3][9] ;
 wire \core.keymem.key_mem[4][0] ;
 wire \core.keymem.key_mem[4][100] ;
 wire \core.keymem.key_mem[4][101] ;
 wire \core.keymem.key_mem[4][102] ;
 wire \core.keymem.key_mem[4][103] ;
 wire \core.keymem.key_mem[4][104] ;
 wire \core.keymem.key_mem[4][105] ;
 wire \core.keymem.key_mem[4][106] ;
 wire \core.keymem.key_mem[4][107] ;
 wire \core.keymem.key_mem[4][108] ;
 wire \core.keymem.key_mem[4][109] ;
 wire \core.keymem.key_mem[4][10] ;
 wire \core.keymem.key_mem[4][110] ;
 wire \core.keymem.key_mem[4][111] ;
 wire \core.keymem.key_mem[4][112] ;
 wire \core.keymem.key_mem[4][113] ;
 wire \core.keymem.key_mem[4][114] ;
 wire \core.keymem.key_mem[4][115] ;
 wire \core.keymem.key_mem[4][116] ;
 wire \core.keymem.key_mem[4][117] ;
 wire \core.keymem.key_mem[4][118] ;
 wire \core.keymem.key_mem[4][119] ;
 wire \core.keymem.key_mem[4][11] ;
 wire \core.keymem.key_mem[4][120] ;
 wire \core.keymem.key_mem[4][121] ;
 wire \core.keymem.key_mem[4][122] ;
 wire \core.keymem.key_mem[4][123] ;
 wire \core.keymem.key_mem[4][124] ;
 wire \core.keymem.key_mem[4][125] ;
 wire \core.keymem.key_mem[4][126] ;
 wire \core.keymem.key_mem[4][127] ;
 wire \core.keymem.key_mem[4][12] ;
 wire \core.keymem.key_mem[4][13] ;
 wire \core.keymem.key_mem[4][14] ;
 wire \core.keymem.key_mem[4][15] ;
 wire \core.keymem.key_mem[4][16] ;
 wire \core.keymem.key_mem[4][17] ;
 wire \core.keymem.key_mem[4][18] ;
 wire \core.keymem.key_mem[4][19] ;
 wire \core.keymem.key_mem[4][1] ;
 wire \core.keymem.key_mem[4][20] ;
 wire \core.keymem.key_mem[4][21] ;
 wire \core.keymem.key_mem[4][22] ;
 wire \core.keymem.key_mem[4][23] ;
 wire \core.keymem.key_mem[4][24] ;
 wire \core.keymem.key_mem[4][25] ;
 wire \core.keymem.key_mem[4][26] ;
 wire \core.keymem.key_mem[4][27] ;
 wire \core.keymem.key_mem[4][28] ;
 wire \core.keymem.key_mem[4][29] ;
 wire \core.keymem.key_mem[4][2] ;
 wire \core.keymem.key_mem[4][30] ;
 wire \core.keymem.key_mem[4][31] ;
 wire \core.keymem.key_mem[4][32] ;
 wire \core.keymem.key_mem[4][33] ;
 wire \core.keymem.key_mem[4][34] ;
 wire \core.keymem.key_mem[4][35] ;
 wire \core.keymem.key_mem[4][36] ;
 wire \core.keymem.key_mem[4][37] ;
 wire \core.keymem.key_mem[4][38] ;
 wire \core.keymem.key_mem[4][39] ;
 wire \core.keymem.key_mem[4][3] ;
 wire \core.keymem.key_mem[4][40] ;
 wire \core.keymem.key_mem[4][41] ;
 wire \core.keymem.key_mem[4][42] ;
 wire \core.keymem.key_mem[4][43] ;
 wire \core.keymem.key_mem[4][44] ;
 wire \core.keymem.key_mem[4][45] ;
 wire \core.keymem.key_mem[4][46] ;
 wire \core.keymem.key_mem[4][47] ;
 wire \core.keymem.key_mem[4][48] ;
 wire \core.keymem.key_mem[4][49] ;
 wire \core.keymem.key_mem[4][4] ;
 wire \core.keymem.key_mem[4][50] ;
 wire \core.keymem.key_mem[4][51] ;
 wire \core.keymem.key_mem[4][52] ;
 wire \core.keymem.key_mem[4][53] ;
 wire \core.keymem.key_mem[4][54] ;
 wire \core.keymem.key_mem[4][55] ;
 wire \core.keymem.key_mem[4][56] ;
 wire \core.keymem.key_mem[4][57] ;
 wire \core.keymem.key_mem[4][58] ;
 wire \core.keymem.key_mem[4][59] ;
 wire \core.keymem.key_mem[4][5] ;
 wire \core.keymem.key_mem[4][60] ;
 wire \core.keymem.key_mem[4][61] ;
 wire \core.keymem.key_mem[4][62] ;
 wire \core.keymem.key_mem[4][63] ;
 wire \core.keymem.key_mem[4][64] ;
 wire \core.keymem.key_mem[4][65] ;
 wire \core.keymem.key_mem[4][66] ;
 wire \core.keymem.key_mem[4][67] ;
 wire \core.keymem.key_mem[4][68] ;
 wire \core.keymem.key_mem[4][69] ;
 wire \core.keymem.key_mem[4][6] ;
 wire \core.keymem.key_mem[4][70] ;
 wire \core.keymem.key_mem[4][71] ;
 wire \core.keymem.key_mem[4][72] ;
 wire \core.keymem.key_mem[4][73] ;
 wire \core.keymem.key_mem[4][74] ;
 wire \core.keymem.key_mem[4][75] ;
 wire \core.keymem.key_mem[4][76] ;
 wire \core.keymem.key_mem[4][77] ;
 wire \core.keymem.key_mem[4][78] ;
 wire \core.keymem.key_mem[4][79] ;
 wire \core.keymem.key_mem[4][7] ;
 wire \core.keymem.key_mem[4][80] ;
 wire \core.keymem.key_mem[4][81] ;
 wire \core.keymem.key_mem[4][82] ;
 wire \core.keymem.key_mem[4][83] ;
 wire \core.keymem.key_mem[4][84] ;
 wire \core.keymem.key_mem[4][85] ;
 wire \core.keymem.key_mem[4][86] ;
 wire \core.keymem.key_mem[4][87] ;
 wire \core.keymem.key_mem[4][88] ;
 wire \core.keymem.key_mem[4][89] ;
 wire \core.keymem.key_mem[4][8] ;
 wire \core.keymem.key_mem[4][90] ;
 wire \core.keymem.key_mem[4][91] ;
 wire \core.keymem.key_mem[4][92] ;
 wire \core.keymem.key_mem[4][93] ;
 wire \core.keymem.key_mem[4][94] ;
 wire \core.keymem.key_mem[4][95] ;
 wire \core.keymem.key_mem[4][96] ;
 wire \core.keymem.key_mem[4][97] ;
 wire \core.keymem.key_mem[4][98] ;
 wire \core.keymem.key_mem[4][99] ;
 wire \core.keymem.key_mem[4][9] ;
 wire \core.keymem.key_mem[5][0] ;
 wire \core.keymem.key_mem[5][100] ;
 wire \core.keymem.key_mem[5][101] ;
 wire \core.keymem.key_mem[5][102] ;
 wire \core.keymem.key_mem[5][103] ;
 wire \core.keymem.key_mem[5][104] ;
 wire \core.keymem.key_mem[5][105] ;
 wire \core.keymem.key_mem[5][106] ;
 wire \core.keymem.key_mem[5][107] ;
 wire \core.keymem.key_mem[5][108] ;
 wire \core.keymem.key_mem[5][109] ;
 wire \core.keymem.key_mem[5][10] ;
 wire \core.keymem.key_mem[5][110] ;
 wire \core.keymem.key_mem[5][111] ;
 wire \core.keymem.key_mem[5][112] ;
 wire \core.keymem.key_mem[5][113] ;
 wire \core.keymem.key_mem[5][114] ;
 wire \core.keymem.key_mem[5][115] ;
 wire \core.keymem.key_mem[5][116] ;
 wire \core.keymem.key_mem[5][117] ;
 wire \core.keymem.key_mem[5][118] ;
 wire \core.keymem.key_mem[5][119] ;
 wire \core.keymem.key_mem[5][11] ;
 wire \core.keymem.key_mem[5][120] ;
 wire \core.keymem.key_mem[5][121] ;
 wire \core.keymem.key_mem[5][122] ;
 wire \core.keymem.key_mem[5][123] ;
 wire \core.keymem.key_mem[5][124] ;
 wire \core.keymem.key_mem[5][125] ;
 wire \core.keymem.key_mem[5][126] ;
 wire \core.keymem.key_mem[5][127] ;
 wire \core.keymem.key_mem[5][12] ;
 wire \core.keymem.key_mem[5][13] ;
 wire \core.keymem.key_mem[5][14] ;
 wire \core.keymem.key_mem[5][15] ;
 wire \core.keymem.key_mem[5][16] ;
 wire \core.keymem.key_mem[5][17] ;
 wire \core.keymem.key_mem[5][18] ;
 wire \core.keymem.key_mem[5][19] ;
 wire \core.keymem.key_mem[5][1] ;
 wire \core.keymem.key_mem[5][20] ;
 wire \core.keymem.key_mem[5][21] ;
 wire \core.keymem.key_mem[5][22] ;
 wire \core.keymem.key_mem[5][23] ;
 wire \core.keymem.key_mem[5][24] ;
 wire \core.keymem.key_mem[5][25] ;
 wire \core.keymem.key_mem[5][26] ;
 wire \core.keymem.key_mem[5][27] ;
 wire \core.keymem.key_mem[5][28] ;
 wire \core.keymem.key_mem[5][29] ;
 wire \core.keymem.key_mem[5][2] ;
 wire \core.keymem.key_mem[5][30] ;
 wire \core.keymem.key_mem[5][31] ;
 wire \core.keymem.key_mem[5][32] ;
 wire \core.keymem.key_mem[5][33] ;
 wire \core.keymem.key_mem[5][34] ;
 wire \core.keymem.key_mem[5][35] ;
 wire \core.keymem.key_mem[5][36] ;
 wire \core.keymem.key_mem[5][37] ;
 wire \core.keymem.key_mem[5][38] ;
 wire \core.keymem.key_mem[5][39] ;
 wire \core.keymem.key_mem[5][3] ;
 wire \core.keymem.key_mem[5][40] ;
 wire \core.keymem.key_mem[5][41] ;
 wire \core.keymem.key_mem[5][42] ;
 wire \core.keymem.key_mem[5][43] ;
 wire \core.keymem.key_mem[5][44] ;
 wire \core.keymem.key_mem[5][45] ;
 wire \core.keymem.key_mem[5][46] ;
 wire \core.keymem.key_mem[5][47] ;
 wire \core.keymem.key_mem[5][48] ;
 wire \core.keymem.key_mem[5][49] ;
 wire \core.keymem.key_mem[5][4] ;
 wire \core.keymem.key_mem[5][50] ;
 wire \core.keymem.key_mem[5][51] ;
 wire \core.keymem.key_mem[5][52] ;
 wire \core.keymem.key_mem[5][53] ;
 wire \core.keymem.key_mem[5][54] ;
 wire \core.keymem.key_mem[5][55] ;
 wire \core.keymem.key_mem[5][56] ;
 wire \core.keymem.key_mem[5][57] ;
 wire \core.keymem.key_mem[5][58] ;
 wire \core.keymem.key_mem[5][59] ;
 wire \core.keymem.key_mem[5][5] ;
 wire \core.keymem.key_mem[5][60] ;
 wire \core.keymem.key_mem[5][61] ;
 wire \core.keymem.key_mem[5][62] ;
 wire \core.keymem.key_mem[5][63] ;
 wire \core.keymem.key_mem[5][64] ;
 wire \core.keymem.key_mem[5][65] ;
 wire \core.keymem.key_mem[5][66] ;
 wire \core.keymem.key_mem[5][67] ;
 wire \core.keymem.key_mem[5][68] ;
 wire \core.keymem.key_mem[5][69] ;
 wire \core.keymem.key_mem[5][6] ;
 wire \core.keymem.key_mem[5][70] ;
 wire \core.keymem.key_mem[5][71] ;
 wire \core.keymem.key_mem[5][72] ;
 wire \core.keymem.key_mem[5][73] ;
 wire \core.keymem.key_mem[5][74] ;
 wire \core.keymem.key_mem[5][75] ;
 wire \core.keymem.key_mem[5][76] ;
 wire \core.keymem.key_mem[5][77] ;
 wire \core.keymem.key_mem[5][78] ;
 wire \core.keymem.key_mem[5][79] ;
 wire \core.keymem.key_mem[5][7] ;
 wire \core.keymem.key_mem[5][80] ;
 wire \core.keymem.key_mem[5][81] ;
 wire \core.keymem.key_mem[5][82] ;
 wire \core.keymem.key_mem[5][83] ;
 wire \core.keymem.key_mem[5][84] ;
 wire \core.keymem.key_mem[5][85] ;
 wire \core.keymem.key_mem[5][86] ;
 wire \core.keymem.key_mem[5][87] ;
 wire \core.keymem.key_mem[5][88] ;
 wire \core.keymem.key_mem[5][89] ;
 wire \core.keymem.key_mem[5][8] ;
 wire \core.keymem.key_mem[5][90] ;
 wire \core.keymem.key_mem[5][91] ;
 wire \core.keymem.key_mem[5][92] ;
 wire \core.keymem.key_mem[5][93] ;
 wire \core.keymem.key_mem[5][94] ;
 wire \core.keymem.key_mem[5][95] ;
 wire \core.keymem.key_mem[5][96] ;
 wire \core.keymem.key_mem[5][97] ;
 wire \core.keymem.key_mem[5][98] ;
 wire \core.keymem.key_mem[5][99] ;
 wire \core.keymem.key_mem[5][9] ;
 wire \core.keymem.key_mem[6][0] ;
 wire \core.keymem.key_mem[6][100] ;
 wire \core.keymem.key_mem[6][101] ;
 wire \core.keymem.key_mem[6][102] ;
 wire \core.keymem.key_mem[6][103] ;
 wire \core.keymem.key_mem[6][104] ;
 wire \core.keymem.key_mem[6][105] ;
 wire \core.keymem.key_mem[6][106] ;
 wire \core.keymem.key_mem[6][107] ;
 wire \core.keymem.key_mem[6][108] ;
 wire \core.keymem.key_mem[6][109] ;
 wire \core.keymem.key_mem[6][10] ;
 wire \core.keymem.key_mem[6][110] ;
 wire \core.keymem.key_mem[6][111] ;
 wire \core.keymem.key_mem[6][112] ;
 wire \core.keymem.key_mem[6][113] ;
 wire \core.keymem.key_mem[6][114] ;
 wire \core.keymem.key_mem[6][115] ;
 wire \core.keymem.key_mem[6][116] ;
 wire \core.keymem.key_mem[6][117] ;
 wire \core.keymem.key_mem[6][118] ;
 wire \core.keymem.key_mem[6][119] ;
 wire \core.keymem.key_mem[6][11] ;
 wire \core.keymem.key_mem[6][120] ;
 wire \core.keymem.key_mem[6][121] ;
 wire \core.keymem.key_mem[6][122] ;
 wire \core.keymem.key_mem[6][123] ;
 wire \core.keymem.key_mem[6][124] ;
 wire \core.keymem.key_mem[6][125] ;
 wire \core.keymem.key_mem[6][126] ;
 wire \core.keymem.key_mem[6][127] ;
 wire \core.keymem.key_mem[6][12] ;
 wire \core.keymem.key_mem[6][13] ;
 wire \core.keymem.key_mem[6][14] ;
 wire \core.keymem.key_mem[6][15] ;
 wire \core.keymem.key_mem[6][16] ;
 wire \core.keymem.key_mem[6][17] ;
 wire \core.keymem.key_mem[6][18] ;
 wire \core.keymem.key_mem[6][19] ;
 wire \core.keymem.key_mem[6][1] ;
 wire \core.keymem.key_mem[6][20] ;
 wire \core.keymem.key_mem[6][21] ;
 wire \core.keymem.key_mem[6][22] ;
 wire \core.keymem.key_mem[6][23] ;
 wire \core.keymem.key_mem[6][24] ;
 wire \core.keymem.key_mem[6][25] ;
 wire \core.keymem.key_mem[6][26] ;
 wire \core.keymem.key_mem[6][27] ;
 wire \core.keymem.key_mem[6][28] ;
 wire \core.keymem.key_mem[6][29] ;
 wire \core.keymem.key_mem[6][2] ;
 wire \core.keymem.key_mem[6][30] ;
 wire \core.keymem.key_mem[6][31] ;
 wire \core.keymem.key_mem[6][32] ;
 wire \core.keymem.key_mem[6][33] ;
 wire \core.keymem.key_mem[6][34] ;
 wire \core.keymem.key_mem[6][35] ;
 wire \core.keymem.key_mem[6][36] ;
 wire \core.keymem.key_mem[6][37] ;
 wire \core.keymem.key_mem[6][38] ;
 wire \core.keymem.key_mem[6][39] ;
 wire \core.keymem.key_mem[6][3] ;
 wire \core.keymem.key_mem[6][40] ;
 wire \core.keymem.key_mem[6][41] ;
 wire \core.keymem.key_mem[6][42] ;
 wire \core.keymem.key_mem[6][43] ;
 wire \core.keymem.key_mem[6][44] ;
 wire \core.keymem.key_mem[6][45] ;
 wire \core.keymem.key_mem[6][46] ;
 wire \core.keymem.key_mem[6][47] ;
 wire \core.keymem.key_mem[6][48] ;
 wire \core.keymem.key_mem[6][49] ;
 wire \core.keymem.key_mem[6][4] ;
 wire \core.keymem.key_mem[6][50] ;
 wire \core.keymem.key_mem[6][51] ;
 wire \core.keymem.key_mem[6][52] ;
 wire \core.keymem.key_mem[6][53] ;
 wire \core.keymem.key_mem[6][54] ;
 wire \core.keymem.key_mem[6][55] ;
 wire \core.keymem.key_mem[6][56] ;
 wire \core.keymem.key_mem[6][57] ;
 wire \core.keymem.key_mem[6][58] ;
 wire \core.keymem.key_mem[6][59] ;
 wire \core.keymem.key_mem[6][5] ;
 wire \core.keymem.key_mem[6][60] ;
 wire \core.keymem.key_mem[6][61] ;
 wire \core.keymem.key_mem[6][62] ;
 wire \core.keymem.key_mem[6][63] ;
 wire \core.keymem.key_mem[6][64] ;
 wire \core.keymem.key_mem[6][65] ;
 wire \core.keymem.key_mem[6][66] ;
 wire \core.keymem.key_mem[6][67] ;
 wire \core.keymem.key_mem[6][68] ;
 wire \core.keymem.key_mem[6][69] ;
 wire \core.keymem.key_mem[6][6] ;
 wire \core.keymem.key_mem[6][70] ;
 wire \core.keymem.key_mem[6][71] ;
 wire \core.keymem.key_mem[6][72] ;
 wire \core.keymem.key_mem[6][73] ;
 wire \core.keymem.key_mem[6][74] ;
 wire \core.keymem.key_mem[6][75] ;
 wire \core.keymem.key_mem[6][76] ;
 wire \core.keymem.key_mem[6][77] ;
 wire \core.keymem.key_mem[6][78] ;
 wire \core.keymem.key_mem[6][79] ;
 wire \core.keymem.key_mem[6][7] ;
 wire \core.keymem.key_mem[6][80] ;
 wire \core.keymem.key_mem[6][81] ;
 wire \core.keymem.key_mem[6][82] ;
 wire \core.keymem.key_mem[6][83] ;
 wire \core.keymem.key_mem[6][84] ;
 wire \core.keymem.key_mem[6][85] ;
 wire \core.keymem.key_mem[6][86] ;
 wire \core.keymem.key_mem[6][87] ;
 wire \core.keymem.key_mem[6][88] ;
 wire \core.keymem.key_mem[6][89] ;
 wire \core.keymem.key_mem[6][8] ;
 wire \core.keymem.key_mem[6][90] ;
 wire \core.keymem.key_mem[6][91] ;
 wire \core.keymem.key_mem[6][92] ;
 wire \core.keymem.key_mem[6][93] ;
 wire \core.keymem.key_mem[6][94] ;
 wire \core.keymem.key_mem[6][95] ;
 wire \core.keymem.key_mem[6][96] ;
 wire \core.keymem.key_mem[6][97] ;
 wire \core.keymem.key_mem[6][98] ;
 wire \core.keymem.key_mem[6][99] ;
 wire \core.keymem.key_mem[6][9] ;
 wire \core.keymem.key_mem[7][0] ;
 wire \core.keymem.key_mem[7][100] ;
 wire \core.keymem.key_mem[7][101] ;
 wire \core.keymem.key_mem[7][102] ;
 wire \core.keymem.key_mem[7][103] ;
 wire \core.keymem.key_mem[7][104] ;
 wire \core.keymem.key_mem[7][105] ;
 wire \core.keymem.key_mem[7][106] ;
 wire \core.keymem.key_mem[7][107] ;
 wire \core.keymem.key_mem[7][108] ;
 wire \core.keymem.key_mem[7][109] ;
 wire \core.keymem.key_mem[7][10] ;
 wire \core.keymem.key_mem[7][110] ;
 wire \core.keymem.key_mem[7][111] ;
 wire \core.keymem.key_mem[7][112] ;
 wire \core.keymem.key_mem[7][113] ;
 wire \core.keymem.key_mem[7][114] ;
 wire \core.keymem.key_mem[7][115] ;
 wire \core.keymem.key_mem[7][116] ;
 wire \core.keymem.key_mem[7][117] ;
 wire \core.keymem.key_mem[7][118] ;
 wire \core.keymem.key_mem[7][119] ;
 wire \core.keymem.key_mem[7][11] ;
 wire \core.keymem.key_mem[7][120] ;
 wire \core.keymem.key_mem[7][121] ;
 wire \core.keymem.key_mem[7][122] ;
 wire \core.keymem.key_mem[7][123] ;
 wire \core.keymem.key_mem[7][124] ;
 wire \core.keymem.key_mem[7][125] ;
 wire \core.keymem.key_mem[7][126] ;
 wire \core.keymem.key_mem[7][127] ;
 wire \core.keymem.key_mem[7][12] ;
 wire \core.keymem.key_mem[7][13] ;
 wire \core.keymem.key_mem[7][14] ;
 wire \core.keymem.key_mem[7][15] ;
 wire \core.keymem.key_mem[7][16] ;
 wire \core.keymem.key_mem[7][17] ;
 wire \core.keymem.key_mem[7][18] ;
 wire \core.keymem.key_mem[7][19] ;
 wire \core.keymem.key_mem[7][1] ;
 wire \core.keymem.key_mem[7][20] ;
 wire \core.keymem.key_mem[7][21] ;
 wire \core.keymem.key_mem[7][22] ;
 wire \core.keymem.key_mem[7][23] ;
 wire \core.keymem.key_mem[7][24] ;
 wire \core.keymem.key_mem[7][25] ;
 wire \core.keymem.key_mem[7][26] ;
 wire \core.keymem.key_mem[7][27] ;
 wire \core.keymem.key_mem[7][28] ;
 wire \core.keymem.key_mem[7][29] ;
 wire \core.keymem.key_mem[7][2] ;
 wire \core.keymem.key_mem[7][30] ;
 wire \core.keymem.key_mem[7][31] ;
 wire \core.keymem.key_mem[7][32] ;
 wire \core.keymem.key_mem[7][33] ;
 wire \core.keymem.key_mem[7][34] ;
 wire \core.keymem.key_mem[7][35] ;
 wire \core.keymem.key_mem[7][36] ;
 wire \core.keymem.key_mem[7][37] ;
 wire \core.keymem.key_mem[7][38] ;
 wire \core.keymem.key_mem[7][39] ;
 wire \core.keymem.key_mem[7][3] ;
 wire \core.keymem.key_mem[7][40] ;
 wire \core.keymem.key_mem[7][41] ;
 wire \core.keymem.key_mem[7][42] ;
 wire \core.keymem.key_mem[7][43] ;
 wire \core.keymem.key_mem[7][44] ;
 wire \core.keymem.key_mem[7][45] ;
 wire \core.keymem.key_mem[7][46] ;
 wire \core.keymem.key_mem[7][47] ;
 wire \core.keymem.key_mem[7][48] ;
 wire \core.keymem.key_mem[7][49] ;
 wire \core.keymem.key_mem[7][4] ;
 wire \core.keymem.key_mem[7][50] ;
 wire \core.keymem.key_mem[7][51] ;
 wire \core.keymem.key_mem[7][52] ;
 wire \core.keymem.key_mem[7][53] ;
 wire \core.keymem.key_mem[7][54] ;
 wire \core.keymem.key_mem[7][55] ;
 wire \core.keymem.key_mem[7][56] ;
 wire \core.keymem.key_mem[7][57] ;
 wire \core.keymem.key_mem[7][58] ;
 wire \core.keymem.key_mem[7][59] ;
 wire \core.keymem.key_mem[7][5] ;
 wire \core.keymem.key_mem[7][60] ;
 wire \core.keymem.key_mem[7][61] ;
 wire \core.keymem.key_mem[7][62] ;
 wire \core.keymem.key_mem[7][63] ;
 wire \core.keymem.key_mem[7][64] ;
 wire \core.keymem.key_mem[7][65] ;
 wire \core.keymem.key_mem[7][66] ;
 wire \core.keymem.key_mem[7][67] ;
 wire \core.keymem.key_mem[7][68] ;
 wire \core.keymem.key_mem[7][69] ;
 wire \core.keymem.key_mem[7][6] ;
 wire \core.keymem.key_mem[7][70] ;
 wire \core.keymem.key_mem[7][71] ;
 wire \core.keymem.key_mem[7][72] ;
 wire \core.keymem.key_mem[7][73] ;
 wire \core.keymem.key_mem[7][74] ;
 wire \core.keymem.key_mem[7][75] ;
 wire \core.keymem.key_mem[7][76] ;
 wire \core.keymem.key_mem[7][77] ;
 wire \core.keymem.key_mem[7][78] ;
 wire \core.keymem.key_mem[7][79] ;
 wire \core.keymem.key_mem[7][7] ;
 wire \core.keymem.key_mem[7][80] ;
 wire \core.keymem.key_mem[7][81] ;
 wire \core.keymem.key_mem[7][82] ;
 wire \core.keymem.key_mem[7][83] ;
 wire \core.keymem.key_mem[7][84] ;
 wire \core.keymem.key_mem[7][85] ;
 wire \core.keymem.key_mem[7][86] ;
 wire \core.keymem.key_mem[7][87] ;
 wire \core.keymem.key_mem[7][88] ;
 wire \core.keymem.key_mem[7][89] ;
 wire \core.keymem.key_mem[7][8] ;
 wire \core.keymem.key_mem[7][90] ;
 wire \core.keymem.key_mem[7][91] ;
 wire \core.keymem.key_mem[7][92] ;
 wire \core.keymem.key_mem[7][93] ;
 wire \core.keymem.key_mem[7][94] ;
 wire \core.keymem.key_mem[7][95] ;
 wire \core.keymem.key_mem[7][96] ;
 wire \core.keymem.key_mem[7][97] ;
 wire \core.keymem.key_mem[7][98] ;
 wire \core.keymem.key_mem[7][99] ;
 wire \core.keymem.key_mem[7][9] ;
 wire \core.keymem.key_mem[8][0] ;
 wire \core.keymem.key_mem[8][100] ;
 wire \core.keymem.key_mem[8][101] ;
 wire \core.keymem.key_mem[8][102] ;
 wire \core.keymem.key_mem[8][103] ;
 wire \core.keymem.key_mem[8][104] ;
 wire \core.keymem.key_mem[8][105] ;
 wire \core.keymem.key_mem[8][106] ;
 wire \core.keymem.key_mem[8][107] ;
 wire \core.keymem.key_mem[8][108] ;
 wire \core.keymem.key_mem[8][109] ;
 wire \core.keymem.key_mem[8][10] ;
 wire \core.keymem.key_mem[8][110] ;
 wire \core.keymem.key_mem[8][111] ;
 wire \core.keymem.key_mem[8][112] ;
 wire \core.keymem.key_mem[8][113] ;
 wire \core.keymem.key_mem[8][114] ;
 wire \core.keymem.key_mem[8][115] ;
 wire \core.keymem.key_mem[8][116] ;
 wire \core.keymem.key_mem[8][117] ;
 wire \core.keymem.key_mem[8][118] ;
 wire \core.keymem.key_mem[8][119] ;
 wire \core.keymem.key_mem[8][11] ;
 wire \core.keymem.key_mem[8][120] ;
 wire \core.keymem.key_mem[8][121] ;
 wire \core.keymem.key_mem[8][122] ;
 wire \core.keymem.key_mem[8][123] ;
 wire \core.keymem.key_mem[8][124] ;
 wire \core.keymem.key_mem[8][125] ;
 wire \core.keymem.key_mem[8][126] ;
 wire \core.keymem.key_mem[8][127] ;
 wire \core.keymem.key_mem[8][12] ;
 wire \core.keymem.key_mem[8][13] ;
 wire \core.keymem.key_mem[8][14] ;
 wire \core.keymem.key_mem[8][15] ;
 wire \core.keymem.key_mem[8][16] ;
 wire \core.keymem.key_mem[8][17] ;
 wire \core.keymem.key_mem[8][18] ;
 wire \core.keymem.key_mem[8][19] ;
 wire \core.keymem.key_mem[8][1] ;
 wire \core.keymem.key_mem[8][20] ;
 wire \core.keymem.key_mem[8][21] ;
 wire \core.keymem.key_mem[8][22] ;
 wire \core.keymem.key_mem[8][23] ;
 wire \core.keymem.key_mem[8][24] ;
 wire \core.keymem.key_mem[8][25] ;
 wire \core.keymem.key_mem[8][26] ;
 wire \core.keymem.key_mem[8][27] ;
 wire \core.keymem.key_mem[8][28] ;
 wire \core.keymem.key_mem[8][29] ;
 wire \core.keymem.key_mem[8][2] ;
 wire \core.keymem.key_mem[8][30] ;
 wire \core.keymem.key_mem[8][31] ;
 wire \core.keymem.key_mem[8][32] ;
 wire \core.keymem.key_mem[8][33] ;
 wire \core.keymem.key_mem[8][34] ;
 wire \core.keymem.key_mem[8][35] ;
 wire \core.keymem.key_mem[8][36] ;
 wire \core.keymem.key_mem[8][37] ;
 wire \core.keymem.key_mem[8][38] ;
 wire \core.keymem.key_mem[8][39] ;
 wire \core.keymem.key_mem[8][3] ;
 wire \core.keymem.key_mem[8][40] ;
 wire \core.keymem.key_mem[8][41] ;
 wire \core.keymem.key_mem[8][42] ;
 wire \core.keymem.key_mem[8][43] ;
 wire \core.keymem.key_mem[8][44] ;
 wire \core.keymem.key_mem[8][45] ;
 wire \core.keymem.key_mem[8][46] ;
 wire \core.keymem.key_mem[8][47] ;
 wire \core.keymem.key_mem[8][48] ;
 wire \core.keymem.key_mem[8][49] ;
 wire \core.keymem.key_mem[8][4] ;
 wire \core.keymem.key_mem[8][50] ;
 wire \core.keymem.key_mem[8][51] ;
 wire \core.keymem.key_mem[8][52] ;
 wire \core.keymem.key_mem[8][53] ;
 wire \core.keymem.key_mem[8][54] ;
 wire \core.keymem.key_mem[8][55] ;
 wire \core.keymem.key_mem[8][56] ;
 wire \core.keymem.key_mem[8][57] ;
 wire \core.keymem.key_mem[8][58] ;
 wire \core.keymem.key_mem[8][59] ;
 wire \core.keymem.key_mem[8][5] ;
 wire \core.keymem.key_mem[8][60] ;
 wire \core.keymem.key_mem[8][61] ;
 wire \core.keymem.key_mem[8][62] ;
 wire \core.keymem.key_mem[8][63] ;
 wire \core.keymem.key_mem[8][64] ;
 wire \core.keymem.key_mem[8][65] ;
 wire \core.keymem.key_mem[8][66] ;
 wire \core.keymem.key_mem[8][67] ;
 wire \core.keymem.key_mem[8][68] ;
 wire \core.keymem.key_mem[8][69] ;
 wire \core.keymem.key_mem[8][6] ;
 wire \core.keymem.key_mem[8][70] ;
 wire \core.keymem.key_mem[8][71] ;
 wire \core.keymem.key_mem[8][72] ;
 wire \core.keymem.key_mem[8][73] ;
 wire \core.keymem.key_mem[8][74] ;
 wire \core.keymem.key_mem[8][75] ;
 wire \core.keymem.key_mem[8][76] ;
 wire \core.keymem.key_mem[8][77] ;
 wire \core.keymem.key_mem[8][78] ;
 wire \core.keymem.key_mem[8][79] ;
 wire \core.keymem.key_mem[8][7] ;
 wire \core.keymem.key_mem[8][80] ;
 wire \core.keymem.key_mem[8][81] ;
 wire \core.keymem.key_mem[8][82] ;
 wire \core.keymem.key_mem[8][83] ;
 wire \core.keymem.key_mem[8][84] ;
 wire \core.keymem.key_mem[8][85] ;
 wire \core.keymem.key_mem[8][86] ;
 wire \core.keymem.key_mem[8][87] ;
 wire \core.keymem.key_mem[8][88] ;
 wire \core.keymem.key_mem[8][89] ;
 wire \core.keymem.key_mem[8][8] ;
 wire \core.keymem.key_mem[8][90] ;
 wire \core.keymem.key_mem[8][91] ;
 wire \core.keymem.key_mem[8][92] ;
 wire \core.keymem.key_mem[8][93] ;
 wire \core.keymem.key_mem[8][94] ;
 wire \core.keymem.key_mem[8][95] ;
 wire \core.keymem.key_mem[8][96] ;
 wire \core.keymem.key_mem[8][97] ;
 wire \core.keymem.key_mem[8][98] ;
 wire \core.keymem.key_mem[8][99] ;
 wire \core.keymem.key_mem[8][9] ;
 wire \core.keymem.key_mem[9][0] ;
 wire \core.keymem.key_mem[9][100] ;
 wire \core.keymem.key_mem[9][101] ;
 wire \core.keymem.key_mem[9][102] ;
 wire \core.keymem.key_mem[9][103] ;
 wire \core.keymem.key_mem[9][104] ;
 wire \core.keymem.key_mem[9][105] ;
 wire \core.keymem.key_mem[9][106] ;
 wire \core.keymem.key_mem[9][107] ;
 wire \core.keymem.key_mem[9][108] ;
 wire \core.keymem.key_mem[9][109] ;
 wire \core.keymem.key_mem[9][10] ;
 wire \core.keymem.key_mem[9][110] ;
 wire \core.keymem.key_mem[9][111] ;
 wire \core.keymem.key_mem[9][112] ;
 wire \core.keymem.key_mem[9][113] ;
 wire \core.keymem.key_mem[9][114] ;
 wire \core.keymem.key_mem[9][115] ;
 wire \core.keymem.key_mem[9][116] ;
 wire \core.keymem.key_mem[9][117] ;
 wire \core.keymem.key_mem[9][118] ;
 wire \core.keymem.key_mem[9][119] ;
 wire \core.keymem.key_mem[9][11] ;
 wire \core.keymem.key_mem[9][120] ;
 wire \core.keymem.key_mem[9][121] ;
 wire \core.keymem.key_mem[9][122] ;
 wire \core.keymem.key_mem[9][123] ;
 wire \core.keymem.key_mem[9][124] ;
 wire \core.keymem.key_mem[9][125] ;
 wire \core.keymem.key_mem[9][126] ;
 wire \core.keymem.key_mem[9][127] ;
 wire \core.keymem.key_mem[9][12] ;
 wire \core.keymem.key_mem[9][13] ;
 wire \core.keymem.key_mem[9][14] ;
 wire \core.keymem.key_mem[9][15] ;
 wire \core.keymem.key_mem[9][16] ;
 wire \core.keymem.key_mem[9][17] ;
 wire \core.keymem.key_mem[9][18] ;
 wire \core.keymem.key_mem[9][19] ;
 wire \core.keymem.key_mem[9][1] ;
 wire \core.keymem.key_mem[9][20] ;
 wire \core.keymem.key_mem[9][21] ;
 wire \core.keymem.key_mem[9][22] ;
 wire \core.keymem.key_mem[9][23] ;
 wire \core.keymem.key_mem[9][24] ;
 wire \core.keymem.key_mem[9][25] ;
 wire \core.keymem.key_mem[9][26] ;
 wire \core.keymem.key_mem[9][27] ;
 wire \core.keymem.key_mem[9][28] ;
 wire \core.keymem.key_mem[9][29] ;
 wire \core.keymem.key_mem[9][2] ;
 wire \core.keymem.key_mem[9][30] ;
 wire \core.keymem.key_mem[9][31] ;
 wire \core.keymem.key_mem[9][32] ;
 wire \core.keymem.key_mem[9][33] ;
 wire \core.keymem.key_mem[9][34] ;
 wire \core.keymem.key_mem[9][35] ;
 wire \core.keymem.key_mem[9][36] ;
 wire \core.keymem.key_mem[9][37] ;
 wire \core.keymem.key_mem[9][38] ;
 wire \core.keymem.key_mem[9][39] ;
 wire \core.keymem.key_mem[9][3] ;
 wire \core.keymem.key_mem[9][40] ;
 wire \core.keymem.key_mem[9][41] ;
 wire \core.keymem.key_mem[9][42] ;
 wire \core.keymem.key_mem[9][43] ;
 wire \core.keymem.key_mem[9][44] ;
 wire \core.keymem.key_mem[9][45] ;
 wire \core.keymem.key_mem[9][46] ;
 wire \core.keymem.key_mem[9][47] ;
 wire \core.keymem.key_mem[9][48] ;
 wire \core.keymem.key_mem[9][49] ;
 wire \core.keymem.key_mem[9][4] ;
 wire \core.keymem.key_mem[9][50] ;
 wire \core.keymem.key_mem[9][51] ;
 wire \core.keymem.key_mem[9][52] ;
 wire \core.keymem.key_mem[9][53] ;
 wire \core.keymem.key_mem[9][54] ;
 wire \core.keymem.key_mem[9][55] ;
 wire \core.keymem.key_mem[9][56] ;
 wire \core.keymem.key_mem[9][57] ;
 wire \core.keymem.key_mem[9][58] ;
 wire \core.keymem.key_mem[9][59] ;
 wire \core.keymem.key_mem[9][5] ;
 wire \core.keymem.key_mem[9][60] ;
 wire \core.keymem.key_mem[9][61] ;
 wire \core.keymem.key_mem[9][62] ;
 wire \core.keymem.key_mem[9][63] ;
 wire \core.keymem.key_mem[9][64] ;
 wire \core.keymem.key_mem[9][65] ;
 wire \core.keymem.key_mem[9][66] ;
 wire \core.keymem.key_mem[9][67] ;
 wire \core.keymem.key_mem[9][68] ;
 wire \core.keymem.key_mem[9][69] ;
 wire \core.keymem.key_mem[9][6] ;
 wire \core.keymem.key_mem[9][70] ;
 wire \core.keymem.key_mem[9][71] ;
 wire \core.keymem.key_mem[9][72] ;
 wire \core.keymem.key_mem[9][73] ;
 wire \core.keymem.key_mem[9][74] ;
 wire \core.keymem.key_mem[9][75] ;
 wire \core.keymem.key_mem[9][76] ;
 wire \core.keymem.key_mem[9][77] ;
 wire \core.keymem.key_mem[9][78] ;
 wire \core.keymem.key_mem[9][79] ;
 wire \core.keymem.key_mem[9][7] ;
 wire \core.keymem.key_mem[9][80] ;
 wire \core.keymem.key_mem[9][81] ;
 wire \core.keymem.key_mem[9][82] ;
 wire \core.keymem.key_mem[9][83] ;
 wire \core.keymem.key_mem[9][84] ;
 wire \core.keymem.key_mem[9][85] ;
 wire \core.keymem.key_mem[9][86] ;
 wire \core.keymem.key_mem[9][87] ;
 wire \core.keymem.key_mem[9][88] ;
 wire \core.keymem.key_mem[9][89] ;
 wire \core.keymem.key_mem[9][8] ;
 wire \core.keymem.key_mem[9][90] ;
 wire \core.keymem.key_mem[9][91] ;
 wire \core.keymem.key_mem[9][92] ;
 wire \core.keymem.key_mem[9][93] ;
 wire \core.keymem.key_mem[9][94] ;
 wire \core.keymem.key_mem[9][95] ;
 wire \core.keymem.key_mem[9][96] ;
 wire \core.keymem.key_mem[9][97] ;
 wire \core.keymem.key_mem[9][98] ;
 wire \core.keymem.key_mem[9][99] ;
 wire \core.keymem.key_mem[9][9] ;
 wire \core.keymem.key_mem_ctrl_reg[0] ;
 wire \core.keymem.key_mem_ctrl_reg[1] ;
 wire \core.keymem.key_mem_ctrl_reg[2] ;
 wire \core.keymem.key_mem_ctrl_reg[3] ;
 wire \core.keymem.prev_key0_reg[0] ;
 wire \core.keymem.prev_key0_reg[100] ;
 wire \core.keymem.prev_key0_reg[101] ;
 wire \core.keymem.prev_key0_reg[102] ;
 wire \core.keymem.prev_key0_reg[103] ;
 wire \core.keymem.prev_key0_reg[104] ;
 wire \core.keymem.prev_key0_reg[105] ;
 wire \core.keymem.prev_key0_reg[106] ;
 wire \core.keymem.prev_key0_reg[107] ;
 wire \core.keymem.prev_key0_reg[108] ;
 wire \core.keymem.prev_key0_reg[109] ;
 wire \core.keymem.prev_key0_reg[10] ;
 wire \core.keymem.prev_key0_reg[110] ;
 wire \core.keymem.prev_key0_reg[111] ;
 wire \core.keymem.prev_key0_reg[112] ;
 wire \core.keymem.prev_key0_reg[113] ;
 wire \core.keymem.prev_key0_reg[114] ;
 wire \core.keymem.prev_key0_reg[115] ;
 wire \core.keymem.prev_key0_reg[116] ;
 wire \core.keymem.prev_key0_reg[117] ;
 wire \core.keymem.prev_key0_reg[118] ;
 wire \core.keymem.prev_key0_reg[119] ;
 wire \core.keymem.prev_key0_reg[11] ;
 wire \core.keymem.prev_key0_reg[120] ;
 wire \core.keymem.prev_key0_reg[121] ;
 wire \core.keymem.prev_key0_reg[122] ;
 wire \core.keymem.prev_key0_reg[123] ;
 wire \core.keymem.prev_key0_reg[124] ;
 wire \core.keymem.prev_key0_reg[125] ;
 wire \core.keymem.prev_key0_reg[126] ;
 wire \core.keymem.prev_key0_reg[127] ;
 wire \core.keymem.prev_key0_reg[12] ;
 wire \core.keymem.prev_key0_reg[13] ;
 wire \core.keymem.prev_key0_reg[14] ;
 wire \core.keymem.prev_key0_reg[15] ;
 wire \core.keymem.prev_key0_reg[16] ;
 wire \core.keymem.prev_key0_reg[17] ;
 wire \core.keymem.prev_key0_reg[18] ;
 wire \core.keymem.prev_key0_reg[19] ;
 wire \core.keymem.prev_key0_reg[1] ;
 wire \core.keymem.prev_key0_reg[20] ;
 wire \core.keymem.prev_key0_reg[21] ;
 wire \core.keymem.prev_key0_reg[22] ;
 wire \core.keymem.prev_key0_reg[23] ;
 wire \core.keymem.prev_key0_reg[24] ;
 wire \core.keymem.prev_key0_reg[25] ;
 wire \core.keymem.prev_key0_reg[26] ;
 wire \core.keymem.prev_key0_reg[27] ;
 wire \core.keymem.prev_key0_reg[28] ;
 wire \core.keymem.prev_key0_reg[29] ;
 wire \core.keymem.prev_key0_reg[2] ;
 wire \core.keymem.prev_key0_reg[30] ;
 wire \core.keymem.prev_key0_reg[31] ;
 wire \core.keymem.prev_key0_reg[32] ;
 wire \core.keymem.prev_key0_reg[33] ;
 wire \core.keymem.prev_key0_reg[34] ;
 wire \core.keymem.prev_key0_reg[35] ;
 wire \core.keymem.prev_key0_reg[36] ;
 wire \core.keymem.prev_key0_reg[37] ;
 wire \core.keymem.prev_key0_reg[38] ;
 wire \core.keymem.prev_key0_reg[39] ;
 wire \core.keymem.prev_key0_reg[3] ;
 wire \core.keymem.prev_key0_reg[40] ;
 wire \core.keymem.prev_key0_reg[41] ;
 wire \core.keymem.prev_key0_reg[42] ;
 wire \core.keymem.prev_key0_reg[43] ;
 wire \core.keymem.prev_key0_reg[44] ;
 wire \core.keymem.prev_key0_reg[45] ;
 wire \core.keymem.prev_key0_reg[46] ;
 wire \core.keymem.prev_key0_reg[47] ;
 wire \core.keymem.prev_key0_reg[48] ;
 wire \core.keymem.prev_key0_reg[49] ;
 wire \core.keymem.prev_key0_reg[4] ;
 wire \core.keymem.prev_key0_reg[50] ;
 wire \core.keymem.prev_key0_reg[51] ;
 wire \core.keymem.prev_key0_reg[52] ;
 wire \core.keymem.prev_key0_reg[53] ;
 wire \core.keymem.prev_key0_reg[54] ;
 wire \core.keymem.prev_key0_reg[55] ;
 wire \core.keymem.prev_key0_reg[56] ;
 wire \core.keymem.prev_key0_reg[57] ;
 wire \core.keymem.prev_key0_reg[58] ;
 wire \core.keymem.prev_key0_reg[59] ;
 wire \core.keymem.prev_key0_reg[5] ;
 wire \core.keymem.prev_key0_reg[60] ;
 wire \core.keymem.prev_key0_reg[61] ;
 wire \core.keymem.prev_key0_reg[62] ;
 wire \core.keymem.prev_key0_reg[63] ;
 wire \core.keymem.prev_key0_reg[64] ;
 wire \core.keymem.prev_key0_reg[65] ;
 wire \core.keymem.prev_key0_reg[66] ;
 wire \core.keymem.prev_key0_reg[67] ;
 wire \core.keymem.prev_key0_reg[68] ;
 wire \core.keymem.prev_key0_reg[69] ;
 wire \core.keymem.prev_key0_reg[6] ;
 wire \core.keymem.prev_key0_reg[70] ;
 wire \core.keymem.prev_key0_reg[71] ;
 wire \core.keymem.prev_key0_reg[72] ;
 wire \core.keymem.prev_key0_reg[73] ;
 wire \core.keymem.prev_key0_reg[74] ;
 wire \core.keymem.prev_key0_reg[75] ;
 wire \core.keymem.prev_key0_reg[76] ;
 wire \core.keymem.prev_key0_reg[77] ;
 wire \core.keymem.prev_key0_reg[78] ;
 wire \core.keymem.prev_key0_reg[79] ;
 wire \core.keymem.prev_key0_reg[7] ;
 wire \core.keymem.prev_key0_reg[80] ;
 wire \core.keymem.prev_key0_reg[81] ;
 wire \core.keymem.prev_key0_reg[82] ;
 wire \core.keymem.prev_key0_reg[83] ;
 wire \core.keymem.prev_key0_reg[84] ;
 wire \core.keymem.prev_key0_reg[85] ;
 wire \core.keymem.prev_key0_reg[86] ;
 wire \core.keymem.prev_key0_reg[87] ;
 wire \core.keymem.prev_key0_reg[88] ;
 wire \core.keymem.prev_key0_reg[89] ;
 wire \core.keymem.prev_key0_reg[8] ;
 wire \core.keymem.prev_key0_reg[90] ;
 wire \core.keymem.prev_key0_reg[91] ;
 wire \core.keymem.prev_key0_reg[92] ;
 wire \core.keymem.prev_key0_reg[93] ;
 wire \core.keymem.prev_key0_reg[94] ;
 wire \core.keymem.prev_key0_reg[95] ;
 wire \core.keymem.prev_key0_reg[96] ;
 wire \core.keymem.prev_key0_reg[97] ;
 wire \core.keymem.prev_key0_reg[98] ;
 wire \core.keymem.prev_key0_reg[99] ;
 wire \core.keymem.prev_key0_reg[9] ;
 wire \core.keymem.prev_key1_reg[0] ;
 wire \core.keymem.prev_key1_reg[100] ;
 wire \core.keymem.prev_key1_reg[101] ;
 wire \core.keymem.prev_key1_reg[102] ;
 wire \core.keymem.prev_key1_reg[103] ;
 wire \core.keymem.prev_key1_reg[104] ;
 wire \core.keymem.prev_key1_reg[105] ;
 wire \core.keymem.prev_key1_reg[106] ;
 wire \core.keymem.prev_key1_reg[107] ;
 wire \core.keymem.prev_key1_reg[108] ;
 wire \core.keymem.prev_key1_reg[109] ;
 wire \core.keymem.prev_key1_reg[10] ;
 wire \core.keymem.prev_key1_reg[110] ;
 wire \core.keymem.prev_key1_reg[111] ;
 wire \core.keymem.prev_key1_reg[112] ;
 wire \core.keymem.prev_key1_reg[113] ;
 wire \core.keymem.prev_key1_reg[114] ;
 wire \core.keymem.prev_key1_reg[115] ;
 wire \core.keymem.prev_key1_reg[116] ;
 wire \core.keymem.prev_key1_reg[117] ;
 wire \core.keymem.prev_key1_reg[118] ;
 wire \core.keymem.prev_key1_reg[119] ;
 wire \core.keymem.prev_key1_reg[11] ;
 wire \core.keymem.prev_key1_reg[120] ;
 wire \core.keymem.prev_key1_reg[121] ;
 wire \core.keymem.prev_key1_reg[122] ;
 wire \core.keymem.prev_key1_reg[123] ;
 wire \core.keymem.prev_key1_reg[124] ;
 wire \core.keymem.prev_key1_reg[125] ;
 wire \core.keymem.prev_key1_reg[126] ;
 wire \core.keymem.prev_key1_reg[127] ;
 wire \core.keymem.prev_key1_reg[12] ;
 wire \core.keymem.prev_key1_reg[13] ;
 wire \core.keymem.prev_key1_reg[14] ;
 wire \core.keymem.prev_key1_reg[15] ;
 wire \core.keymem.prev_key1_reg[16] ;
 wire \core.keymem.prev_key1_reg[17] ;
 wire \core.keymem.prev_key1_reg[18] ;
 wire \core.keymem.prev_key1_reg[19] ;
 wire \core.keymem.prev_key1_reg[1] ;
 wire \core.keymem.prev_key1_reg[20] ;
 wire \core.keymem.prev_key1_reg[21] ;
 wire \core.keymem.prev_key1_reg[22] ;
 wire \core.keymem.prev_key1_reg[23] ;
 wire \core.keymem.prev_key1_reg[24] ;
 wire \core.keymem.prev_key1_reg[25] ;
 wire \core.keymem.prev_key1_reg[26] ;
 wire \core.keymem.prev_key1_reg[27] ;
 wire \core.keymem.prev_key1_reg[28] ;
 wire \core.keymem.prev_key1_reg[29] ;
 wire \core.keymem.prev_key1_reg[2] ;
 wire \core.keymem.prev_key1_reg[30] ;
 wire \core.keymem.prev_key1_reg[31] ;
 wire \core.keymem.prev_key1_reg[32] ;
 wire \core.keymem.prev_key1_reg[33] ;
 wire \core.keymem.prev_key1_reg[34] ;
 wire \core.keymem.prev_key1_reg[35] ;
 wire \core.keymem.prev_key1_reg[36] ;
 wire \core.keymem.prev_key1_reg[37] ;
 wire \core.keymem.prev_key1_reg[38] ;
 wire \core.keymem.prev_key1_reg[39] ;
 wire \core.keymem.prev_key1_reg[3] ;
 wire \core.keymem.prev_key1_reg[40] ;
 wire \core.keymem.prev_key1_reg[41] ;
 wire \core.keymem.prev_key1_reg[42] ;
 wire \core.keymem.prev_key1_reg[43] ;
 wire \core.keymem.prev_key1_reg[44] ;
 wire \core.keymem.prev_key1_reg[45] ;
 wire \core.keymem.prev_key1_reg[46] ;
 wire \core.keymem.prev_key1_reg[47] ;
 wire \core.keymem.prev_key1_reg[48] ;
 wire \core.keymem.prev_key1_reg[49] ;
 wire \core.keymem.prev_key1_reg[4] ;
 wire \core.keymem.prev_key1_reg[50] ;
 wire \core.keymem.prev_key1_reg[51] ;
 wire \core.keymem.prev_key1_reg[52] ;
 wire \core.keymem.prev_key1_reg[53] ;
 wire \core.keymem.prev_key1_reg[54] ;
 wire \core.keymem.prev_key1_reg[55] ;
 wire \core.keymem.prev_key1_reg[56] ;
 wire \core.keymem.prev_key1_reg[57] ;
 wire \core.keymem.prev_key1_reg[58] ;
 wire \core.keymem.prev_key1_reg[59] ;
 wire \core.keymem.prev_key1_reg[5] ;
 wire \core.keymem.prev_key1_reg[60] ;
 wire \core.keymem.prev_key1_reg[61] ;
 wire \core.keymem.prev_key1_reg[62] ;
 wire \core.keymem.prev_key1_reg[63] ;
 wire \core.keymem.prev_key1_reg[64] ;
 wire \core.keymem.prev_key1_reg[65] ;
 wire \core.keymem.prev_key1_reg[66] ;
 wire \core.keymem.prev_key1_reg[67] ;
 wire \core.keymem.prev_key1_reg[68] ;
 wire \core.keymem.prev_key1_reg[69] ;
 wire \core.keymem.prev_key1_reg[6] ;
 wire \core.keymem.prev_key1_reg[70] ;
 wire \core.keymem.prev_key1_reg[71] ;
 wire \core.keymem.prev_key1_reg[72] ;
 wire \core.keymem.prev_key1_reg[73] ;
 wire \core.keymem.prev_key1_reg[74] ;
 wire \core.keymem.prev_key1_reg[75] ;
 wire \core.keymem.prev_key1_reg[76] ;
 wire \core.keymem.prev_key1_reg[77] ;
 wire \core.keymem.prev_key1_reg[78] ;
 wire \core.keymem.prev_key1_reg[79] ;
 wire \core.keymem.prev_key1_reg[7] ;
 wire \core.keymem.prev_key1_reg[80] ;
 wire \core.keymem.prev_key1_reg[81] ;
 wire \core.keymem.prev_key1_reg[82] ;
 wire \core.keymem.prev_key1_reg[83] ;
 wire \core.keymem.prev_key1_reg[84] ;
 wire \core.keymem.prev_key1_reg[85] ;
 wire \core.keymem.prev_key1_reg[86] ;
 wire \core.keymem.prev_key1_reg[87] ;
 wire \core.keymem.prev_key1_reg[88] ;
 wire \core.keymem.prev_key1_reg[89] ;
 wire \core.keymem.prev_key1_reg[8] ;
 wire \core.keymem.prev_key1_reg[90] ;
 wire \core.keymem.prev_key1_reg[91] ;
 wire \core.keymem.prev_key1_reg[92] ;
 wire \core.keymem.prev_key1_reg[93] ;
 wire \core.keymem.prev_key1_reg[94] ;
 wire \core.keymem.prev_key1_reg[95] ;
 wire \core.keymem.prev_key1_reg[96] ;
 wire \core.keymem.prev_key1_reg[97] ;
 wire \core.keymem.prev_key1_reg[98] ;
 wire \core.keymem.prev_key1_reg[99] ;
 wire \core.keymem.prev_key1_reg[9] ;
 wire \core.keymem.rcon_logic.tmp_rcon[0] ;
 wire \core.keymem.rcon_logic.tmp_rcon[2] ;
 wire \core.keymem.rcon_logic.tmp_rcon[5] ;
 wire \core.keymem.rcon_logic.tmp_rcon[6] ;
 wire \core.keymem.rcon_logic.tmp_rcon[7] ;
 wire \core.keymem.rcon_reg[0] ;
 wire \core.keymem.rcon_reg[2] ;
 wire \core.keymem.rcon_reg[3] ;
 wire \core.keymem.round_ctr_reg[0] ;
 wire \core.keymem.round_ctr_reg[1] ;
 wire \core.keymem.round_ctr_reg[2] ;
 wire \core.keymem.round_ctr_reg[3] ;
 wire \core.muxed_new_block[0] ;
 wire \core.muxed_new_block[100] ;
 wire \core.muxed_new_block[101] ;
 wire \core.muxed_new_block[102] ;
 wire \core.muxed_new_block[103] ;
 wire \core.muxed_new_block[104] ;
 wire \core.muxed_new_block[105] ;
 wire \core.muxed_new_block[106] ;
 wire \core.muxed_new_block[107] ;
 wire \core.muxed_new_block[108] ;
 wire \core.muxed_new_block[109] ;
 wire \core.muxed_new_block[10] ;
 wire \core.muxed_new_block[110] ;
 wire \core.muxed_new_block[111] ;
 wire \core.muxed_new_block[112] ;
 wire \core.muxed_new_block[113] ;
 wire \core.muxed_new_block[114] ;
 wire \core.muxed_new_block[115] ;
 wire \core.muxed_new_block[116] ;
 wire \core.muxed_new_block[117] ;
 wire \core.muxed_new_block[118] ;
 wire \core.muxed_new_block[119] ;
 wire \core.muxed_new_block[11] ;
 wire \core.muxed_new_block[120] ;
 wire \core.muxed_new_block[121] ;
 wire \core.muxed_new_block[122] ;
 wire \core.muxed_new_block[123] ;
 wire \core.muxed_new_block[124] ;
 wire \core.muxed_new_block[125] ;
 wire \core.muxed_new_block[126] ;
 wire \core.muxed_new_block[127] ;
 wire \core.muxed_new_block[12] ;
 wire \core.muxed_new_block[13] ;
 wire \core.muxed_new_block[14] ;
 wire \core.muxed_new_block[15] ;
 wire \core.muxed_new_block[16] ;
 wire \core.muxed_new_block[17] ;
 wire \core.muxed_new_block[18] ;
 wire \core.muxed_new_block[19] ;
 wire \core.muxed_new_block[1] ;
 wire \core.muxed_new_block[20] ;
 wire \core.muxed_new_block[21] ;
 wire \core.muxed_new_block[22] ;
 wire \core.muxed_new_block[23] ;
 wire \core.muxed_new_block[24] ;
 wire \core.muxed_new_block[25] ;
 wire \core.muxed_new_block[26] ;
 wire \core.muxed_new_block[27] ;
 wire \core.muxed_new_block[28] ;
 wire \core.muxed_new_block[29] ;
 wire \core.muxed_new_block[2] ;
 wire \core.muxed_new_block[30] ;
 wire \core.muxed_new_block[31] ;
 wire \core.muxed_new_block[32] ;
 wire \core.muxed_new_block[33] ;
 wire \core.muxed_new_block[34] ;
 wire \core.muxed_new_block[35] ;
 wire \core.muxed_new_block[36] ;
 wire \core.muxed_new_block[37] ;
 wire \core.muxed_new_block[38] ;
 wire \core.muxed_new_block[39] ;
 wire \core.muxed_new_block[3] ;
 wire \core.muxed_new_block[40] ;
 wire \core.muxed_new_block[41] ;
 wire \core.muxed_new_block[42] ;
 wire \core.muxed_new_block[43] ;
 wire \core.muxed_new_block[44] ;
 wire \core.muxed_new_block[45] ;
 wire \core.muxed_new_block[46] ;
 wire \core.muxed_new_block[47] ;
 wire \core.muxed_new_block[48] ;
 wire \core.muxed_new_block[49] ;
 wire \core.muxed_new_block[4] ;
 wire \core.muxed_new_block[50] ;
 wire \core.muxed_new_block[51] ;
 wire \core.muxed_new_block[52] ;
 wire \core.muxed_new_block[53] ;
 wire \core.muxed_new_block[54] ;
 wire \core.muxed_new_block[55] ;
 wire \core.muxed_new_block[56] ;
 wire \core.muxed_new_block[57] ;
 wire \core.muxed_new_block[58] ;
 wire \core.muxed_new_block[59] ;
 wire \core.muxed_new_block[5] ;
 wire \core.muxed_new_block[60] ;
 wire \core.muxed_new_block[61] ;
 wire \core.muxed_new_block[62] ;
 wire \core.muxed_new_block[63] ;
 wire \core.muxed_new_block[64] ;
 wire \core.muxed_new_block[65] ;
 wire \core.muxed_new_block[66] ;
 wire \core.muxed_new_block[67] ;
 wire \core.muxed_new_block[68] ;
 wire \core.muxed_new_block[69] ;
 wire \core.muxed_new_block[6] ;
 wire \core.muxed_new_block[70] ;
 wire \core.muxed_new_block[71] ;
 wire \core.muxed_new_block[72] ;
 wire \core.muxed_new_block[73] ;
 wire \core.muxed_new_block[74] ;
 wire \core.muxed_new_block[75] ;
 wire \core.muxed_new_block[76] ;
 wire \core.muxed_new_block[77] ;
 wire \core.muxed_new_block[78] ;
 wire \core.muxed_new_block[79] ;
 wire \core.muxed_new_block[7] ;
 wire \core.muxed_new_block[80] ;
 wire \core.muxed_new_block[81] ;
 wire \core.muxed_new_block[82] ;
 wire \core.muxed_new_block[83] ;
 wire \core.muxed_new_block[84] ;
 wire \core.muxed_new_block[85] ;
 wire \core.muxed_new_block[86] ;
 wire \core.muxed_new_block[87] ;
 wire \core.muxed_new_block[88] ;
 wire \core.muxed_new_block[89] ;
 wire \core.muxed_new_block[8] ;
 wire \core.muxed_new_block[90] ;
 wire \core.muxed_new_block[91] ;
 wire \core.muxed_new_block[92] ;
 wire \core.muxed_new_block[93] ;
 wire \core.muxed_new_block[94] ;
 wire \core.muxed_new_block[95] ;
 wire \core.muxed_new_block[96] ;
 wire \core.muxed_new_block[97] ;
 wire \core.muxed_new_block[98] ;
 wire \core.muxed_new_block[99] ;
 wire \core.muxed_new_block[9] ;
 wire \core.next ;
 wire \core.ready ;
 wire \core.result_valid ;
 wire init_new;
 wire next_new;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire ready_reg;
 wire \result_reg[0] ;
 wire \result_reg[100] ;
 wire \result_reg[101] ;
 wire \result_reg[102] ;
 wire \result_reg[103] ;
 wire \result_reg[104] ;
 wire \result_reg[105] ;
 wire \result_reg[106] ;
 wire \result_reg[107] ;
 wire \result_reg[108] ;
 wire \result_reg[109] ;
 wire \result_reg[10] ;
 wire \result_reg[110] ;
 wire \result_reg[111] ;
 wire \result_reg[112] ;
 wire \result_reg[113] ;
 wire \result_reg[114] ;
 wire \result_reg[115] ;
 wire \result_reg[116] ;
 wire \result_reg[117] ;
 wire \result_reg[118] ;
 wire \result_reg[119] ;
 wire \result_reg[11] ;
 wire \result_reg[120] ;
 wire \result_reg[121] ;
 wire \result_reg[122] ;
 wire \result_reg[123] ;
 wire \result_reg[124] ;
 wire \result_reg[125] ;
 wire \result_reg[126] ;
 wire \result_reg[127] ;
 wire \result_reg[12] ;
 wire \result_reg[13] ;
 wire \result_reg[14] ;
 wire \result_reg[15] ;
 wire \result_reg[16] ;
 wire \result_reg[17] ;
 wire \result_reg[18] ;
 wire \result_reg[19] ;
 wire \result_reg[1] ;
 wire \result_reg[20] ;
 wire \result_reg[21] ;
 wire \result_reg[22] ;
 wire \result_reg[23] ;
 wire \result_reg[24] ;
 wire \result_reg[25] ;
 wire \result_reg[26] ;
 wire \result_reg[27] ;
 wire \result_reg[28] ;
 wire \result_reg[29] ;
 wire \result_reg[2] ;
 wire \result_reg[30] ;
 wire \result_reg[31] ;
 wire \result_reg[32] ;
 wire \result_reg[33] ;
 wire \result_reg[34] ;
 wire \result_reg[35] ;
 wire \result_reg[36] ;
 wire \result_reg[37] ;
 wire \result_reg[38] ;
 wire \result_reg[39] ;
 wire \result_reg[3] ;
 wire \result_reg[40] ;
 wire \result_reg[41] ;
 wire \result_reg[42] ;
 wire \result_reg[43] ;
 wire \result_reg[44] ;
 wire \result_reg[45] ;
 wire \result_reg[46] ;
 wire \result_reg[47] ;
 wire \result_reg[48] ;
 wire \result_reg[49] ;
 wire \result_reg[4] ;
 wire \result_reg[50] ;
 wire \result_reg[51] ;
 wire \result_reg[52] ;
 wire \result_reg[53] ;
 wire \result_reg[54] ;
 wire \result_reg[55] ;
 wire \result_reg[56] ;
 wire \result_reg[57] ;
 wire \result_reg[58] ;
 wire \result_reg[59] ;
 wire \result_reg[5] ;
 wire \result_reg[60] ;
 wire \result_reg[61] ;
 wire \result_reg[62] ;
 wire \result_reg[63] ;
 wire \result_reg[64] ;
 wire \result_reg[65] ;
 wire \result_reg[66] ;
 wire \result_reg[67] ;
 wire \result_reg[68] ;
 wire \result_reg[69] ;
 wire \result_reg[6] ;
 wire \result_reg[70] ;
 wire \result_reg[71] ;
 wire \result_reg[72] ;
 wire \result_reg[73] ;
 wire \result_reg[74] ;
 wire \result_reg[75] ;
 wire \result_reg[76] ;
 wire \result_reg[77] ;
 wire \result_reg[78] ;
 wire \result_reg[79] ;
 wire \result_reg[7] ;
 wire \result_reg[80] ;
 wire \result_reg[81] ;
 wire \result_reg[82] ;
 wire \result_reg[83] ;
 wire \result_reg[84] ;
 wire \result_reg[85] ;
 wire \result_reg[86] ;
 wire \result_reg[87] ;
 wire \result_reg[88] ;
 wire \result_reg[89] ;
 wire \result_reg[8] ;
 wire \result_reg[90] ;
 wire \result_reg[91] ;
 wire \result_reg[92] ;
 wire \result_reg[93] ;
 wire \result_reg[94] ;
 wire \result_reg[95] ;
 wire \result_reg[96] ;
 wire \result_reg[97] ;
 wire \result_reg[98] ;
 wire \result_reg[99] ;
 wire \result_reg[9] ;
 wire valid_reg;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_leaf_327_clk;
 wire clknet_leaf_328_clk;
 wire clknet_leaf_329_clk;
 wire clknet_leaf_330_clk;
 wire clknet_leaf_331_clk;
 wire clknet_leaf_332_clk;
 wire clknet_leaf_333_clk;
 wire clknet_leaf_334_clk;
 wire clknet_leaf_335_clk;
 wire clknet_leaf_336_clk;
 wire clknet_leaf_337_clk;
 wire clknet_leaf_338_clk;
 wire clknet_leaf_339_clk;
 wire clknet_leaf_340_clk;
 wire clknet_leaf_341_clk;
 wire clknet_leaf_342_clk;
 wire clknet_leaf_343_clk;
 wire clknet_leaf_344_clk;
 wire clknet_leaf_345_clk;
 wire clknet_leaf_346_clk;
 wire clknet_leaf_347_clk;
 wire clknet_leaf_348_clk;
 wire clknet_leaf_349_clk;
 wire clknet_leaf_350_clk;
 wire clknet_leaf_351_clk;
 wire clknet_leaf_352_clk;
 wire clknet_leaf_353_clk;
 wire clknet_leaf_354_clk;
 wire clknet_leaf_355_clk;
 wire clknet_leaf_356_clk;
 wire clknet_leaf_357_clk;
 wire clknet_leaf_358_clk;
 wire clknet_leaf_359_clk;
 wire clknet_leaf_360_clk;
 wire clknet_leaf_361_clk;
 wire clknet_leaf_362_clk;
 wire clknet_leaf_363_clk;
 wire clknet_leaf_364_clk;
 wire clknet_leaf_365_clk;
 wire clknet_leaf_366_clk;
 wire clknet_leaf_367_clk;
 wire clknet_leaf_368_clk;
 wire clknet_leaf_369_clk;
 wire clknet_leaf_370_clk;
 wire clknet_leaf_371_clk;
 wire clknet_leaf_372_clk;
 wire clknet_leaf_373_clk;
 wire clknet_leaf_374_clk;
 wire clknet_leaf_375_clk;
 wire clknet_leaf_376_clk;
 wire clknet_leaf_377_clk;
 wire clknet_leaf_378_clk;
 wire clknet_leaf_379_clk;
 wire clknet_leaf_380_clk;
 wire clknet_leaf_381_clk;
 wire clknet_leaf_382_clk;
 wire clknet_leaf_383_clk;
 wire clknet_leaf_384_clk;
 wire clknet_leaf_385_clk;
 wire clknet_leaf_386_clk;
 wire clknet_leaf_387_clk;
 wire clknet_leaf_388_clk;
 wire clknet_leaf_389_clk;
 wire clknet_leaf_390_clk;
 wire clknet_leaf_391_clk;
 wire clknet_leaf_392_clk;
 wire clknet_leaf_393_clk;
 wire clknet_leaf_394_clk;
 wire clknet_leaf_395_clk;
 wire clknet_leaf_396_clk;
 wire clknet_leaf_397_clk;
 wire clknet_leaf_398_clk;
 wire clknet_leaf_399_clk;
 wire clknet_leaf_400_clk;
 wire clknet_leaf_401_clk;
 wire clknet_leaf_402_clk;
 wire clknet_leaf_403_clk;
 wire clknet_leaf_404_clk;
 wire clknet_leaf_405_clk;
 wire clknet_leaf_406_clk;
 wire clknet_leaf_407_clk;
 wire clknet_leaf_408_clk;
 wire clknet_leaf_409_clk;
 wire clknet_leaf_410_clk;
 wire clknet_leaf_411_clk;
 wire clknet_leaf_412_clk;
 wire clknet_leaf_413_clk;
 wire clknet_leaf_414_clk;
 wire clknet_leaf_415_clk;
 wire clknet_leaf_416_clk;
 wire clknet_leaf_417_clk;
 wire clknet_leaf_418_clk;
 wire clknet_leaf_419_clk;
 wire clknet_leaf_420_clk;
 wire clknet_leaf_421_clk;
 wire clknet_leaf_422_clk;
 wire clknet_leaf_423_clk;
 wire clknet_leaf_424_clk;
 wire clknet_leaf_425_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 BUF_X2 _22140_ (.A(\core.aes_core_ctrl_reg[2] ),
    .Z(_16200_));
 BUF_X2 _22141_ (.A(\core.encdec ),
    .Z(_16201_));
 BUF_X4 _22142_ (.A(_16201_),
    .Z(_16202_));
 BUF_X8 _22143_ (.A(_16202_),
    .Z(_16203_));
 MUX2_X2 _22144_ (.A(\core.dec_block.ready ),
    .B(\core.enc_block.ready ),
    .S(_16203_),
    .Z(_16204_));
 AOI22_X4 _22145_ (.A1(\core.key_ready ),
    .A2(_16200_),
    .B1(\core.aes_core_ctrl_reg[1] ),
    .B2(_16204_),
    .ZN(_16205_));
 BUF_X4 _22146_ (.A(\core.next ),
    .Z(_16206_));
 NAND2_X1 _22147_ (.A1(_16206_),
    .A2(\core.aes_core_ctrl_reg[0] ),
    .ZN(_16207_));
 NAND3_X1 _22148_ (.A1(_16200_),
    .A2(_16205_),
    .A3(_16207_),
    .ZN(_16208_));
 INV_X1 _22149_ (.A(\core.aes_core_ctrl_reg[0] ),
    .ZN(_16209_));
 BUF_X4 _22150_ (.A(\core.init ),
    .Z(_16210_));
 INV_X2 _22151_ (.A(_16210_),
    .ZN(_16211_));
 OAI21_X1 _22152_ (.A(_16208_),
    .B1(_16209_),
    .B2(_16211_),
    .ZN(_00008_));
 AND2_X1 _22153_ (.A1(_16210_),
    .A2(\core.aes_core_ctrl_reg[0] ),
    .ZN(_16212_));
 NAND2_X1 _22154_ (.A1(\core.aes_core_ctrl_reg[1] ),
    .A2(_16205_),
    .ZN(_16213_));
 AOI21_X1 _22155_ (.A(_16212_),
    .B1(_16207_),
    .B2(_16213_),
    .ZN(_00007_));
 INV_X2 _22156_ (.A(net2),
    .ZN(_22094_));
 NAND2_X1 _22157_ (.A1(_16210_),
    .A2(\core.keymem.key_mem_ctrl_reg[0] ),
    .ZN(_16214_));
 INV_X1 _22158_ (.A(_16214_),
    .ZN(_00004_));
 INV_X1 _22159_ (.A(\core.keymem.key_mem_ctrl_reg[2] ),
    .ZN(_16215_));
 BUF_X2 _22160_ (.A(_22108_),
    .Z(_16216_));
 INV_X1 _22161_ (.A(_16216_),
    .ZN(_16217_));
 BUF_X4 _22162_ (.A(\core.keymem.round_ctr_reg[2] ),
    .Z(_16218_));
 BUF_X8 _22163_ (.A(\core.dec_block.keylen ),
    .Z(_16219_));
 XOR2_X2 _22164_ (.A(_16218_),
    .B(_16219_),
    .Z(_16220_));
 NOR3_X2 _22165_ (.A1(_00319_),
    .A2(_16217_),
    .A3(_16220_),
    .ZN(_16221_));
 BUF_X4 _22166_ (.A(\core.keymem.key_mem_ctrl_reg[1] ),
    .Z(_16222_));
 AOI21_X1 _22167_ (.A(_00004_),
    .B1(_16221_),
    .B2(_16222_),
    .ZN(_16223_));
 BUF_X4 _22168_ (.A(_00318_),
    .Z(_16224_));
 AOI21_X1 _22169_ (.A(_16223_),
    .B1(_00320_),
    .B2(_16224_),
    .ZN(_16225_));
 OR3_X1 _22170_ (.A1(\core.keymem.key_mem_ctrl_reg[2] ),
    .A2(\core.keymem.key_mem_ctrl_reg[3] ),
    .A3(_16225_),
    .ZN(_16226_));
 OAI21_X1 _22171_ (.A(_16215_),
    .B1(_16226_),
    .B2(_16224_),
    .ZN(_00014_));
 INV_X1 _22172_ (.A(_16221_),
    .ZN(_16227_));
 BUF_X8 _22173_ (.A(_16222_),
    .Z(_16228_));
 BUF_X8 _22174_ (.A(_16228_),
    .Z(_16229_));
 AOI221_X1 _22175_ (.A(\core.keymem.key_mem_ctrl_reg[3] ),
    .B1(\core.keymem.key_mem_ctrl_reg[0] ),
    .B2(_16211_),
    .C1(_16227_),
    .C2(_16229_),
    .ZN(_16230_));
 MUX2_X1 _22176_ (.A(_00320_),
    .B(_16230_),
    .S(_16226_),
    .Z(_16231_));
 INV_X1 _22177_ (.A(_16231_),
    .ZN(_00013_));
 CLKBUF_X3 _22178_ (.A(\core.enc_block.enc_ctrl_reg[2] ),
    .Z(_16232_));
 INV_X1 _22179_ (.A(_16232_),
    .ZN(_16233_));
 BUF_X4 _22180_ (.A(\core.enc_block.enc_ctrl_reg[3] ),
    .Z(_16234_));
 INV_X4 _22181_ (.A(_16234_),
    .ZN(_16235_));
 BUF_X4 _22182_ (.A(\core.enc_block.round[1] ),
    .Z(_16236_));
 AOI21_X2 _22183_ (.A(_22092_),
    .B1(_22093_),
    .B2(_16236_),
    .ZN(_16237_));
 NOR3_X2 _22184_ (.A1(_16235_),
    .A2(_00323_),
    .A3(_16237_),
    .ZN(_16238_));
 BUF_X4 _22185_ (.A(_00321_),
    .Z(_16239_));
 INV_X2 _22186_ (.A(_16239_),
    .ZN(_16240_));
 AND3_X4 _22187_ (.A1(_16203_),
    .A2(_16206_),
    .A3(\core.enc_block.enc_ctrl_reg[0] ),
    .ZN(_16241_));
 BUF_X2 _22188_ (.A(_22124_),
    .Z(_16242_));
 BUF_X2 _22189_ (.A(\core.enc_block.enc_ctrl_reg[1] ),
    .Z(_16243_));
 AOI21_X2 _22190_ (.A(_16241_),
    .B1(_16242_),
    .B2(_16243_),
    .ZN(_16244_));
 AOI21_X1 _22191_ (.A(_16234_),
    .B1(_16240_),
    .B2(_16244_),
    .ZN(_16245_));
 OAI21_X1 _22192_ (.A(_16233_),
    .B1(_16238_),
    .B2(_16245_),
    .ZN(_00012_));
 INV_X2 _22193_ (.A(_16238_),
    .ZN(_16246_));
 INV_X1 _22194_ (.A(\core.enc_block.enc_ctrl_reg[0] ),
    .ZN(_16247_));
 AOI21_X1 _22195_ (.A(_16247_),
    .B1(_16206_),
    .B2(_16203_),
    .ZN(_16248_));
 NOR2_X4 _22196_ (.A1(_16234_),
    .A2(_16232_),
    .ZN(_16249_));
 INV_X2 _22197_ (.A(_16242_),
    .ZN(_16250_));
 BUF_X4 _22198_ (.A(_16250_),
    .Z(_16251_));
 BUF_X4 _22199_ (.A(_16251_),
    .Z(_16252_));
 AOI221_X2 _22200_ (.A(_16248_),
    .B1(_16249_),
    .B2(_16244_),
    .C1(_16243_),
    .C2(_16252_),
    .ZN(_16253_));
 OR2_X1 _22201_ (.A1(_16239_),
    .A2(_16244_),
    .ZN(_16254_));
 AND3_X1 _22202_ (.A1(_00322_),
    .A2(_16249_),
    .A3(_16254_),
    .ZN(_16255_));
 OAI21_X1 _22203_ (.A(_16246_),
    .B1(_16253_),
    .B2(_16255_),
    .ZN(_00011_));
 NOR2_X1 _22204_ (.A1(_16210_),
    .A2(_16206_),
    .ZN(_16256_));
 NOR3_X1 _22205_ (.A1(_16200_),
    .A2(\core.aes_core_ctrl_reg[1] ),
    .A3(_16256_),
    .ZN(_16257_));
 OAI21_X1 _22206_ (.A(_16205_),
    .B1(_16257_),
    .B2(_16209_),
    .ZN(_00006_));
 BUF_X4 _22207_ (.A(\core.dec_block.dec_ctrl_reg[3] ),
    .Z(_16258_));
 INV_X4 _22208_ (.A(_16258_),
    .ZN(_16259_));
 BUF_X4 _22209_ (.A(_00324_),
    .Z(_16260_));
 INV_X2 _22210_ (.A(_16260_),
    .ZN(_16261_));
 INV_X4 _22211_ (.A(_16201_),
    .ZN(_16262_));
 AND2_X2 _22212_ (.A1(_16262_),
    .A2(_16206_),
    .ZN(_16263_));
 NAND2_X4 _22213_ (.A1(\core.dec_block.dec_ctrl_reg[0] ),
    .A2(_16263_),
    .ZN(_16264_));
 BUF_X4 _22214_ (.A(_22138_),
    .Z(_16265_));
 BUF_X4 _22215_ (.A(_16265_),
    .Z(_16266_));
 BUF_X4 _22216_ (.A(_16266_),
    .Z(_16267_));
 BUF_X4 _22217_ (.A(_16267_),
    .Z(_16268_));
 NAND2_X4 _22218_ (.A1(\core.dec_block.dec_ctrl_reg[1] ),
    .A2(_16268_),
    .ZN(_16269_));
 NAND4_X1 _22219_ (.A1(_16259_),
    .A2(_16261_),
    .A3(_16264_),
    .A4(_16269_),
    .ZN(_16270_));
 CLKBUF_X2 _22220_ (.A(\core.dec_block.dec_ctrl_reg[2] ),
    .Z(_16271_));
 BUF_X4 _22221_ (.A(\core.dec_block.round[2] ),
    .Z(_16272_));
 BUF_X4 _22222_ (.A(\core.dec_block.round[3] ),
    .Z(_16273_));
 NOR2_X2 _22223_ (.A1(_16272_),
    .A2(_16273_),
    .ZN(_16274_));
 AND2_X2 _22224_ (.A1(_22128_),
    .A2(_16274_),
    .ZN(_16275_));
 NOR2_X2 _22225_ (.A1(_16259_),
    .A2(_16275_),
    .ZN(_16276_));
 NOR2_X1 _22226_ (.A1(_16271_),
    .A2(_16276_),
    .ZN(_16277_));
 NAND2_X1 _22227_ (.A1(_16270_),
    .A2(_16277_),
    .ZN(_00010_));
 INV_X2 _22228_ (.A(\core.dec_block.dec_ctrl_reg[1] ),
    .ZN(_16278_));
 NOR2_X1 _22229_ (.A1(_16278_),
    .A2(_16268_),
    .ZN(_16279_));
 INV_X1 _22230_ (.A(_16263_),
    .ZN(_16280_));
 AOI21_X1 _22231_ (.A(_16279_),
    .B1(_16280_),
    .B2(\core.dec_block.dec_ctrl_reg[0] ),
    .ZN(_16281_));
 AOI22_X2 _22232_ (.A1(_00325_),
    .A2(_16260_),
    .B1(_16264_),
    .B2(_16269_),
    .ZN(_16282_));
 NOR2_X1 _22233_ (.A1(_16271_),
    .A2(_16282_),
    .ZN(_16283_));
 MUX2_X1 _22234_ (.A(_16281_),
    .B(_00325_),
    .S(_16283_),
    .Z(_16284_));
 AOI22_X1 _22235_ (.A1(_16276_),
    .A2(_16281_),
    .B1(_16284_),
    .B2(_16259_),
    .ZN(_00009_));
 BUF_X4 _22236_ (.A(_16229_),
    .Z(_16285_));
 CLKBUF_X3 _22237_ (.A(_16285_),
    .Z(_16286_));
 AND3_X1 _22238_ (.A1(_16286_),
    .A2(_16221_),
    .A3(_16226_),
    .ZN(_00005_));
 NAND3_X1 _22239_ (.A1(_00322_),
    .A2(_16239_),
    .A3(_16249_),
    .ZN(_16287_));
 AND3_X1 _22240_ (.A1(_16243_),
    .A2(_16242_),
    .A3(_16287_),
    .ZN(_00003_));
 AND2_X1 _22241_ (.A1(_16241_),
    .A2(_16287_),
    .ZN(_00002_));
 NOR3_X1 _22242_ (.A1(_16258_),
    .A2(_16271_),
    .A3(_16282_),
    .ZN(_16288_));
 NOR2_X1 _22243_ (.A1(_16269_),
    .A2(_16288_),
    .ZN(_00001_));
 NOR2_X1 _22244_ (.A1(_16264_),
    .A2(_16288_),
    .ZN(_00000_));
 INV_X2 _22245_ (.A(net3),
    .ZN(_22095_));
 BUF_X4 _22246_ (.A(net18),
    .Z(_16289_));
 INV_X1 _22247_ (.A(net5),
    .ZN(_16290_));
 INV_X2 _22248_ (.A(net1),
    .ZN(_16291_));
 BUF_X4 _22249_ (.A(address[0]),
    .Z(_16292_));
 INV_X4 _22250_ (.A(_16292_),
    .ZN(_16293_));
 NOR2_X4 _22251_ (.A1(_16291_),
    .A2(_16293_),
    .ZN(_16294_));
 AOI21_X1 _22252_ (.A(_22098_),
    .B1(_22096_),
    .B2(_16294_),
    .ZN(_16295_));
 OR4_X4 _22253_ (.A1(net6),
    .A2(net7),
    .A3(_16290_),
    .A4(_16295_),
    .ZN(_16296_));
 NAND2_X4 _22254_ (.A1(net17),
    .A2(net8),
    .ZN(_16297_));
 NOR3_X4 _22255_ (.A1(net4),
    .A2(_16296_),
    .A3(_16297_),
    .ZN(_16298_));
 NOR2_X4 _22256_ (.A1(net1),
    .A2(_16292_),
    .ZN(_16299_));
 NAND2_X4 _22257_ (.A1(_16298_),
    .A2(_16299_),
    .ZN(_16300_));
 BUF_X4 _22258_ (.A(_16300_),
    .Z(_16301_));
 MUX2_X1 _22259_ (.A(_16289_),
    .B(\block_reg[0][0] ),
    .S(_16301_),
    .Z(_00439_));
 BUF_X4 _22260_ (.A(net19),
    .Z(_16302_));
 MUX2_X1 _22261_ (.A(_16302_),
    .B(\block_reg[0][10] ),
    .S(_16301_),
    .Z(_00440_));
 BUF_X4 _22262_ (.A(net20),
    .Z(_16303_));
 MUX2_X1 _22263_ (.A(_16303_),
    .B(\block_reg[0][11] ),
    .S(_16301_),
    .Z(_00441_));
 BUF_X4 _22264_ (.A(net21),
    .Z(_16304_));
 MUX2_X1 _22265_ (.A(_16304_),
    .B(\block_reg[0][12] ),
    .S(_16301_),
    .Z(_00442_));
 BUF_X4 _22266_ (.A(net22),
    .Z(_16305_));
 MUX2_X1 _22267_ (.A(_16305_),
    .B(\block_reg[0][13] ),
    .S(_16301_),
    .Z(_00443_));
 BUF_X4 _22268_ (.A(net23),
    .Z(_16306_));
 MUX2_X1 _22269_ (.A(_16306_),
    .B(\block_reg[0][14] ),
    .S(_16301_),
    .Z(_00444_));
 CLKBUF_X3 _22270_ (.A(net24),
    .Z(_16307_));
 MUX2_X1 _22271_ (.A(_16307_),
    .B(\block_reg[0][15] ),
    .S(_16301_),
    .Z(_00445_));
 BUF_X4 _22272_ (.A(net25),
    .Z(_16308_));
 MUX2_X1 _22273_ (.A(_16308_),
    .B(\block_reg[0][16] ),
    .S(_16301_),
    .Z(_00446_));
 CLKBUF_X3 _22274_ (.A(net26),
    .Z(_16309_));
 MUX2_X1 _22275_ (.A(_16309_),
    .B(\block_reg[0][17] ),
    .S(_16301_),
    .Z(_00447_));
 BUF_X4 _22276_ (.A(net27),
    .Z(_16310_));
 MUX2_X1 _22277_ (.A(_16310_),
    .B(\block_reg[0][18] ),
    .S(_16301_),
    .Z(_00448_));
 BUF_X4 _22278_ (.A(net28),
    .Z(_16311_));
 CLKBUF_X3 _22279_ (.A(_16300_),
    .Z(_16312_));
 MUX2_X1 _22280_ (.A(_16311_),
    .B(\block_reg[0][19] ),
    .S(_16312_),
    .Z(_00449_));
 BUF_X4 _22281_ (.A(net29),
    .Z(_16313_));
 MUX2_X1 _22282_ (.A(_16313_),
    .B(\block_reg[0][1] ),
    .S(_16312_),
    .Z(_00450_));
 BUF_X4 _22283_ (.A(net30),
    .Z(_16314_));
 MUX2_X1 _22284_ (.A(_16314_),
    .B(\block_reg[0][20] ),
    .S(_16312_),
    .Z(_00451_));
 BUF_X4 _22285_ (.A(net31),
    .Z(_16315_));
 MUX2_X1 _22286_ (.A(_16315_),
    .B(\block_reg[0][21] ),
    .S(_16312_),
    .Z(_00452_));
 CLKBUF_X3 _22287_ (.A(net32),
    .Z(_16316_));
 MUX2_X1 _22288_ (.A(_16316_),
    .B(\block_reg[0][22] ),
    .S(_16312_),
    .Z(_00453_));
 BUF_X4 _22289_ (.A(net33),
    .Z(_16317_));
 MUX2_X1 _22290_ (.A(_16317_),
    .B(\block_reg[0][23] ),
    .S(_16312_),
    .Z(_00454_));
 BUF_X4 _22291_ (.A(net34),
    .Z(_16318_));
 MUX2_X1 _22292_ (.A(_16318_),
    .B(\block_reg[0][24] ),
    .S(_16312_),
    .Z(_00455_));
 BUF_X4 _22293_ (.A(net35),
    .Z(_16319_));
 MUX2_X1 _22294_ (.A(_16319_),
    .B(\block_reg[0][25] ),
    .S(_16312_),
    .Z(_00456_));
 BUF_X4 _22295_ (.A(net36),
    .Z(_16320_));
 MUX2_X1 _22296_ (.A(_16320_),
    .B(\block_reg[0][26] ),
    .S(_16312_),
    .Z(_00457_));
 BUF_X4 _22297_ (.A(net37),
    .Z(_16321_));
 MUX2_X1 _22298_ (.A(_16321_),
    .B(\block_reg[0][27] ),
    .S(_16312_),
    .Z(_00458_));
 BUF_X4 _22299_ (.A(net38),
    .Z(_16322_));
 BUF_X4 _22300_ (.A(_16300_),
    .Z(_16323_));
 MUX2_X1 _22301_ (.A(_16322_),
    .B(\block_reg[0][28] ),
    .S(_16323_),
    .Z(_00459_));
 BUF_X4 _22302_ (.A(net39),
    .Z(_16324_));
 MUX2_X1 _22303_ (.A(_16324_),
    .B(\block_reg[0][29] ),
    .S(_16323_),
    .Z(_00460_));
 BUF_X4 _22304_ (.A(net40),
    .Z(_16325_));
 MUX2_X1 _22305_ (.A(_16325_),
    .B(\block_reg[0][2] ),
    .S(_16323_),
    .Z(_00461_));
 BUF_X4 _22306_ (.A(net41),
    .Z(_16326_));
 MUX2_X1 _22307_ (.A(_16326_),
    .B(\block_reg[0][30] ),
    .S(_16323_),
    .Z(_00462_));
 BUF_X4 _22308_ (.A(net42),
    .Z(_16327_));
 MUX2_X1 _22309_ (.A(_16327_),
    .B(\block_reg[0][31] ),
    .S(_16323_),
    .Z(_00463_));
 BUF_X4 _22310_ (.A(net43),
    .Z(_16328_));
 MUX2_X1 _22311_ (.A(_16328_),
    .B(\block_reg[0][3] ),
    .S(_16323_),
    .Z(_00464_));
 BUF_X4 _22312_ (.A(net44),
    .Z(_16329_));
 MUX2_X1 _22313_ (.A(_16329_),
    .B(\block_reg[0][4] ),
    .S(_16323_),
    .Z(_00465_));
 BUF_X4 _22314_ (.A(net45),
    .Z(_16330_));
 MUX2_X1 _22315_ (.A(_16330_),
    .B(\block_reg[0][5] ),
    .S(_16323_),
    .Z(_00466_));
 BUF_X4 _22316_ (.A(net46),
    .Z(_16331_));
 MUX2_X1 _22317_ (.A(_16331_),
    .B(\block_reg[0][6] ),
    .S(_16323_),
    .Z(_00467_));
 BUF_X4 _22318_ (.A(net47),
    .Z(_16332_));
 MUX2_X1 _22319_ (.A(_16332_),
    .B(\block_reg[0][7] ),
    .S(_16323_),
    .Z(_00468_));
 BUF_X4 _22320_ (.A(net48),
    .Z(_16333_));
 MUX2_X1 _22321_ (.A(_16333_),
    .B(\block_reg[0][8] ),
    .S(_16300_),
    .Z(_00469_));
 BUF_X4 _22322_ (.A(net49),
    .Z(_16334_));
 MUX2_X1 _22323_ (.A(_16334_),
    .B(\block_reg[0][9] ),
    .S(_16300_),
    .Z(_00470_));
 BUF_X4 _22324_ (.A(net1),
    .Z(_16335_));
 NOR2_X2 _22325_ (.A1(_16335_),
    .A2(_16293_),
    .ZN(_16336_));
 NAND2_X4 _22326_ (.A1(_16298_),
    .A2(_16336_),
    .ZN(_16337_));
 BUF_X4 _22327_ (.A(_16337_),
    .Z(_16338_));
 MUX2_X1 _22328_ (.A(_16289_),
    .B(\block_reg[1][0] ),
    .S(_16338_),
    .Z(_00471_));
 MUX2_X1 _22329_ (.A(_16302_),
    .B(\block_reg[1][10] ),
    .S(_16338_),
    .Z(_00472_));
 MUX2_X1 _22330_ (.A(_16303_),
    .B(\block_reg[1][11] ),
    .S(_16338_),
    .Z(_00473_));
 MUX2_X1 _22331_ (.A(_16304_),
    .B(\block_reg[1][12] ),
    .S(_16338_),
    .Z(_00474_));
 MUX2_X1 _22332_ (.A(_16305_),
    .B(\block_reg[1][13] ),
    .S(_16338_),
    .Z(_00475_));
 MUX2_X1 _22333_ (.A(_16306_),
    .B(\block_reg[1][14] ),
    .S(_16338_),
    .Z(_00476_));
 MUX2_X1 _22334_ (.A(_16307_),
    .B(\block_reg[1][15] ),
    .S(_16338_),
    .Z(_00477_));
 MUX2_X1 _22335_ (.A(_16308_),
    .B(\block_reg[1][16] ),
    .S(_16338_),
    .Z(_00478_));
 MUX2_X1 _22336_ (.A(_16309_),
    .B(\block_reg[1][17] ),
    .S(_16338_),
    .Z(_00479_));
 MUX2_X1 _22337_ (.A(_16310_),
    .B(\block_reg[1][18] ),
    .S(_16338_),
    .Z(_00480_));
 CLKBUF_X3 _22338_ (.A(_16337_),
    .Z(_16339_));
 MUX2_X1 _22339_ (.A(_16311_),
    .B(\block_reg[1][19] ),
    .S(_16339_),
    .Z(_00481_));
 MUX2_X1 _22340_ (.A(_16313_),
    .B(\block_reg[1][1] ),
    .S(_16339_),
    .Z(_00482_));
 MUX2_X1 _22341_ (.A(_16314_),
    .B(\block_reg[1][20] ),
    .S(_16339_),
    .Z(_00483_));
 MUX2_X1 _22342_ (.A(_16315_),
    .B(\block_reg[1][21] ),
    .S(_16339_),
    .Z(_00484_));
 MUX2_X1 _22343_ (.A(_16316_),
    .B(\block_reg[1][22] ),
    .S(_16339_),
    .Z(_00485_));
 MUX2_X1 _22344_ (.A(_16317_),
    .B(\block_reg[1][23] ),
    .S(_16339_),
    .Z(_00486_));
 MUX2_X1 _22345_ (.A(_16318_),
    .B(\block_reg[1][24] ),
    .S(_16339_),
    .Z(_00487_));
 MUX2_X1 _22346_ (.A(_16319_),
    .B(\block_reg[1][25] ),
    .S(_16339_),
    .Z(_00488_));
 MUX2_X1 _22347_ (.A(_16320_),
    .B(\block_reg[1][26] ),
    .S(_16339_),
    .Z(_00489_));
 MUX2_X1 _22348_ (.A(_16321_),
    .B(\block_reg[1][27] ),
    .S(_16339_),
    .Z(_00490_));
 BUF_X4 _22349_ (.A(_16337_),
    .Z(_16340_));
 MUX2_X1 _22350_ (.A(_16322_),
    .B(\block_reg[1][28] ),
    .S(_16340_),
    .Z(_00491_));
 MUX2_X1 _22351_ (.A(_16324_),
    .B(\block_reg[1][29] ),
    .S(_16340_),
    .Z(_00492_));
 MUX2_X1 _22352_ (.A(_16325_),
    .B(\block_reg[1][2] ),
    .S(_16340_),
    .Z(_00493_));
 MUX2_X1 _22353_ (.A(_16326_),
    .B(\block_reg[1][30] ),
    .S(_16340_),
    .Z(_00494_));
 MUX2_X1 _22354_ (.A(_16327_),
    .B(\block_reg[1][31] ),
    .S(_16340_),
    .Z(_00495_));
 MUX2_X1 _22355_ (.A(_16328_),
    .B(\block_reg[1][3] ),
    .S(_16340_),
    .Z(_00496_));
 MUX2_X1 _22356_ (.A(_16329_),
    .B(\block_reg[1][4] ),
    .S(_16340_),
    .Z(_00497_));
 MUX2_X1 _22357_ (.A(_16330_),
    .B(\block_reg[1][5] ),
    .S(_16340_),
    .Z(_00498_));
 MUX2_X1 _22358_ (.A(_16331_),
    .B(\block_reg[1][6] ),
    .S(_16340_),
    .Z(_00499_));
 MUX2_X1 _22359_ (.A(_16332_),
    .B(\block_reg[1][7] ),
    .S(_16340_),
    .Z(_00500_));
 MUX2_X1 _22360_ (.A(_16333_),
    .B(\block_reg[1][8] ),
    .S(_16337_),
    .Z(_00501_));
 MUX2_X1 _22361_ (.A(_16334_),
    .B(\block_reg[1][9] ),
    .S(_16337_),
    .Z(_00502_));
 BUF_X4 _22362_ (.A(_16292_),
    .Z(_16341_));
 NOR2_X2 _22363_ (.A1(_16291_),
    .A2(_16341_),
    .ZN(_16342_));
 NAND2_X4 _22364_ (.A1(_16298_),
    .A2(_16342_),
    .ZN(_16343_));
 BUF_X4 _22365_ (.A(_16343_),
    .Z(_16344_));
 MUX2_X1 _22366_ (.A(_16289_),
    .B(\block_reg[2][0] ),
    .S(_16344_),
    .Z(_00503_));
 MUX2_X1 _22367_ (.A(_16302_),
    .B(\block_reg[2][10] ),
    .S(_16344_),
    .Z(_00504_));
 MUX2_X1 _22368_ (.A(_16303_),
    .B(\block_reg[2][11] ),
    .S(_16344_),
    .Z(_00505_));
 MUX2_X1 _22369_ (.A(_16304_),
    .B(\block_reg[2][12] ),
    .S(_16344_),
    .Z(_00506_));
 MUX2_X1 _22370_ (.A(_16305_),
    .B(\block_reg[2][13] ),
    .S(_16344_),
    .Z(_00507_));
 MUX2_X1 _22371_ (.A(_16306_),
    .B(\block_reg[2][14] ),
    .S(_16344_),
    .Z(_00508_));
 MUX2_X1 _22372_ (.A(_16307_),
    .B(\block_reg[2][15] ),
    .S(_16344_),
    .Z(_00509_));
 MUX2_X1 _22373_ (.A(_16308_),
    .B(\block_reg[2][16] ),
    .S(_16344_),
    .Z(_00510_));
 MUX2_X1 _22374_ (.A(_16309_),
    .B(\block_reg[2][17] ),
    .S(_16344_),
    .Z(_00511_));
 MUX2_X1 _22375_ (.A(_16310_),
    .B(\block_reg[2][18] ),
    .S(_16344_),
    .Z(_00512_));
 CLKBUF_X3 _22376_ (.A(_16343_),
    .Z(_16345_));
 MUX2_X1 _22377_ (.A(_16311_),
    .B(\block_reg[2][19] ),
    .S(_16345_),
    .Z(_00513_));
 MUX2_X1 _22378_ (.A(_16313_),
    .B(\block_reg[2][1] ),
    .S(_16345_),
    .Z(_00514_));
 MUX2_X1 _22379_ (.A(_16314_),
    .B(\block_reg[2][20] ),
    .S(_16345_),
    .Z(_00515_));
 MUX2_X1 _22380_ (.A(_16315_),
    .B(\block_reg[2][21] ),
    .S(_16345_),
    .Z(_00516_));
 MUX2_X1 _22381_ (.A(_16316_),
    .B(\block_reg[2][22] ),
    .S(_16345_),
    .Z(_00517_));
 MUX2_X1 _22382_ (.A(_16317_),
    .B(\block_reg[2][23] ),
    .S(_16345_),
    .Z(_00518_));
 MUX2_X1 _22383_ (.A(_16318_),
    .B(\block_reg[2][24] ),
    .S(_16345_),
    .Z(_00519_));
 MUX2_X1 _22384_ (.A(_16319_),
    .B(\block_reg[2][25] ),
    .S(_16345_),
    .Z(_00520_));
 MUX2_X1 _22385_ (.A(_16320_),
    .B(\block_reg[2][26] ),
    .S(_16345_),
    .Z(_00521_));
 MUX2_X1 _22386_ (.A(_16321_),
    .B(\block_reg[2][27] ),
    .S(_16345_),
    .Z(_00522_));
 BUF_X4 _22387_ (.A(_16343_),
    .Z(_16346_));
 MUX2_X1 _22388_ (.A(_16322_),
    .B(\block_reg[2][28] ),
    .S(_16346_),
    .Z(_00523_));
 MUX2_X1 _22389_ (.A(_16324_),
    .B(\block_reg[2][29] ),
    .S(_16346_),
    .Z(_00524_));
 MUX2_X1 _22390_ (.A(_16325_),
    .B(\block_reg[2][2] ),
    .S(_16346_),
    .Z(_00525_));
 MUX2_X1 _22391_ (.A(_16326_),
    .B(\block_reg[2][30] ),
    .S(_16346_),
    .Z(_00526_));
 MUX2_X1 _22392_ (.A(_16327_),
    .B(\block_reg[2][31] ),
    .S(_16346_),
    .Z(_00527_));
 MUX2_X1 _22393_ (.A(_16328_),
    .B(\block_reg[2][3] ),
    .S(_16346_),
    .Z(_00528_));
 MUX2_X1 _22394_ (.A(_16329_),
    .B(\block_reg[2][4] ),
    .S(_16346_),
    .Z(_00529_));
 MUX2_X1 _22395_ (.A(_16330_),
    .B(\block_reg[2][5] ),
    .S(_16346_),
    .Z(_00530_));
 MUX2_X1 _22396_ (.A(_16331_),
    .B(\block_reg[2][6] ),
    .S(_16346_),
    .Z(_00531_));
 MUX2_X1 _22397_ (.A(_16332_),
    .B(\block_reg[2][7] ),
    .S(_16346_),
    .Z(_00532_));
 MUX2_X1 _22398_ (.A(_16333_),
    .B(\block_reg[2][8] ),
    .S(_16343_),
    .Z(_00533_));
 MUX2_X1 _22399_ (.A(_16334_),
    .B(\block_reg[2][9] ),
    .S(_16343_),
    .Z(_00534_));
 NAND2_X4 _22400_ (.A1(_16294_),
    .A2(_16298_),
    .ZN(_16347_));
 BUF_X4 _22401_ (.A(_16347_),
    .Z(_16348_));
 MUX2_X1 _22402_ (.A(_16289_),
    .B(\block_reg[3][0] ),
    .S(_16348_),
    .Z(_00535_));
 MUX2_X1 _22403_ (.A(_16302_),
    .B(\block_reg[3][10] ),
    .S(_16348_),
    .Z(_00536_));
 MUX2_X1 _22404_ (.A(_16303_),
    .B(\block_reg[3][11] ),
    .S(_16348_),
    .Z(_00537_));
 MUX2_X1 _22405_ (.A(_16304_),
    .B(\block_reg[3][12] ),
    .S(_16348_),
    .Z(_00538_));
 MUX2_X1 _22406_ (.A(_16305_),
    .B(\block_reg[3][13] ),
    .S(_16348_),
    .Z(_00539_));
 MUX2_X1 _22407_ (.A(_16306_),
    .B(\block_reg[3][14] ),
    .S(_16348_),
    .Z(_00540_));
 MUX2_X1 _22408_ (.A(_16307_),
    .B(\block_reg[3][15] ),
    .S(_16348_),
    .Z(_00541_));
 MUX2_X1 _22409_ (.A(_16308_),
    .B(\block_reg[3][16] ),
    .S(_16348_),
    .Z(_00542_));
 MUX2_X1 _22410_ (.A(_16309_),
    .B(\block_reg[3][17] ),
    .S(_16348_),
    .Z(_00543_));
 MUX2_X1 _22411_ (.A(_16310_),
    .B(\block_reg[3][18] ),
    .S(_16348_),
    .Z(_00544_));
 CLKBUF_X3 _22412_ (.A(_16347_),
    .Z(_16349_));
 MUX2_X1 _22413_ (.A(_16311_),
    .B(\block_reg[3][19] ),
    .S(_16349_),
    .Z(_00545_));
 MUX2_X1 _22414_ (.A(_16313_),
    .B(\block_reg[3][1] ),
    .S(_16349_),
    .Z(_00546_));
 MUX2_X1 _22415_ (.A(_16314_),
    .B(\block_reg[3][20] ),
    .S(_16349_),
    .Z(_00547_));
 MUX2_X1 _22416_ (.A(_16315_),
    .B(\block_reg[3][21] ),
    .S(_16349_),
    .Z(_00548_));
 MUX2_X1 _22417_ (.A(_16316_),
    .B(\block_reg[3][22] ),
    .S(_16349_),
    .Z(_00549_));
 MUX2_X1 _22418_ (.A(_16317_),
    .B(\block_reg[3][23] ),
    .S(_16349_),
    .Z(_00550_));
 MUX2_X1 _22419_ (.A(_16318_),
    .B(\block_reg[3][24] ),
    .S(_16349_),
    .Z(_00551_));
 MUX2_X1 _22420_ (.A(_16319_),
    .B(\block_reg[3][25] ),
    .S(_16349_),
    .Z(_00552_));
 MUX2_X1 _22421_ (.A(_16320_),
    .B(\block_reg[3][26] ),
    .S(_16349_),
    .Z(_00553_));
 MUX2_X1 _22422_ (.A(_16321_),
    .B(\block_reg[3][27] ),
    .S(_16349_),
    .Z(_00554_));
 CLKBUF_X3 _22423_ (.A(_16347_),
    .Z(_16350_));
 MUX2_X1 _22424_ (.A(_16322_),
    .B(\block_reg[3][28] ),
    .S(_16350_),
    .Z(_00555_));
 MUX2_X1 _22425_ (.A(_16324_),
    .B(\block_reg[3][29] ),
    .S(_16350_),
    .Z(_00556_));
 MUX2_X1 _22426_ (.A(_16325_),
    .B(\block_reg[3][2] ),
    .S(_16350_),
    .Z(_00557_));
 MUX2_X1 _22427_ (.A(_16326_),
    .B(\block_reg[3][30] ),
    .S(_16350_),
    .Z(_00558_));
 MUX2_X1 _22428_ (.A(_16327_),
    .B(\block_reg[3][31] ),
    .S(_16350_),
    .Z(_00559_));
 MUX2_X1 _22429_ (.A(_16328_),
    .B(\block_reg[3][3] ),
    .S(_16350_),
    .Z(_00560_));
 MUX2_X1 _22430_ (.A(_16329_),
    .B(\block_reg[3][4] ),
    .S(_16350_),
    .Z(_00561_));
 MUX2_X1 _22431_ (.A(_16330_),
    .B(\block_reg[3][5] ),
    .S(_16350_),
    .Z(_00562_));
 MUX2_X1 _22432_ (.A(_16331_),
    .B(\block_reg[3][6] ),
    .S(_16350_),
    .Z(_00563_));
 MUX2_X1 _22433_ (.A(_16332_),
    .B(\block_reg[3][7] ),
    .S(_16350_),
    .Z(_00564_));
 MUX2_X1 _22434_ (.A(_16333_),
    .B(\block_reg[3][8] ),
    .S(_16347_),
    .Z(_00565_));
 MUX2_X1 _22435_ (.A(_16334_),
    .B(\block_reg[3][9] ),
    .S(_16347_),
    .Z(_00566_));
 CLKBUF_X3 _22436_ (.A(_00174_),
    .Z(_16351_));
 NAND2_X2 _22437_ (.A1(_16260_),
    .A2(_16351_),
    .ZN(_16352_));
 AOI21_X4 _22438_ (.A(_16259_),
    .B1(_16275_),
    .B2(_16352_),
    .ZN(_16353_));
 INV_X2 _22439_ (.A(_16351_),
    .ZN(_16354_));
 BUF_X4 _22440_ (.A(_22132_),
    .Z(_16355_));
 BUF_X4 _22441_ (.A(_16355_),
    .Z(_16356_));
 BUF_X4 _22442_ (.A(_16356_),
    .Z(_16357_));
 BUF_X4 _22443_ (.A(_16357_),
    .Z(_16358_));
 BUF_X4 _22444_ (.A(_16358_),
    .Z(_16359_));
 NOR2_X4 _22445_ (.A1(_16278_),
    .A2(_16260_),
    .ZN(_16360_));
 AOI21_X1 _22446_ (.A(_16354_),
    .B1(_16359_),
    .B2(_16360_),
    .ZN(_16361_));
 NOR2_X2 _22447_ (.A1(_16258_),
    .A2(_16361_),
    .ZN(_16362_));
 OR2_X1 _22448_ (.A1(_16353_),
    .A2(_16362_),
    .ZN(_16363_));
 BUF_X4 _22449_ (.A(_16363_),
    .Z(_16364_));
 CLKBUF_X3 _22450_ (.A(_16364_),
    .Z(_16365_));
 BUF_X4 _22451_ (.A(_16365_),
    .Z(_16366_));
 NOR2_X4 _22452_ (.A1(_16353_),
    .A2(_16362_),
    .ZN(_16367_));
 NOR2_X2 _22453_ (.A1(_16258_),
    .A2(_16351_),
    .ZN(_16368_));
 INV_X1 _22454_ (.A(_16368_),
    .ZN(_16369_));
 NOR2_X2 _22455_ (.A1(_16261_),
    .A2(_16369_),
    .ZN(_16370_));
 BUF_X4 _22456_ (.A(_16370_),
    .Z(_16371_));
 BUF_X4 _22457_ (.A(_16371_),
    .Z(_16372_));
 CLKBUF_X3 _22458_ (.A(\core.enc_block.round[0] ),
    .Z(_16373_));
 NAND2_X1 _22459_ (.A1(_16236_),
    .A2(_16373_),
    .ZN(_16374_));
 BUF_X4 _22460_ (.A(\core.dec_block.round[0] ),
    .Z(_16375_));
 BUF_X4 _22461_ (.A(\core.dec_block.round[1] ),
    .Z(_16376_));
 NAND2_X1 _22462_ (.A1(_16375_),
    .A2(_16376_),
    .ZN(_16377_));
 MUX2_X2 _22463_ (.A(_16374_),
    .B(_16377_),
    .S(_16262_),
    .Z(_16378_));
 NOR3_X2 _22464_ (.A1(_16202_),
    .A2(_16272_),
    .A3(_16273_),
    .ZN(_16379_));
 BUF_X4 _22465_ (.A(\core.enc_block.round[2] ),
    .Z(_16380_));
 BUF_X4 _22466_ (.A(\core.enc_block.round[3] ),
    .Z(_16381_));
 NOR2_X2 _22467_ (.A1(_16380_),
    .A2(_16381_),
    .ZN(_16382_));
 AOI21_X4 _22468_ (.A(_16379_),
    .B1(_16382_),
    .B2(_16202_),
    .ZN(_16383_));
 NOR2_X4 _22469_ (.A1(_16378_),
    .A2(_16383_),
    .ZN(_16384_));
 BUF_X8 _22470_ (.A(_16384_),
    .Z(_16385_));
 BUF_X8 _22471_ (.A(_16385_),
    .Z(_16386_));
 BUF_X4 _22472_ (.A(_16386_),
    .Z(_16387_));
 NAND2_X1 _22473_ (.A1(_16380_),
    .A2(_16381_),
    .ZN(_16388_));
 NAND2_X1 _22474_ (.A1(_16272_),
    .A2(_16273_),
    .ZN(_16389_));
 MUX2_X2 _22475_ (.A(_16388_),
    .B(_16389_),
    .S(_16262_),
    .Z(_16390_));
 NOR3_X2 _22476_ (.A1(_16202_),
    .A2(_16375_),
    .A3(_16376_),
    .ZN(_16391_));
 NOR2_X2 _22477_ (.A1(_16236_),
    .A2(_16373_),
    .ZN(_16392_));
 BUF_X4 _22478_ (.A(_16202_),
    .Z(_16393_));
 AOI21_X4 _22479_ (.A(_16391_),
    .B1(_16392_),
    .B2(_16393_),
    .ZN(_16394_));
 NOR2_X2 _22480_ (.A1(_16390_),
    .A2(_16394_),
    .ZN(_16395_));
 BUF_X4 _22481_ (.A(_16395_),
    .Z(_16396_));
 BUF_X8 _22482_ (.A(_16396_),
    .Z(_16397_));
 BUF_X8 _22483_ (.A(_16397_),
    .Z(_16398_));
 BUF_X8 _22484_ (.A(_16398_),
    .Z(_16399_));
 AOI22_X1 _22485_ (.A1(\core.keymem.key_mem[3][64] ),
    .A2(_16387_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][64] ),
    .ZN(_16400_));
 NAND2_X2 _22486_ (.A1(_16202_),
    .A2(_16380_),
    .ZN(_16401_));
 OR2_X4 _22487_ (.A1(_16381_),
    .A2(_16401_),
    .ZN(_16402_));
 INV_X1 _22488_ (.A(_16272_),
    .ZN(_16403_));
 OR3_X4 _22489_ (.A1(_16393_),
    .A2(_16403_),
    .A3(_16273_),
    .ZN(_16404_));
 AOI21_X4 _22490_ (.A(_16378_),
    .B1(_16402_),
    .B2(_16404_),
    .ZN(_16405_));
 BUF_X8 _22491_ (.A(_16405_),
    .Z(_16406_));
 BUF_X8 _22492_ (.A(_16406_),
    .Z(_16407_));
 BUF_X8 _22493_ (.A(_16407_),
    .Z(_16408_));
 INV_X2 _22494_ (.A(_16373_),
    .ZN(_16409_));
 OR3_X1 _22495_ (.A1(_16262_),
    .A2(_16236_),
    .A3(_16409_),
    .ZN(_16410_));
 BUF_X4 _22496_ (.A(_16410_),
    .Z(_16411_));
 INV_X2 _22497_ (.A(_16376_),
    .ZN(_16412_));
 NAND3_X4 _22498_ (.A1(_16262_),
    .A2(_16375_),
    .A3(_16412_),
    .ZN(_16413_));
 AOI21_X4 _22499_ (.A(_16383_),
    .B1(_16411_),
    .B2(_16413_),
    .ZN(_16414_));
 BUF_X8 _22500_ (.A(_16414_),
    .Z(_16415_));
 BUF_X8 _22501_ (.A(_16415_),
    .Z(_16416_));
 BUF_X8 _22502_ (.A(_16416_),
    .Z(_16417_));
 AOI22_X1 _22503_ (.A1(\core.keymem.key_mem[7][64] ),
    .A2(_16408_),
    .B1(_16417_),
    .B2(\core.keymem.key_mem[1][64] ),
    .ZN(_16418_));
 AND2_X1 _22504_ (.A1(_16201_),
    .A2(_16236_),
    .ZN(_16419_));
 NOR2_X1 _22505_ (.A1(_16201_),
    .A2(_16375_),
    .ZN(_16420_));
 AOI22_X4 _22506_ (.A1(_16409_),
    .A2(_16419_),
    .B1(_16420_),
    .B2(_16376_),
    .ZN(_16421_));
 NOR2_X4 _22507_ (.A1(_16383_),
    .A2(_16421_),
    .ZN(_16422_));
 BUF_X8 _22508_ (.A(_16422_),
    .Z(_16423_));
 BUF_X8 _22509_ (.A(_16423_),
    .Z(_16424_));
 BUF_X8 _22510_ (.A(_16424_),
    .Z(_16425_));
 INV_X2 _22511_ (.A(_16380_),
    .ZN(_16426_));
 NAND3_X4 _22512_ (.A1(_16393_),
    .A2(_16426_),
    .A3(_16381_),
    .ZN(_16427_));
 NOR2_X2 _22513_ (.A1(_16202_),
    .A2(_16272_),
    .ZN(_16428_));
 NAND2_X4 _22514_ (.A1(_16273_),
    .A2(_16428_),
    .ZN(_16429_));
 AOI21_X4 _22515_ (.A(_16421_),
    .B1(_16427_),
    .B2(_16429_),
    .ZN(_16430_));
 BUF_X8 _22516_ (.A(_16430_),
    .Z(_16431_));
 BUF_X8 _22517_ (.A(_16431_),
    .Z(_16432_));
 BUF_X8 _22518_ (.A(_16432_),
    .Z(_16433_));
 AOI22_X1 _22519_ (.A1(\core.keymem.key_mem[2][64] ),
    .A2(_16425_),
    .B1(_16433_),
    .B2(\core.keymem.key_mem[10][64] ),
    .ZN(_16434_));
 NOR2_X4 _22520_ (.A1(_16390_),
    .A2(_16421_),
    .ZN(_16435_));
 BUF_X8 _22521_ (.A(_16435_),
    .Z(_16436_));
 BUF_X8 _22522_ (.A(_16436_),
    .Z(_16437_));
 BUF_X8 _22523_ (.A(_16437_),
    .Z(_16438_));
 BUF_X8 _22524_ (.A(_16438_),
    .Z(_16439_));
 AOI21_X4 _22525_ (.A(_16378_),
    .B1(_16427_),
    .B2(_16429_),
    .ZN(_16440_));
 BUF_X8 _22526_ (.A(_16440_),
    .Z(_16441_));
 BUF_X8 _22527_ (.A(_16441_),
    .Z(_16442_));
 BUF_X8 _22528_ (.A(_16442_),
    .Z(_16443_));
 AOI22_X1 _22529_ (.A1(\core.keymem.key_mem[14][64] ),
    .A2(_16439_),
    .B1(_16443_),
    .B2(\core.keymem.key_mem[11][64] ),
    .ZN(_16444_));
 NAND4_X1 _22530_ (.A1(_16400_),
    .A2(_16418_),
    .A3(_16434_),
    .A4(_16444_),
    .ZN(_16445_));
 AOI21_X4 _22531_ (.A(_16421_),
    .B1(_16404_),
    .B2(_16402_),
    .ZN(_16446_));
 BUF_X8 _22532_ (.A(_16446_),
    .Z(_16447_));
 BUF_X4 _22533_ (.A(_16447_),
    .Z(_16448_));
 BUF_X8 _22534_ (.A(_16448_),
    .Z(_16449_));
 AOI21_X4 _22535_ (.A(_16394_),
    .B1(_16427_),
    .B2(_16429_),
    .ZN(_16450_));
 BUF_X8 _22536_ (.A(_16450_),
    .Z(_16451_));
 BUF_X8 _22537_ (.A(_16451_),
    .Z(_16452_));
 BUF_X8 _22538_ (.A(_16452_),
    .Z(_16453_));
 AOI22_X1 _22539_ (.A1(\core.keymem.key_mem[6][64] ),
    .A2(_16449_),
    .B1(_16453_),
    .B2(\core.keymem.key_mem[8][64] ),
    .ZN(_16454_));
 AOI21_X4 _22540_ (.A(_16394_),
    .B1(_16402_),
    .B2(_16404_),
    .ZN(_16455_));
 BUF_X8 _22541_ (.A(_16455_),
    .Z(_16456_));
 BUF_X8 _22542_ (.A(_16456_),
    .Z(_16457_));
 BUF_X8 _22543_ (.A(_16457_),
    .Z(_16458_));
 AOI22_X4 _22544_ (.A1(_16427_),
    .A2(_16429_),
    .B1(_16411_),
    .B2(_16413_),
    .ZN(_16459_));
 BUF_X4 _22545_ (.A(_16459_),
    .Z(_16460_));
 BUF_X8 _22546_ (.A(_16460_),
    .Z(_16461_));
 BUF_X8 _22547_ (.A(_16461_),
    .Z(_16462_));
 BUF_X8 _22548_ (.A(_16462_),
    .Z(_16463_));
 AOI22_X1 _22549_ (.A1(\core.keymem.key_mem[4][64] ),
    .A2(_16458_),
    .B1(_16463_),
    .B2(\core.keymem.key_mem[9][64] ),
    .ZN(_16464_));
 AOI22_X4 _22550_ (.A1(_16402_),
    .A2(_16404_),
    .B1(_16411_),
    .B2(_16413_),
    .ZN(_16465_));
 BUF_X4 _22551_ (.A(_16465_),
    .Z(_16466_));
 BUF_X8 _22552_ (.A(_16466_),
    .Z(_16467_));
 BUF_X8 _22553_ (.A(_16467_),
    .Z(_16468_));
 BUF_X8 _22554_ (.A(_16468_),
    .Z(_16469_));
 AOI21_X4 _22555_ (.A(_16390_),
    .B1(_16411_),
    .B2(_16413_),
    .ZN(_16470_));
 BUF_X8 _22556_ (.A(_16470_),
    .Z(_16471_));
 BUF_X8 _22557_ (.A(_16471_),
    .Z(_16472_));
 BUF_X8 _22558_ (.A(_16472_),
    .Z(_16473_));
 AOI22_X1 _22559_ (.A1(\core.keymem.key_mem[5][64] ),
    .A2(_16469_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][64] ),
    .ZN(_16474_));
 NAND3_X1 _22560_ (.A1(_16454_),
    .A2(_16464_),
    .A3(_16474_),
    .ZN(_16475_));
 NOR2_X1 _22561_ (.A1(_16445_),
    .A2(_16475_),
    .ZN(_16476_));
 INV_X2 _22562_ (.A(_16381_),
    .ZN(_16477_));
 OAI22_X4 _22563_ (.A1(_16477_),
    .A2(_16401_),
    .B1(_16389_),
    .B2(_16393_),
    .ZN(_16478_));
 NAND3_X1 _22564_ (.A1(_16393_),
    .A2(_16236_),
    .A3(_16373_),
    .ZN(_16479_));
 OAI21_X4 _22565_ (.A(_16479_),
    .B1(_16377_),
    .B2(_16203_),
    .ZN(_16480_));
 BUF_X4 _22566_ (.A(_16480_),
    .Z(_16481_));
 NOR2_X1 _22567_ (.A1(_16375_),
    .A2(_16376_),
    .ZN(_16482_));
 MUX2_X2 _22568_ (.A(_16482_),
    .B(_16392_),
    .S(_16393_),
    .Z(_16483_));
 BUF_X4 _22569_ (.A(_16483_),
    .Z(_16484_));
 MUX2_X2 _22570_ (.A(_16274_),
    .B(_16382_),
    .S(_16393_),
    .Z(_16485_));
 AOI22_X4 _22571_ (.A1(_16478_),
    .A2(_16481_),
    .B1(_16484_),
    .B2(_16485_),
    .ZN(_16486_));
 BUF_X8 _22572_ (.A(_16486_),
    .Z(_16487_));
 BUF_X8 _22573_ (.A(_16487_),
    .Z(_16488_));
 BUF_X8 _22574_ (.A(_16488_),
    .Z(_16489_));
 MUX2_X2 _22575_ (.A(_00225_),
    .B(_16476_),
    .S(_16489_),
    .Z(_16490_));
 XNOR2_X1 _22576_ (.A(\block_reg[1][0] ),
    .B(_16490_),
    .ZN(_16491_));
 AOI21_X1 _22577_ (.A(_16367_),
    .B1(_16372_),
    .B2(_16491_),
    .ZN(_16492_));
 OAI22_X4 _22578_ (.A1(_16390_),
    .A2(_16378_),
    .B1(_16394_),
    .B2(_16383_),
    .ZN(_16493_));
 BUF_X8 _22579_ (.A(_16493_),
    .Z(_16494_));
 BUF_X8 _22580_ (.A(_16494_),
    .Z(_16495_));
 BUF_X8 _22581_ (.A(_16495_),
    .Z(_16496_));
 BUF_X8 _22582_ (.A(_16496_),
    .Z(_16497_));
 BUF_X8 _22583_ (.A(_16497_),
    .Z(_16498_));
 BUF_X8 _22584_ (.A(_16455_),
    .Z(_16499_));
 BUF_X8 _22585_ (.A(_16499_),
    .Z(_16500_));
 BUF_X8 _22586_ (.A(_16500_),
    .Z(_16501_));
 BUF_X8 _22587_ (.A(_16438_),
    .Z(_16502_));
 AOI22_X2 _22588_ (.A1(\core.keymem.key_mem[4][96] ),
    .A2(_16501_),
    .B1(_16502_),
    .B2(\core.keymem.key_mem[14][96] ),
    .ZN(_16503_));
 BUF_X8 _22589_ (.A(_16440_),
    .Z(_16504_));
 BUF_X8 _22590_ (.A(_16504_),
    .Z(_16505_));
 BUF_X8 _22591_ (.A(_16505_),
    .Z(_16506_));
 BUF_X8 _22592_ (.A(_16506_),
    .Z(_16507_));
 AOI22_X2 _22593_ (.A1(\core.keymem.key_mem[2][96] ),
    .A2(_16425_),
    .B1(_16507_),
    .B2(\core.keymem.key_mem[11][96] ),
    .ZN(_16508_));
 BUF_X8 _22594_ (.A(_16467_),
    .Z(_16509_));
 BUF_X8 _22595_ (.A(_16509_),
    .Z(_16510_));
 AOI22_X2 _22596_ (.A1(\core.keymem.key_mem[3][96] ),
    .A2(_16387_),
    .B1(_16510_),
    .B2(\core.keymem.key_mem[5][96] ),
    .ZN(_16511_));
 BUF_X8 _22597_ (.A(_16406_),
    .Z(_16512_));
 BUF_X8 _22598_ (.A(_16512_),
    .Z(_16513_));
 BUF_X8 _22599_ (.A(_16430_),
    .Z(_16514_));
 BUF_X8 _22600_ (.A(_16514_),
    .Z(_16515_));
 BUF_X8 _22601_ (.A(_16515_),
    .Z(_16516_));
 AOI22_X2 _22602_ (.A1(\core.keymem.key_mem[7][96] ),
    .A2(_16513_),
    .B1(_16516_),
    .B2(\core.keymem.key_mem[10][96] ),
    .ZN(_16517_));
 NAND4_X2 _22603_ (.A1(_16503_),
    .A2(_16508_),
    .A3(_16511_),
    .A4(_16517_),
    .ZN(_16518_));
 BUF_X8 _22604_ (.A(_16446_),
    .Z(_16519_));
 BUF_X8 _22605_ (.A(_16519_),
    .Z(_16520_));
 BUF_X4 _22606_ (.A(_16520_),
    .Z(_16521_));
 BUF_X8 _22607_ (.A(_16521_),
    .Z(_16522_));
 BUF_X4 _22608_ (.A(_16414_),
    .Z(_16523_));
 BUF_X8 _22609_ (.A(_16523_),
    .Z(_16524_));
 BUF_X4 _22610_ (.A(_16524_),
    .Z(_16525_));
 BUF_X8 _22611_ (.A(_16525_),
    .Z(_16526_));
 AOI22_X1 _22612_ (.A1(\core.keymem.key_mem[6][96] ),
    .A2(_16522_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][96] ),
    .ZN(_16527_));
 BUF_X8 _22613_ (.A(_16450_),
    .Z(_16528_));
 BUF_X8 _22614_ (.A(_16528_),
    .Z(_16529_));
 BUF_X8 _22615_ (.A(_16529_),
    .Z(_16530_));
 BUF_X8 _22616_ (.A(_16470_),
    .Z(_16531_));
 BUF_X8 _22617_ (.A(_16531_),
    .Z(_16532_));
 BUF_X8 _22618_ (.A(_16532_),
    .Z(_16533_));
 AOI22_X2 _22619_ (.A1(\core.keymem.key_mem[8][96] ),
    .A2(_16530_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][96] ),
    .ZN(_16534_));
 BUF_X8 _22620_ (.A(_16460_),
    .Z(_16535_));
 BUF_X8 _22621_ (.A(_16535_),
    .Z(_16536_));
 BUF_X8 _22622_ (.A(_16536_),
    .Z(_16537_));
 BUF_X8 _22623_ (.A(_16396_),
    .Z(_16538_));
 BUF_X8 _22624_ (.A(_16538_),
    .Z(_16539_));
 BUF_X8 _22625_ (.A(_16539_),
    .Z(_16540_));
 AOI22_X2 _22626_ (.A1(\core.keymem.key_mem[9][96] ),
    .A2(_16537_),
    .B1(_16540_),
    .B2(\core.keymem.key_mem[12][96] ),
    .ZN(_16541_));
 NAND3_X2 _22627_ (.A1(_16527_),
    .A2(_16534_),
    .A3(_16541_),
    .ZN(_16542_));
 NOR3_X4 _22628_ (.A1(_16498_),
    .A2(_16518_),
    .A3(_16542_),
    .ZN(_16543_));
 BUF_X8 _22629_ (.A(_16493_),
    .Z(_16544_));
 BUF_X8 _22630_ (.A(_16544_),
    .Z(_16545_));
 BUF_X8 _22631_ (.A(_16545_),
    .Z(_16546_));
 BUF_X8 _22632_ (.A(_16546_),
    .Z(_16547_));
 BUF_X8 _22633_ (.A(_16547_),
    .Z(_16548_));
 BUF_X8 _22634_ (.A(_16548_),
    .Z(_16549_));
 AOI21_X4 _22635_ (.A(_16543_),
    .B1(_16549_),
    .B2(_00186_),
    .ZN(_16550_));
 XNOR2_X2 _22636_ (.A(\core.dec_block.block_w0_reg[0] ),
    .B(_16550_),
    .ZN(_16551_));
 NAND2_X1 _22637_ (.A1(_22128_),
    .A2(_16274_),
    .ZN(_16552_));
 OR3_X2 _22638_ (.A1(_16259_),
    .A2(_16552_),
    .A3(_16352_),
    .ZN(_16553_));
 BUF_X4 _22639_ (.A(_16553_),
    .Z(_16554_));
 BUF_X4 _22640_ (.A(_16554_),
    .Z(_16555_));
 BUF_X4 _22641_ (.A(_16555_),
    .Z(_16556_));
 OAI21_X1 _22642_ (.A(_16492_),
    .B1(_16551_),
    .B2(_16556_),
    .ZN(_16557_));
 NOR4_X4 _22643_ (.A1(_16258_),
    .A2(_16278_),
    .A3(_00324_),
    .A4(_16354_),
    .ZN(_16558_));
 BUF_X8 _22644_ (.A(_16558_),
    .Z(_16559_));
 BUF_X4 _22645_ (.A(_16559_),
    .Z(_16560_));
 BUF_X4 _22646_ (.A(_16560_),
    .Z(_16561_));
 BUF_X4 _22647_ (.A(_16561_),
    .Z(_16562_));
 NAND2_X1 _22648_ (.A1(_16358_),
    .A2(\core.dec_block.block_w0_reg[2] ),
    .ZN(_16563_));
 BUF_X4 _22649_ (.A(_22134_),
    .Z(_16564_));
 BUF_X4 _22650_ (.A(_16564_),
    .Z(_16565_));
 BUF_X4 _22651_ (.A(_16565_),
    .Z(_16566_));
 BUF_X4 _22652_ (.A(_22136_),
    .Z(_16567_));
 BUF_X4 _22653_ (.A(_16567_),
    .Z(_16568_));
 BUF_X4 _22654_ (.A(_16568_),
    .Z(_16569_));
 AOI222_X2 _22655_ (.A1(\core.dec_block.block_w2_reg[2] ),
    .A2(_16566_),
    .B1(_16569_),
    .B2(\core.dec_block.block_w1_reg[2] ),
    .C1(_16267_),
    .C2(\core.dec_block.block_w3_reg[2] ),
    .ZN(_16570_));
 OAI21_X4 _22656_ (.A(_16563_),
    .B1(_16570_),
    .B2(_16358_),
    .ZN(_16571_));
 NAND2_X1 _22657_ (.A1(_16358_),
    .A2(\core.dec_block.block_w0_reg[3] ),
    .ZN(_16572_));
 AOI222_X2 _22658_ (.A1(\core.dec_block.block_w2_reg[3] ),
    .A2(_16566_),
    .B1(_16569_),
    .B2(\core.dec_block.block_w1_reg[3] ),
    .C1(_16267_),
    .C2(\core.dec_block.block_w3_reg[3] ),
    .ZN(_16573_));
 OAI21_X4 _22659_ (.A(_16572_),
    .B1(_16573_),
    .B2(_16358_),
    .ZN(_16574_));
 OAI21_X4 _22660_ (.A(_16562_),
    .B1(_16571_),
    .B2(_16574_),
    .ZN(_16575_));
 BUF_X4 _22661_ (.A(_16560_),
    .Z(_16576_));
 NAND2_X1 _22662_ (.A1(_16358_),
    .A2(\core.dec_block.block_w0_reg[1] ),
    .ZN(_16577_));
 AOI222_X2 _22663_ (.A1(\core.dec_block.block_w2_reg[1] ),
    .A2(_16566_),
    .B1(_16569_),
    .B2(\core.dec_block.block_w1_reg[1] ),
    .C1(_16267_),
    .C2(\core.dec_block.block_w3_reg[1] ),
    .ZN(_16578_));
 OAI21_X2 _22664_ (.A(_16577_),
    .B1(_16578_),
    .B2(_16358_),
    .ZN(_16579_));
 AND2_X2 _22665_ (.A1(_16576_),
    .A2(_16579_),
    .ZN(_16580_));
 BUF_X2 _22666_ (.A(\core.dec_block.block_w0_reg[7] ),
    .Z(_16581_));
 NAND2_X1 _22667_ (.A1(_16581_),
    .A2(_16357_),
    .ZN(_16582_));
 AOI222_X2 _22668_ (.A1(\core.dec_block.block_w2_reg[7] ),
    .A2(_16566_),
    .B1(_16569_),
    .B2(\core.dec_block.block_w1_reg[7] ),
    .C1(_16266_),
    .C2(\core.dec_block.block_w3_reg[7] ),
    .ZN(_16583_));
 BUF_X4 _22669_ (.A(_16356_),
    .Z(_16584_));
 OAI21_X2 _22670_ (.A(_16582_),
    .B1(_16583_),
    .B2(_16584_),
    .ZN(_16585_));
 NAND2_X2 _22671_ (.A1(_16561_),
    .A2(_16585_),
    .ZN(_16586_));
 BUF_X4 _22672_ (.A(_16586_),
    .Z(_16587_));
 NAND2_X1 _22673_ (.A1(\core.dec_block.block_w0_reg[6] ),
    .A2(_16356_),
    .ZN(_16588_));
 BUF_X2 _22674_ (.A(\core.dec_block.block_w2_reg[6] ),
    .Z(_16589_));
 AOI222_X2 _22675_ (.A1(_16589_),
    .A2(_16565_),
    .B1(_16568_),
    .B2(\core.dec_block.block_w1_reg[6] ),
    .C1(_16266_),
    .C2(\core.dec_block.block_w3_reg[6] ),
    .ZN(_16590_));
 OAI21_X4 _22676_ (.A(_16588_),
    .B1(_16590_),
    .B2(_16357_),
    .ZN(_16591_));
 NAND2_X4 _22677_ (.A1(_16576_),
    .A2(_16591_),
    .ZN(_16592_));
 NAND2_X4 _22678_ (.A1(_16587_),
    .A2(_16592_),
    .ZN(_16593_));
 NAND2_X1 _22679_ (.A1(\core.dec_block.block_w0_reg[5] ),
    .A2(_16357_),
    .ZN(_16594_));
 AOI222_X2 _22680_ (.A1(\core.dec_block.block_w2_reg[5] ),
    .A2(_16565_),
    .B1(_16568_),
    .B2(\core.dec_block.block_w1_reg[5] ),
    .C1(_16266_),
    .C2(\core.dec_block.block_w3_reg[5] ),
    .ZN(_16595_));
 OAI21_X4 _22681_ (.A(_16594_),
    .B1(_16595_),
    .B2(_16584_),
    .ZN(_16596_));
 AND2_X2 _22682_ (.A1(_16561_),
    .A2(_16596_),
    .ZN(_16597_));
 NAND2_X1 _22683_ (.A1(_16356_),
    .A2(\core.dec_block.block_w0_reg[4] ),
    .ZN(_16598_));
 AOI222_X2 _22684_ (.A1(\core.dec_block.block_w2_reg[4] ),
    .A2(_16565_),
    .B1(_16568_),
    .B2(\core.dec_block.block_w1_reg[4] ),
    .C1(_16266_),
    .C2(\core.dec_block.block_w3_reg[4] ),
    .ZN(_16599_));
 OAI21_X4 _22685_ (.A(_16598_),
    .B1(_16599_),
    .B2(_16356_),
    .ZN(_16600_));
 NAND2_X4 _22686_ (.A1(_16561_),
    .A2(_16600_),
    .ZN(_16601_));
 NAND2_X4 _22687_ (.A1(_16597_),
    .A2(_16601_),
    .ZN(_16602_));
 NOR2_X4 _22688_ (.A1(_16593_),
    .A2(_16602_),
    .ZN(_16603_));
 NAND2_X1 _22689_ (.A1(_16580_),
    .A2(_16603_),
    .ZN(_16604_));
 AND2_X1 _22690_ (.A1(_16576_),
    .A2(_16574_),
    .ZN(_16605_));
 BUF_X4 _22691_ (.A(_16605_),
    .Z(_16606_));
 AND2_X1 _22692_ (.A1(_16560_),
    .A2(_16600_),
    .ZN(_16607_));
 BUF_X4 _22693_ (.A(_16607_),
    .Z(_16608_));
 NAND2_X4 _22694_ (.A1(_16597_),
    .A2(_16608_),
    .ZN(_16609_));
 AND2_X1 _22695_ (.A1(_16560_),
    .A2(_16591_),
    .ZN(_16610_));
 BUF_X4 _22696_ (.A(_16610_),
    .Z(_16611_));
 NAND2_X4 _22697_ (.A1(_16586_),
    .A2(_16611_),
    .ZN(_16612_));
 NOR2_X4 _22698_ (.A1(_16609_),
    .A2(_16612_),
    .ZN(_16613_));
 AND2_X2 _22699_ (.A1(_16562_),
    .A2(_16571_),
    .ZN(_16614_));
 OAI21_X1 _22700_ (.A(_16606_),
    .B1(_16613_),
    .B2(_16614_),
    .ZN(_16615_));
 AND2_X1 _22701_ (.A1(_16576_),
    .A2(_16585_),
    .ZN(_16616_));
 BUF_X4 _22702_ (.A(_16616_),
    .Z(_16617_));
 NOR2_X2 _22703_ (.A1(_16617_),
    .A2(_16611_),
    .ZN(_16618_));
 NAND2_X4 _22704_ (.A1(_16576_),
    .A2(_16596_),
    .ZN(_16619_));
 NOR2_X4 _22705_ (.A1(_16619_),
    .A2(_16601_),
    .ZN(_16620_));
 NAND2_X1 _22706_ (.A1(_16618_),
    .A2(_16620_),
    .ZN(_16621_));
 BUF_X4 _22707_ (.A(_16576_),
    .Z(_16622_));
 NAND2_X4 _22708_ (.A1(_16622_),
    .A2(_16571_),
    .ZN(_16623_));
 NAND2_X4 _22709_ (.A1(_16562_),
    .A2(_16574_),
    .ZN(_16624_));
 BUF_X4 _22710_ (.A(_16624_),
    .Z(_16625_));
 NOR2_X4 _22711_ (.A1(_16623_),
    .A2(_16625_),
    .ZN(_16626_));
 AOI221_X2 _22712_ (.A(_16575_),
    .B1(_16604_),
    .B2(_16615_),
    .C1(_16621_),
    .C2(_16626_),
    .ZN(_16627_));
 NOR2_X4 _22713_ (.A1(_16619_),
    .A2(_16608_),
    .ZN(_16628_));
 NOR2_X4 _22714_ (.A1(_16587_),
    .A2(_16592_),
    .ZN(_16629_));
 NAND2_X2 _22715_ (.A1(_16628_),
    .A2(_16629_),
    .ZN(_16630_));
 NAND2_X4 _22716_ (.A1(_16620_),
    .A2(_16629_),
    .ZN(_16631_));
 BUF_X4 _22717_ (.A(_16580_),
    .Z(_16632_));
 OAI21_X1 _22718_ (.A(_16630_),
    .B1(_16631_),
    .B2(_16632_),
    .ZN(_16633_));
 BUF_X4 _22719_ (.A(_16625_),
    .Z(_16634_));
 BUF_X4 _22720_ (.A(_16614_),
    .Z(_16635_));
 BUF_X4 _22721_ (.A(_16619_),
    .Z(_16636_));
 NAND2_X4 _22722_ (.A1(_16636_),
    .A2(_16608_),
    .ZN(_16637_));
 NOR2_X4 _22723_ (.A1(_16593_),
    .A2(_16637_),
    .ZN(_16638_));
 NAND2_X1 _22724_ (.A1(_16635_),
    .A2(_16638_),
    .ZN(_16639_));
 NAND2_X1 _22725_ (.A1(\core.dec_block.block_w0_reg[0] ),
    .A2(_16584_),
    .ZN(_16640_));
 AOI222_X2 _22726_ (.A1(\core.dec_block.block_w2_reg[0] ),
    .A2(_16566_),
    .B1(_16569_),
    .B2(\core.dec_block.block_w1_reg[0] ),
    .C1(_16267_),
    .C2(\core.dec_block.block_w3_reg[0] ),
    .ZN(_16641_));
 OAI21_X2 _22727_ (.A(_16640_),
    .B1(_16641_),
    .B2(_16584_),
    .ZN(_16642_));
 AND2_X1 _22728_ (.A1(_16561_),
    .A2(_16642_),
    .ZN(_16643_));
 BUF_X4 _22729_ (.A(_16643_),
    .Z(_16644_));
 NAND2_X1 _22730_ (.A1(_16576_),
    .A2(_16579_),
    .ZN(_16645_));
 BUF_X4 _22731_ (.A(_16645_),
    .Z(_16646_));
 NAND2_X4 _22732_ (.A1(_16644_),
    .A2(_16646_),
    .ZN(_16647_));
 BUF_X4 _22733_ (.A(_16623_),
    .Z(_16648_));
 NAND2_X4 _22734_ (.A1(_16636_),
    .A2(_16601_),
    .ZN(_16649_));
 NOR2_X4 _22735_ (.A1(_16593_),
    .A2(_16649_),
    .ZN(_16650_));
 NAND2_X1 _22736_ (.A1(_16648_),
    .A2(_16650_),
    .ZN(_16651_));
 OAI21_X1 _22737_ (.A(_16639_),
    .B1(_16647_),
    .B2(_16651_),
    .ZN(_16652_));
 AOI221_X2 _22738_ (.A(_16627_),
    .B1(_16633_),
    .B2(_16626_),
    .C1(_16634_),
    .C2(_16652_),
    .ZN(_16653_));
 BUF_X4 _22739_ (.A(_16635_),
    .Z(_16654_));
 CLKBUF_X3 _22740_ (.A(_16654_),
    .Z(_16655_));
 BUF_X4 _22741_ (.A(_16625_),
    .Z(_16656_));
 BUF_X4 _22742_ (.A(_16592_),
    .Z(_16657_));
 NAND2_X4 _22743_ (.A1(_16617_),
    .A2(_16657_),
    .ZN(_16658_));
 NOR2_X4 _22744_ (.A1(_16602_),
    .A2(_16658_),
    .ZN(_16659_));
 NAND2_X1 _22745_ (.A1(_16656_),
    .A2(_16659_),
    .ZN(_16660_));
 NOR2_X4 _22746_ (.A1(_16597_),
    .A2(_16608_),
    .ZN(_16661_));
 NAND2_X2 _22747_ (.A1(_16618_),
    .A2(_16661_),
    .ZN(_16662_));
 BUF_X4 _22748_ (.A(_16662_),
    .Z(_16663_));
 BUF_X4 _22749_ (.A(_16656_),
    .Z(_16664_));
 OAI21_X1 _22750_ (.A(_16660_),
    .B1(_16663_),
    .B2(_16664_),
    .ZN(_16665_));
 NOR2_X4 _22751_ (.A1(_16635_),
    .A2(_16624_),
    .ZN(_16666_));
 BUF_X4 _22752_ (.A(_16644_),
    .Z(_16667_));
 BUF_X4 _22753_ (.A(_16601_),
    .Z(_16668_));
 BUF_X4 _22754_ (.A(_16611_),
    .Z(_16669_));
 BUF_X4 _22755_ (.A(_16597_),
    .Z(_16670_));
 NOR3_X4 _22756_ (.A1(_16587_),
    .A2(_16669_),
    .A3(_16670_),
    .ZN(_16671_));
 NAND2_X2 _22757_ (.A1(_16668_),
    .A2(_16671_),
    .ZN(_16672_));
 NOR2_X1 _22758_ (.A1(_16667_),
    .A2(_16672_),
    .ZN(_16673_));
 AOI22_X1 _22759_ (.A1(_16655_),
    .A2(_16665_),
    .B1(_16666_),
    .B2(_16673_),
    .ZN(_16674_));
 BUF_X4 _22760_ (.A(_16646_),
    .Z(_16675_));
 BUF_X4 _22761_ (.A(_16675_),
    .Z(_16676_));
 CLKBUF_X3 _22762_ (.A(_16676_),
    .Z(_16677_));
 CLKBUF_X3 _22763_ (.A(_16677_),
    .Z(_16678_));
 NOR2_X4 _22764_ (.A1(_16617_),
    .A2(_16657_),
    .ZN(_16679_));
 NAND2_X4 _22765_ (.A1(_16620_),
    .A2(_16679_),
    .ZN(_16680_));
 NAND2_X4 _22766_ (.A1(_16614_),
    .A2(_16606_),
    .ZN(_16681_));
 BUF_X4 _22767_ (.A(_16681_),
    .Z(_16682_));
 NOR2_X4 _22768_ (.A1(_16670_),
    .A2(_16668_),
    .ZN(_16683_));
 NAND2_X1 _22769_ (.A1(_16618_),
    .A2(_16683_),
    .ZN(_16684_));
 BUF_X4 _22770_ (.A(_16684_),
    .Z(_16685_));
 BUF_X4 _22771_ (.A(_16575_),
    .Z(_16686_));
 NAND2_X1 _22772_ (.A1(_16644_),
    .A2(_16686_),
    .ZN(_16687_));
 OAI22_X1 _22773_ (.A1(_16680_),
    .A2(_16682_),
    .B1(_16685_),
    .B2(_16687_),
    .ZN(_16688_));
 NAND2_X4 _22774_ (.A1(_16576_),
    .A2(_16642_),
    .ZN(_16689_));
 NAND2_X1 _22775_ (.A1(_16689_),
    .A2(_16646_),
    .ZN(_16690_));
 CLKBUF_X3 _22776_ (.A(_16690_),
    .Z(_16691_));
 NAND2_X4 _22777_ (.A1(_16623_),
    .A2(_16625_),
    .ZN(_16692_));
 NAND2_X1 _22778_ (.A1(_16683_),
    .A2(_16629_),
    .ZN(_16693_));
 BUF_X4 _22779_ (.A(_16693_),
    .Z(_16694_));
 NOR2_X1 _22780_ (.A1(_16692_),
    .A2(_16694_),
    .ZN(_16695_));
 AOI22_X1 _22781_ (.A1(_16678_),
    .A2(_16688_),
    .B1(_16691_),
    .B2(_16695_),
    .ZN(_16696_));
 NAND2_X1 _22782_ (.A1(_16674_),
    .A2(_16696_),
    .ZN(_16697_));
 BUF_X4 _22783_ (.A(_16606_),
    .Z(_16698_));
 NAND2_X4 _22784_ (.A1(_16628_),
    .A2(_16679_),
    .ZN(_16699_));
 NAND2_X2 _22785_ (.A1(_16689_),
    .A2(_16632_),
    .ZN(_16700_));
 CLKBUF_X3 _22786_ (.A(_16700_),
    .Z(_16701_));
 NOR3_X1 _22787_ (.A1(_16698_),
    .A2(_16699_),
    .A3(_16701_),
    .ZN(_16702_));
 NAND2_X4 _22788_ (.A1(_16623_),
    .A2(_16606_),
    .ZN(_16703_));
 NOR2_X4 _22789_ (.A1(_16703_),
    .A2(_16700_),
    .ZN(_16704_));
 BUF_X4 _22790_ (.A(_16632_),
    .Z(_16705_));
 NOR2_X2 _22791_ (.A1(_16705_),
    .A2(_16692_),
    .ZN(_16706_));
 NAND2_X4 _22792_ (.A1(_16617_),
    .A2(_16611_),
    .ZN(_16707_));
 NOR2_X4 _22793_ (.A1(_16609_),
    .A2(_16707_),
    .ZN(_16708_));
 AOI221_X2 _22794_ (.A(_16702_),
    .B1(_16704_),
    .B2(_16638_),
    .C1(_16706_),
    .C2(_16708_),
    .ZN(_16709_));
 NAND2_X4 _22795_ (.A1(_16647_),
    .A2(_16700_),
    .ZN(_16710_));
 NAND2_X1 _22796_ (.A1(_16664_),
    .A2(_16710_),
    .ZN(_16711_));
 NOR2_X4 _22797_ (.A1(_16649_),
    .A2(_16707_),
    .ZN(_16712_));
 NAND2_X2 _22798_ (.A1(_16654_),
    .A2(_16712_),
    .ZN(_16713_));
 CLKBUF_X3 _22799_ (.A(_16664_),
    .Z(_16714_));
 BUF_X4 _22800_ (.A(_16648_),
    .Z(_16715_));
 NOR2_X2 _22801_ (.A1(_16602_),
    .A2(_16707_),
    .ZN(_16716_));
 BUF_X4 _22802_ (.A(_16716_),
    .Z(_16717_));
 NAND2_X1 _22803_ (.A1(_16715_),
    .A2(_16717_),
    .ZN(_16718_));
 MUX2_X1 _22804_ (.A(_16713_),
    .B(_16718_),
    .S(_16710_),
    .Z(_16719_));
 OAI221_X2 _22805_ (.A(_16709_),
    .B1(_16711_),
    .B2(_16713_),
    .C1(_16714_),
    .C2(_16719_),
    .ZN(_16720_));
 NOR2_X1 _22806_ (.A1(_16697_),
    .A2(_16720_),
    .ZN(_16721_));
 BUF_X4 _22807_ (.A(_16689_),
    .Z(_16722_));
 NOR2_X2 _22808_ (.A1(_16635_),
    .A2(_16722_),
    .ZN(_16723_));
 NAND2_X1 _22809_ (.A1(_16618_),
    .A2(_16628_),
    .ZN(_16724_));
 BUF_X4 _22810_ (.A(_16724_),
    .Z(_16725_));
 NAND2_X2 _22811_ (.A1(_16625_),
    .A2(_16675_),
    .ZN(_16726_));
 NAND2_X2 _22812_ (.A1(_16698_),
    .A2(_16632_),
    .ZN(_16727_));
 NAND2_X4 _22813_ (.A1(_16661_),
    .A2(_16629_),
    .ZN(_16728_));
 OAI22_X1 _22814_ (.A1(_16725_),
    .A2(_16726_),
    .B1(_16727_),
    .B2(_16728_),
    .ZN(_16729_));
 NAND2_X1 _22815_ (.A1(_16723_),
    .A2(_16729_),
    .ZN(_16730_));
 NAND2_X1 _22816_ (.A1(_16626_),
    .A2(_16710_),
    .ZN(_16731_));
 NAND2_X4 _22817_ (.A1(_16679_),
    .A2(_16683_),
    .ZN(_16732_));
 BUF_X4 _22818_ (.A(_16626_),
    .Z(_16733_));
 AOI22_X1 _22819_ (.A1(_16733_),
    .A2(_16638_),
    .B1(_16686_),
    .B2(_16717_),
    .ZN(_16734_));
 OAI221_X2 _22820_ (.A(_16730_),
    .B1(_16731_),
    .B2(_16732_),
    .C1(_16734_),
    .C2(_16678_),
    .ZN(_16735_));
 BUF_X4 _22821_ (.A(_16703_),
    .Z(_16736_));
 BUF_X4 _22822_ (.A(_16722_),
    .Z(_16737_));
 BUF_X4 _22823_ (.A(_16621_),
    .Z(_16738_));
 AOI21_X1 _22824_ (.A(_16737_),
    .B1(_16738_),
    .B2(_16732_),
    .ZN(_16739_));
 NOR2_X4 _22825_ (.A1(_16689_),
    .A2(_16580_),
    .ZN(_16740_));
 NOR2_X4 _22826_ (.A1(_16644_),
    .A2(_16646_),
    .ZN(_16741_));
 NOR2_X2 _22827_ (.A1(_16740_),
    .A2(_16741_),
    .ZN(_16742_));
 NOR2_X4 _22828_ (.A1(_16602_),
    .A2(_16612_),
    .ZN(_16743_));
 AOI21_X1 _22829_ (.A(_16739_),
    .B1(_16742_),
    .B2(_16743_),
    .ZN(_16744_));
 CLKBUF_X3 _22830_ (.A(_16705_),
    .Z(_16745_));
 NOR2_X4 _22831_ (.A1(_16637_),
    .A2(_16707_),
    .ZN(_16746_));
 NOR2_X4 _22832_ (.A1(_16658_),
    .A2(_16609_),
    .ZN(_16747_));
 AOI21_X1 _22833_ (.A(_16746_),
    .B1(_16747_),
    .B2(_16667_),
    .ZN(_16748_));
 NOR2_X1 _22834_ (.A1(_16745_),
    .A2(_16748_),
    .ZN(_16749_));
 NOR2_X1 _22835_ (.A1(_16722_),
    .A2(_16672_),
    .ZN(_16750_));
 AOI21_X1 _22836_ (.A(_16749_),
    .B1(_16750_),
    .B2(_16745_),
    .ZN(_16751_));
 OAI22_X2 _22837_ (.A1(_16736_),
    .A2(_16744_),
    .B1(_16751_),
    .B2(_16682_),
    .ZN(_16752_));
 BUF_X4 _22838_ (.A(_16648_),
    .Z(_16753_));
 BUF_X4 _22839_ (.A(_16698_),
    .Z(_16754_));
 OAI22_X1 _22840_ (.A1(_16663_),
    .A2(_16667_),
    .B1(_16631_),
    .B2(_16741_),
    .ZN(_16755_));
 NAND3_X1 _22841_ (.A1(_16753_),
    .A2(_16754_),
    .A3(_16755_),
    .ZN(_16756_));
 AND2_X1 _22842_ (.A1(_16580_),
    .A2(_16575_),
    .ZN(_16757_));
 BUF_X4 _22843_ (.A(_16757_),
    .Z(_16758_));
 NAND2_X4 _22844_ (.A1(_16689_),
    .A2(_16758_),
    .ZN(_16759_));
 NOR2_X4 _22845_ (.A1(_16612_),
    .A2(_16637_),
    .ZN(_16760_));
 NOR2_X4 _22846_ (.A1(_16689_),
    .A2(_16646_),
    .ZN(_16761_));
 OAI21_X1 _22847_ (.A(_16691_),
    .B1(_16761_),
    .B2(_16698_),
    .ZN(_16762_));
 NOR2_X2 _22848_ (.A1(_16722_),
    .A2(_16680_),
    .ZN(_16763_));
 BUF_X4 _22849_ (.A(_16675_),
    .Z(_16764_));
 NOR2_X1 _22850_ (.A1(_16634_),
    .A2(_16764_),
    .ZN(_16765_));
 AOI22_X1 _22851_ (.A1(_16760_),
    .A2(_16762_),
    .B1(_16763_),
    .B2(_16765_),
    .ZN(_16766_));
 BUF_X4 _22852_ (.A(_16753_),
    .Z(_16767_));
 OAI221_X2 _22853_ (.A(_16756_),
    .B1(_16759_),
    .B2(_16685_),
    .C1(_16766_),
    .C2(_16767_),
    .ZN(_16768_));
 NAND3_X4 _22854_ (.A1(_16617_),
    .A2(_16657_),
    .A3(_16636_),
    .ZN(_16769_));
 CLKBUF_X3 _22855_ (.A(_16668_),
    .Z(_16770_));
 NOR3_X1 _22856_ (.A1(_16770_),
    .A2(_16703_),
    .A3(_16742_),
    .ZN(_16771_));
 AND2_X1 _22857_ (.A1(_16722_),
    .A2(_16758_),
    .ZN(_16772_));
 AOI21_X2 _22858_ (.A(_16771_),
    .B1(_16772_),
    .B2(_16770_),
    .ZN(_16773_));
 MUX2_X1 _22859_ (.A(_16693_),
    .B(_16728_),
    .S(_16648_),
    .Z(_16774_));
 BUF_X4 _22860_ (.A(_16644_),
    .Z(_16775_));
 NAND2_X1 _22861_ (.A1(_16775_),
    .A2(_16712_),
    .ZN(_16776_));
 MUX2_X1 _22862_ (.A(_16774_),
    .B(_16776_),
    .S(_16705_),
    .Z(_16777_));
 OAI22_X4 _22863_ (.A1(_16769_),
    .A2(_16773_),
    .B1(_16777_),
    .B2(_16754_),
    .ZN(_16778_));
 NOR4_X2 _22864_ (.A1(_16735_),
    .A2(_16752_),
    .A3(_16768_),
    .A4(_16778_),
    .ZN(_16779_));
 NAND3_X2 _22865_ (.A1(_16653_),
    .A2(_16721_),
    .A3(_16779_),
    .ZN(_16780_));
 NAND2_X2 _22866_ (.A1(_16666_),
    .A2(_16646_),
    .ZN(_16781_));
 NOR2_X4 _22867_ (.A1(_16623_),
    .A2(_16606_),
    .ZN(_16782_));
 NAND2_X1 _22868_ (.A1(_16761_),
    .A2(_16782_),
    .ZN(_16783_));
 AOI21_X1 _22869_ (.A(_16694_),
    .B1(_16781_),
    .B2(_16783_),
    .ZN(_16784_));
 NAND2_X4 _22870_ (.A1(_16614_),
    .A2(_16624_),
    .ZN(_16785_));
 AOI22_X1 _22871_ (.A1(_16708_),
    .A2(_16740_),
    .B1(_16741_),
    .B2(_16716_),
    .ZN(_16786_));
 NOR2_X1 _22872_ (.A1(_16785_),
    .A2(_16786_),
    .ZN(_16787_));
 OR2_X1 _22873_ (.A1(_16784_),
    .A2(_16787_),
    .ZN(_16788_));
 NOR2_X1 _22874_ (.A1(_16649_),
    .A2(_16612_),
    .ZN(_16789_));
 CLKBUF_X3 _22875_ (.A(_16789_),
    .Z(_16790_));
 NAND2_X1 _22876_ (.A1(_16654_),
    .A2(_16790_),
    .ZN(_16791_));
 OR2_X1 _22877_ (.A1(_16602_),
    .A2(_16658_),
    .ZN(_16792_));
 CLKBUF_X3 _22878_ (.A(_16792_),
    .Z(_16793_));
 BUF_X4 _22879_ (.A(_16654_),
    .Z(_16794_));
 OAI21_X1 _22880_ (.A(_16791_),
    .B1(_16793_),
    .B2(_16794_),
    .ZN(_16795_));
 CLKBUF_X3 _22881_ (.A(_16632_),
    .Z(_16796_));
 NOR2_X1 _22882_ (.A1(_16656_),
    .A2(_16796_),
    .ZN(_16797_));
 BUF_X4 _22883_ (.A(_16775_),
    .Z(_16798_));
 BUF_X4 _22884_ (.A(_16798_),
    .Z(_16799_));
 NAND2_X4 _22885_ (.A1(_16646_),
    .A2(_16782_),
    .ZN(_16800_));
 OAI22_X2 _22886_ (.A1(_16736_),
    .A2(_16694_),
    .B1(_16800_),
    .B2(_16680_),
    .ZN(_16801_));
 AOI221_X2 _22887_ (.A(_16788_),
    .B1(_16795_),
    .B2(_16797_),
    .C1(_16799_),
    .C2(_16801_),
    .ZN(_16802_));
 BUF_X4 _22888_ (.A(_16796_),
    .Z(_16803_));
 AOI21_X2 _22889_ (.A(_16769_),
    .B1(_16803_),
    .B2(_16770_),
    .ZN(_16804_));
 NOR2_X2 _22890_ (.A1(_16775_),
    .A2(_16680_),
    .ZN(_16805_));
 AOI21_X2 _22891_ (.A(_16804_),
    .B1(_16805_),
    .B2(_16803_),
    .ZN(_16806_));
 OAI21_X4 _22892_ (.A(_16802_),
    .B1(_16806_),
    .B2(_16785_),
    .ZN(_16807_));
 CLKBUF_X3 _22893_ (.A(_16617_),
    .Z(_16808_));
 NAND3_X1 _22894_ (.A1(_16808_),
    .A2(_16657_),
    .A3(_16798_),
    .ZN(_16809_));
 CLKBUF_X3 _22895_ (.A(_16669_),
    .Z(_16810_));
 BUF_X4 _22896_ (.A(_16737_),
    .Z(_16811_));
 NAND3_X1 _22897_ (.A1(_16587_),
    .A2(_16810_),
    .A3(_16811_),
    .ZN(_16812_));
 AOI21_X1 _22898_ (.A(_16602_),
    .B1(_16809_),
    .B2(_16812_),
    .ZN(_16813_));
 NOR3_X1 _22899_ (.A1(_16770_),
    .A2(_16811_),
    .A3(_16707_),
    .ZN(_16814_));
 OAI21_X1 _22900_ (.A(_16803_),
    .B1(_16813_),
    .B2(_16814_),
    .ZN(_16815_));
 NAND2_X1 _22901_ (.A1(_16587_),
    .A2(_16668_),
    .ZN(_16816_));
 NAND2_X1 _22902_ (.A1(_16611_),
    .A2(_16670_),
    .ZN(_16817_));
 OR3_X1 _22903_ (.A1(_16647_),
    .A2(_16816_),
    .A3(_16817_),
    .ZN(_16818_));
 AOI21_X2 _22904_ (.A(_16682_),
    .B1(_16815_),
    .B2(_16818_),
    .ZN(_16819_));
 NAND2_X1 _22905_ (.A1(_16745_),
    .A2(_16613_),
    .ZN(_16820_));
 BUF_X4 _22906_ (.A(_16608_),
    .Z(_16821_));
 NOR2_X2 _22907_ (.A1(_16821_),
    .A2(_16769_),
    .ZN(_16822_));
 NAND2_X2 _22908_ (.A1(_16822_),
    .A2(_16764_),
    .ZN(_16823_));
 AOI21_X1 _22909_ (.A(_16687_),
    .B1(_16820_),
    .B2(_16823_),
    .ZN(_16824_));
 NOR2_X4 _22910_ (.A1(_16644_),
    .A2(_16632_),
    .ZN(_16825_));
 NAND2_X2 _22911_ (.A1(_16666_),
    .A2(_16825_),
    .ZN(_16826_));
 NOR2_X1 _22912_ (.A1(_16728_),
    .A2(_16826_),
    .ZN(_16827_));
 NOR2_X4 _22913_ (.A1(_16593_),
    .A2(_16609_),
    .ZN(_16828_));
 AOI21_X1 _22914_ (.A(_16827_),
    .B1(_16772_),
    .B2(_16828_),
    .ZN(_16829_));
 NOR2_X1 _22915_ (.A1(_16682_),
    .A2(_16701_),
    .ZN(_16830_));
 NOR2_X4 _22916_ (.A1(_16668_),
    .A2(_16769_),
    .ZN(_16831_));
 OAI21_X1 _22917_ (.A(_16830_),
    .B1(_16831_),
    .B2(_16603_),
    .ZN(_16832_));
 NAND2_X1 _22918_ (.A1(_16829_),
    .A2(_16832_),
    .ZN(_16833_));
 BUF_X4 _22919_ (.A(_16754_),
    .Z(_16834_));
 XNOR2_X2 _22920_ (.A(_16654_),
    .B(_16775_),
    .ZN(_16835_));
 NOR4_X2 _22921_ (.A1(_16834_),
    .A2(_16663_),
    .A3(_16676_),
    .A4(_16835_),
    .ZN(_16836_));
 NOR3_X2 _22922_ (.A1(_16824_),
    .A2(_16833_),
    .A3(_16836_),
    .ZN(_16837_));
 OAI21_X1 _22923_ (.A(_16793_),
    .B1(_16672_),
    .B2(_16677_),
    .ZN(_16838_));
 NAND3_X1 _22924_ (.A1(_16686_),
    .A2(_16701_),
    .A3(_16838_),
    .ZN(_16839_));
 NAND2_X1 _22925_ (.A1(_16753_),
    .A2(_16747_),
    .ZN(_16840_));
 NAND2_X4 _22926_ (.A1(_16821_),
    .A2(_16671_),
    .ZN(_16841_));
 OAI21_X1 _22927_ (.A(_16840_),
    .B1(_16841_),
    .B2(_16753_),
    .ZN(_16842_));
 NAND3_X1 _22928_ (.A1(_16834_),
    .A2(_16740_),
    .A3(_16842_),
    .ZN(_16843_));
 OR2_X2 _22929_ (.A1(_16658_),
    .A2(_16609_),
    .ZN(_16844_));
 BUF_X4 _22930_ (.A(_16844_),
    .Z(_16845_));
 NAND2_X1 _22931_ (.A1(_16654_),
    .A2(_16676_),
    .ZN(_16846_));
 BUF_X4 _22932_ (.A(_16737_),
    .Z(_16847_));
 OAI33_X1 _22933_ (.A1(_16677_),
    .A2(_16845_),
    .A3(_16835_),
    .B1(_16846_),
    .B2(_16738_),
    .B3(_16847_),
    .ZN(_16848_));
 NAND2_X1 _22934_ (.A1(_16714_),
    .A2(_16848_),
    .ZN(_16849_));
 NAND4_X2 _22935_ (.A1(_16837_),
    .A2(_16839_),
    .A3(_16843_),
    .A4(_16849_),
    .ZN(_16850_));
 NOR4_X4 _22936_ (.A1(_16780_),
    .A2(_16807_),
    .A3(_16819_),
    .A4(_16850_),
    .ZN(_16851_));
 BUF_X8 _22937_ (.A(_16546_),
    .Z(_16852_));
 AOI22_X2 _22938_ (.A1(\core.keymem.key_mem[12][70] ),
    .A2(_16539_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][70] ),
    .ZN(_16853_));
 BUF_X8 _22939_ (.A(_16523_),
    .Z(_16854_));
 BUF_X8 _22940_ (.A(_16854_),
    .Z(_16855_));
 AOI22_X2 _22941_ (.A1(\core.keymem.key_mem[6][70] ),
    .A2(_16448_),
    .B1(_16855_),
    .B2(\core.keymem.key_mem[1][70] ),
    .ZN(_16856_));
 AOI22_X2 _22942_ (.A1(\core.keymem.key_mem[14][70] ),
    .A2(_16438_),
    .B1(_16512_),
    .B2(\core.keymem.key_mem[7][70] ),
    .ZN(_16857_));
 BUF_X8 _22943_ (.A(_16422_),
    .Z(_16858_));
 BUF_X8 _22944_ (.A(_16858_),
    .Z(_16859_));
 BUF_X8 _22945_ (.A(_16859_),
    .Z(_16860_));
 AOI22_X2 _22946_ (.A1(\core.keymem.key_mem[2][70] ),
    .A2(_16860_),
    .B1(_16452_),
    .B2(\core.keymem.key_mem[8][70] ),
    .ZN(_16861_));
 NAND4_X2 _22947_ (.A1(_16853_),
    .A2(_16856_),
    .A3(_16857_),
    .A4(_16861_),
    .ZN(_16862_));
 AOI22_X1 _22948_ (.A1(\core.keymem.key_mem[9][70] ),
    .A2(_16536_),
    .B1(_16515_),
    .B2(\core.keymem.key_mem[10][70] ),
    .ZN(_16863_));
 BUF_X8 _22949_ (.A(_16384_),
    .Z(_16864_));
 BUF_X8 _22950_ (.A(_16864_),
    .Z(_16865_));
 BUF_X8 _22951_ (.A(_16865_),
    .Z(_16866_));
 AOI22_X2 _22952_ (.A1(\core.keymem.key_mem[3][70] ),
    .A2(_16866_),
    .B1(_16532_),
    .B2(\core.keymem.key_mem[13][70] ),
    .ZN(_16867_));
 AOI22_X2 _22953_ (.A1(\core.keymem.key_mem[4][70] ),
    .A2(_16457_),
    .B1(_16442_),
    .B2(\core.keymem.key_mem[11][70] ),
    .ZN(_16868_));
 NAND3_X2 _22954_ (.A1(_16863_),
    .A2(_16867_),
    .A3(_16868_),
    .ZN(_16869_));
 NOR3_X4 _22955_ (.A1(_16852_),
    .A2(_16862_),
    .A3(_16869_),
    .ZN(_16870_));
 BUF_X8 _22956_ (.A(_16545_),
    .Z(_16871_));
 BUF_X8 _22957_ (.A(_16871_),
    .Z(_16872_));
 BUF_X8 _22958_ (.A(_16872_),
    .Z(_16873_));
 AOI21_X4 _22959_ (.A(_16870_),
    .B1(_16873_),
    .B2(_00232_),
    .ZN(_16874_));
 XNOR2_X2 _22960_ (.A(\core.dec_block.block_w1_reg[6] ),
    .B(_16874_),
    .ZN(_16875_));
 INV_X1 _22961_ (.A(\core.dec_block.block_w1_reg[21] ),
    .ZN(_16876_));
 NOR3_X4 _22962_ (.A1(_16262_),
    .A2(_16236_),
    .A3(_16409_),
    .ZN(_16877_));
 INV_X2 _22963_ (.A(_16375_),
    .ZN(_16878_));
 NOR3_X4 _22964_ (.A1(_16393_),
    .A2(_16878_),
    .A3(_16376_),
    .ZN(_16879_));
 NOR2_X4 _22965_ (.A1(_16877_),
    .A2(_16879_),
    .ZN(_16880_));
 BUF_X4 _22966_ (.A(_16478_),
    .Z(_16881_));
 BUF_X4 _22967_ (.A(_16881_),
    .Z(_16882_));
 NAND2_X1 _22968_ (.A1(\core.keymem.key_mem[13][85] ),
    .A2(_16882_),
    .ZN(_16883_));
 NOR3_X4 _22969_ (.A1(_16262_),
    .A2(_16380_),
    .A3(_16477_),
    .ZN(_16884_));
 BUF_X4 _22970_ (.A(_16884_),
    .Z(_16885_));
 BUF_X4 _22971_ (.A(_16885_),
    .Z(_16886_));
 AND2_X1 _22972_ (.A1(_16273_),
    .A2(_16428_),
    .ZN(_16887_));
 BUF_X4 _22973_ (.A(_16887_),
    .Z(_16888_));
 BUF_X4 _22974_ (.A(_16888_),
    .Z(_16889_));
 BUF_X4 _22975_ (.A(_16889_),
    .Z(_16890_));
 OAI21_X1 _22976_ (.A(\core.keymem.key_mem[9][85] ),
    .B1(_16886_),
    .B2(_16890_),
    .ZN(_16891_));
 AOI21_X2 _22977_ (.A(_16880_),
    .B1(_16883_),
    .B2(_16891_),
    .ZN(_16892_));
 BUF_X4 _22978_ (.A(_16484_),
    .Z(_16893_));
 NOR2_X2 _22979_ (.A1(_16381_),
    .A2(_16401_),
    .ZN(_16894_));
 BUF_X4 _22980_ (.A(_16894_),
    .Z(_16895_));
 BUF_X4 _22981_ (.A(_16895_),
    .Z(_16896_));
 NOR3_X2 _22982_ (.A1(_16203_),
    .A2(_16403_),
    .A3(_16273_),
    .ZN(_16897_));
 BUF_X4 _22983_ (.A(_16897_),
    .Z(_16898_));
 BUF_X4 _22984_ (.A(_16898_),
    .Z(_16899_));
 OAI211_X2 _22985_ (.A(\core.keymem.key_mem[4][85] ),
    .B(_16893_),
    .C1(_16896_),
    .C2(_16899_),
    .ZN(_16900_));
 BUF_X4 _22986_ (.A(_16481_),
    .Z(_16901_));
 BUF_X4 _22987_ (.A(_16485_),
    .Z(_16902_));
 NAND3_X1 _22988_ (.A1(\core.keymem.key_mem[3][85] ),
    .A2(_16901_),
    .A3(_16902_),
    .ZN(_16903_));
 NAND2_X1 _22989_ (.A1(_16393_),
    .A2(_16236_),
    .ZN(_16904_));
 OR2_X1 _22990_ (.A1(_16202_),
    .A2(_16375_),
    .ZN(_16905_));
 OAI22_X4 _22991_ (.A1(_16373_),
    .A2(_16904_),
    .B1(_16905_),
    .B2(_16412_),
    .ZN(_16906_));
 BUF_X4 _22992_ (.A(_16906_),
    .Z(_16907_));
 BUF_X4 _22993_ (.A(_16895_),
    .Z(_16908_));
 OAI211_X2 _22994_ (.A(\core.keymem.key_mem[6][85] ),
    .B(_16907_),
    .C1(_16899_),
    .C2(_16908_),
    .ZN(_16909_));
 NAND3_X1 _22995_ (.A1(\core.keymem.key_mem[2][85] ),
    .A2(_16902_),
    .A3(_16907_),
    .ZN(_16910_));
 NAND4_X2 _22996_ (.A1(_16900_),
    .A2(_16903_),
    .A3(_16909_),
    .A4(_16910_),
    .ZN(_16911_));
 BUF_X4 _22997_ (.A(_16877_),
    .Z(_16912_));
 BUF_X4 _22998_ (.A(_16912_),
    .Z(_16913_));
 BUF_X4 _22999_ (.A(_16879_),
    .Z(_16914_));
 BUF_X4 _23000_ (.A(_16914_),
    .Z(_16915_));
 OAI211_X2 _23001_ (.A(\core.keymem.key_mem[1][85] ),
    .B(_16902_),
    .C1(_16913_),
    .C2(_16915_),
    .ZN(_16916_));
 BUF_X4 _23002_ (.A(_16898_),
    .Z(_16917_));
 OAI211_X2 _23003_ (.A(\core.keymem.key_mem[7][85] ),
    .B(_16901_),
    .C1(_16908_),
    .C2(_16917_),
    .ZN(_16918_));
 BUF_X4 _23004_ (.A(_16881_),
    .Z(_16919_));
 NAND3_X1 _23005_ (.A1(\core.keymem.key_mem[14][85] ),
    .A2(_16919_),
    .A3(_16907_),
    .ZN(_16920_));
 BUF_X4 _23006_ (.A(_16484_),
    .Z(_16921_));
 BUF_X4 _23007_ (.A(_16884_),
    .Z(_16922_));
 BUF_X4 _23008_ (.A(_16888_),
    .Z(_16923_));
 OAI211_X2 _23009_ (.A(\core.keymem.key_mem[8][85] ),
    .B(_16921_),
    .C1(_16922_),
    .C2(_16923_),
    .ZN(_16924_));
 NAND4_X2 _23010_ (.A1(_16916_),
    .A2(_16918_),
    .A3(_16920_),
    .A4(_16924_),
    .ZN(_16925_));
 BUF_X4 _23011_ (.A(_16884_),
    .Z(_16926_));
 BUF_X4 _23012_ (.A(_16926_),
    .Z(_16927_));
 BUF_X4 _23013_ (.A(_16888_),
    .Z(_16928_));
 BUF_X4 _23014_ (.A(_16928_),
    .Z(_16929_));
 OAI211_X2 _23015_ (.A(\core.keymem.key_mem[10][85] ),
    .B(_16907_),
    .C1(_16927_),
    .C2(_16929_),
    .ZN(_16930_));
 BUF_X4 _23016_ (.A(_16484_),
    .Z(_16931_));
 NAND3_X1 _23017_ (.A1(\core.keymem.key_mem[12][85] ),
    .A2(_16919_),
    .A3(_16931_),
    .ZN(_16932_));
 BUF_X4 _23018_ (.A(_16894_),
    .Z(_16933_));
 BUF_X4 _23019_ (.A(_16898_),
    .Z(_16934_));
 BUF_X4 _23020_ (.A(_16912_),
    .Z(_16935_));
 BUF_X4 _23021_ (.A(_16914_),
    .Z(_16936_));
 OAI221_X2 _23022_ (.A(\core.keymem.key_mem[5][85] ),
    .B1(_16933_),
    .B2(_16934_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_16937_));
 BUF_X4 _23023_ (.A(_16480_),
    .Z(_16938_));
 OAI211_X2 _23024_ (.A(\core.keymem.key_mem[11][85] ),
    .B(_16938_),
    .C1(_16922_),
    .C2(_16923_),
    .ZN(_16939_));
 NAND4_X2 _23025_ (.A1(_16930_),
    .A2(_16932_),
    .A3(_16937_),
    .A4(_16939_),
    .ZN(_16940_));
 NOR4_X4 _23026_ (.A1(_16892_),
    .A2(_16911_),
    .A3(_16925_),
    .A4(_16940_),
    .ZN(_16941_));
 MUX2_X2 _23027_ (.A(_00218_),
    .B(_16941_),
    .S(_16487_),
    .Z(_16942_));
 XNOR2_X2 _23028_ (.A(_16876_),
    .B(_16942_),
    .ZN(_16943_));
 INV_X1 _23029_ (.A(\core.dec_block.block_w1_reg[22] ),
    .ZN(_16944_));
 NAND2_X1 _23030_ (.A1(_00230_),
    .A2(_16547_),
    .ZN(_16945_));
 BUF_X8 _23031_ (.A(_16455_),
    .Z(_16946_));
 BUF_X8 _23032_ (.A(_16946_),
    .Z(_16947_));
 BUF_X8 _23033_ (.A(_16465_),
    .Z(_16948_));
 BUF_X8 _23034_ (.A(_16948_),
    .Z(_16949_));
 AOI22_X1 _23035_ (.A1(\core.keymem.key_mem[4][86] ),
    .A2(_16947_),
    .B1(_16949_),
    .B2(\core.keymem.key_mem[5][86] ),
    .ZN(_16950_));
 AOI22_X1 _23036_ (.A1(\core.keymem.key_mem[10][86] ),
    .A2(_16432_),
    .B1(_16442_),
    .B2(\core.keymem.key_mem[11][86] ),
    .ZN(_16951_));
 AOI22_X1 _23037_ (.A1(\core.keymem.key_mem[9][86] ),
    .A2(_16462_),
    .B1(_16398_),
    .B2(\core.keymem.key_mem[12][86] ),
    .ZN(_16952_));
 NAND3_X1 _23038_ (.A1(_16950_),
    .A2(_16951_),
    .A3(_16952_),
    .ZN(_16953_));
 BUF_X4 _23039_ (.A(_16405_),
    .Z(_16954_));
 BUF_X8 _23040_ (.A(_16954_),
    .Z(_16955_));
 AOI222_X2 _23041_ (.A1(\core.keymem.key_mem[7][86] ),
    .A2(_16955_),
    .B1(_16385_),
    .B2(\core.keymem.key_mem[3][86] ),
    .C1(_16415_),
    .C2(\core.keymem.key_mem[1][86] ),
    .ZN(_16956_));
 MUX2_X1 _23042_ (.A(_16403_),
    .B(_16426_),
    .S(_16203_),
    .Z(_16957_));
 BUF_X4 _23043_ (.A(_16957_),
    .Z(_16958_));
 AND3_X1 _23044_ (.A1(\core.keymem.key_mem[8][86] ),
    .A2(_16921_),
    .A3(_16958_),
    .ZN(_16959_));
 MUX2_X2 _23045_ (.A(_16272_),
    .B(_16380_),
    .S(_16393_),
    .Z(_16960_));
 BUF_X4 _23046_ (.A(_16960_),
    .Z(_16961_));
 AND2_X1 _23047_ (.A1(\core.keymem.key_mem[13][86] ),
    .A2(_16961_),
    .ZN(_16962_));
 NAND2_X2 _23048_ (.A1(_16411_),
    .A2(_16413_),
    .ZN(_16963_));
 BUF_X4 _23049_ (.A(_16963_),
    .Z(_16964_));
 AOI21_X1 _23050_ (.A(_16959_),
    .B1(_16962_),
    .B2(_16964_),
    .ZN(_16965_));
 AND2_X1 _23051_ (.A1(_16202_),
    .A2(_16381_),
    .ZN(_16966_));
 AOI21_X4 _23052_ (.A(_16966_),
    .B1(_16273_),
    .B2(_16262_),
    .ZN(_16967_));
 BUF_X8 _23053_ (.A(_16421_),
    .Z(_16968_));
 BUF_X4 _23054_ (.A(_16485_),
    .Z(_16969_));
 BUF_X4 _23055_ (.A(_16969_),
    .Z(_16970_));
 MUX2_X1 _23056_ (.A(_16273_),
    .B(_16381_),
    .S(_16202_),
    .Z(_16971_));
 BUF_X4 _23057_ (.A(_16971_),
    .Z(_16972_));
 MUX2_X1 _23058_ (.A(\core.keymem.key_mem[6][86] ),
    .B(\core.keymem.key_mem[14][86] ),
    .S(_16972_),
    .Z(_16973_));
 AOI22_X2 _23059_ (.A1(\core.keymem.key_mem[2][86] ),
    .A2(_16970_),
    .B1(_16961_),
    .B2(_16973_),
    .ZN(_16974_));
 OAI221_X2 _23060_ (.A(_16956_),
    .B1(_16965_),
    .B2(_16967_),
    .C1(_16968_),
    .C2(_16974_),
    .ZN(_16975_));
 OR2_X1 _23061_ (.A1(_16953_),
    .A2(_16975_),
    .ZN(_16976_));
 OAI21_X4 _23062_ (.A(_16945_),
    .B1(_16976_),
    .B2(_16547_),
    .ZN(_16977_));
 XNOR2_X2 _23063_ (.A(_16944_),
    .B(_16977_),
    .ZN(_16978_));
 XNOR2_X2 _23064_ (.A(_16943_),
    .B(_16978_),
    .ZN(_16979_));
 XNOR2_X1 _23065_ (.A(_16875_),
    .B(_16979_),
    .ZN(_16980_));
 INV_X1 _23066_ (.A(\core.dec_block.block_w1_reg[8] ),
    .ZN(_16981_));
 BUF_X8 _23067_ (.A(_16494_),
    .Z(_16982_));
 BUF_X8 _23068_ (.A(_16982_),
    .Z(_16983_));
 BUF_X8 _23069_ (.A(_16983_),
    .Z(_16984_));
 NAND2_X1 _23070_ (.A1(_00226_),
    .A2(_16984_),
    .ZN(_16985_));
 BUF_X8 _23071_ (.A(_16864_),
    .Z(_16986_));
 BUF_X8 _23072_ (.A(_16986_),
    .Z(_16987_));
 BUF_X8 _23073_ (.A(_16431_),
    .Z(_16988_));
 BUF_X8 _23074_ (.A(_16988_),
    .Z(_16989_));
 AOI222_X2 _23075_ (.A1(\core.keymem.key_mem[3][72] ),
    .A2(_16987_),
    .B1(_16989_),
    .B2(\core.keymem.key_mem[10][72] ),
    .C1(\core.keymem.key_mem[13][72] ),
    .C2(_16532_),
    .ZN(_16990_));
 BUF_X8 _23076_ (.A(_16520_),
    .Z(_16991_));
 AOI22_X2 _23077_ (.A1(\core.keymem.key_mem[6][72] ),
    .A2(_16991_),
    .B1(_16453_),
    .B2(\core.keymem.key_mem[8][72] ),
    .ZN(_16992_));
 BUF_X8 _23078_ (.A(_16858_),
    .Z(_16993_));
 BUF_X8 _23079_ (.A(_16993_),
    .Z(_16994_));
 AOI22_X2 _23080_ (.A1(\core.keymem.key_mem[2][72] ),
    .A2(_16994_),
    .B1(_16463_),
    .B2(\core.keymem.key_mem[9][72] ),
    .ZN(_16995_));
 NAND3_X2 _23081_ (.A1(_16990_),
    .A2(_16992_),
    .A3(_16995_),
    .ZN(_16996_));
 AOI21_X1 _23082_ (.A(_16871_),
    .B1(_16408_),
    .B2(\core.keymem.key_mem[7][72] ),
    .ZN(_16997_));
 BUF_X8 _23083_ (.A(_16436_),
    .Z(_16998_));
 BUF_X8 _23084_ (.A(_16998_),
    .Z(_16999_));
 BUF_X8 _23085_ (.A(_16396_),
    .Z(_17000_));
 BUF_X8 _23086_ (.A(_17000_),
    .Z(_17001_));
 AOI22_X2 _23087_ (.A1(\core.keymem.key_mem[14][72] ),
    .A2(_16999_),
    .B1(_17001_),
    .B2(\core.keymem.key_mem[12][72] ),
    .ZN(_17002_));
 BUF_X8 _23088_ (.A(_16416_),
    .Z(_17003_));
 BUF_X4 _23089_ (.A(_16948_),
    .Z(_17004_));
 BUF_X8 _23090_ (.A(_17004_),
    .Z(_17005_));
 AOI22_X2 _23091_ (.A1(\core.keymem.key_mem[1][72] ),
    .A2(_17003_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][72] ),
    .ZN(_17006_));
 BUF_X8 _23092_ (.A(_16504_),
    .Z(_17007_));
 BUF_X8 _23093_ (.A(_17007_),
    .Z(_17008_));
 AOI22_X2 _23094_ (.A1(\core.keymem.key_mem[4][72] ),
    .A2(_16500_),
    .B1(_17008_),
    .B2(\core.keymem.key_mem[11][72] ),
    .ZN(_17009_));
 NAND4_X2 _23095_ (.A1(_16997_),
    .A2(_17002_),
    .A3(_17006_),
    .A4(_17009_),
    .ZN(_17010_));
 OAI21_X4 _23096_ (.A(_16985_),
    .B1(_16996_),
    .B2(_17010_),
    .ZN(_17011_));
 XNOR2_X2 _23097_ (.A(_16981_),
    .B(_17011_),
    .ZN(_17012_));
 BUF_X8 _23098_ (.A(_16545_),
    .Z(_17013_));
 BUF_X8 _23099_ (.A(_17013_),
    .Z(_17014_));
 BUF_X4 _23100_ (.A(_16906_),
    .Z(_17015_));
 BUF_X4 _23101_ (.A(_17015_),
    .Z(_17016_));
 NAND2_X1 _23102_ (.A1(\core.keymem.key_mem[2][77] ),
    .A2(_17016_),
    .ZN(_17017_));
 BUF_X4 _23103_ (.A(_16877_),
    .Z(_17018_));
 BUF_X4 _23104_ (.A(_17018_),
    .Z(_17019_));
 BUF_X4 _23105_ (.A(_16879_),
    .Z(_17020_));
 BUF_X4 _23106_ (.A(_17020_),
    .Z(_17021_));
 OAI21_X1 _23107_ (.A(\core.keymem.key_mem[1][77] ),
    .B1(_17019_),
    .B2(_17021_),
    .ZN(_17022_));
 AOI21_X2 _23108_ (.A(_16383_),
    .B1(_17017_),
    .B2(_17022_),
    .ZN(_17023_));
 BUF_X4 _23109_ (.A(_16881_),
    .Z(_17024_));
 BUF_X4 _23110_ (.A(_16906_),
    .Z(_17025_));
 BUF_X4 _23111_ (.A(_17025_),
    .Z(_17026_));
 NAND3_X1 _23112_ (.A1(\core.keymem.key_mem[14][77] ),
    .A2(_17024_),
    .A3(_17026_),
    .ZN(_17027_));
 BUF_X4 _23113_ (.A(_16921_),
    .Z(_17028_));
 OAI211_X2 _23114_ (.A(\core.keymem.key_mem[8][77] ),
    .B(_17028_),
    .C1(_16886_),
    .C2(_16890_),
    .ZN(_17029_));
 BUF_X4 _23115_ (.A(_16933_),
    .Z(_17030_));
 BUF_X4 _23116_ (.A(_16934_),
    .Z(_17031_));
 OAI211_X2 _23117_ (.A(\core.keymem.key_mem[4][77] ),
    .B(_17028_),
    .C1(_17030_),
    .C2(_17031_),
    .ZN(_17032_));
 NAND4_X2 _23118_ (.A1(_16487_),
    .A2(_17027_),
    .A3(_17029_),
    .A4(_17032_),
    .ZN(_17033_));
 INV_X1 _23119_ (.A(\core.keymem.key_mem[9][77] ),
    .ZN(_17034_));
 BUF_X4 _23120_ (.A(_16926_),
    .Z(_17035_));
 BUF_X4 _23121_ (.A(_16928_),
    .Z(_17036_));
 OAI22_X2 _23122_ (.A1(_17035_),
    .A2(_17036_),
    .B1(_16913_),
    .B2(_16915_),
    .ZN(_17037_));
 OAI21_X4 _23123_ (.A(_17015_),
    .B1(_16885_),
    .B2(_16889_),
    .ZN(_17038_));
 INV_X1 _23124_ (.A(\core.keymem.key_mem[10][77] ),
    .ZN(_17039_));
 OAI22_X2 _23125_ (.A1(_17034_),
    .A2(_17037_),
    .B1(_17038_),
    .B2(_17039_),
    .ZN(_17040_));
 INV_X1 _23126_ (.A(\core.keymem.key_mem[7][77] ),
    .ZN(_17041_));
 NOR2_X4 _23127_ (.A1(_16895_),
    .A2(_16898_),
    .ZN(_17042_));
 BUF_X4 _23128_ (.A(_16958_),
    .Z(_17043_));
 AND2_X1 _23129_ (.A1(\core.keymem.key_mem[13][77] ),
    .A2(_16972_),
    .ZN(_17044_));
 AOI21_X1 _23130_ (.A(_17044_),
    .B1(_16967_),
    .B2(\core.keymem.key_mem[5][77] ),
    .ZN(_17045_));
 OAI33_X1 _23131_ (.A1(_17041_),
    .A2(_16378_),
    .A3(_17042_),
    .B1(_16880_),
    .B2(_17043_),
    .B3(_17045_),
    .ZN(_17046_));
 NOR4_X4 _23132_ (.A1(_17023_),
    .A2(_17033_),
    .A3(_17040_),
    .A4(_17046_),
    .ZN(_17047_));
 BUF_X4 _23133_ (.A(_16938_),
    .Z(_17048_));
 NAND3_X1 _23134_ (.A1(\core.keymem.key_mem[3][77] ),
    .A2(_17048_),
    .A3(_17043_),
    .ZN(_17049_));
 BUF_X4 _23135_ (.A(_16907_),
    .Z(_17050_));
 BUF_X8 _23136_ (.A(_16961_),
    .Z(_17051_));
 NAND3_X1 _23137_ (.A1(\core.keymem.key_mem[6][77] ),
    .A2(_17050_),
    .A3(_17051_),
    .ZN(_17052_));
 NAND3_X1 _23138_ (.A1(_16967_),
    .A2(_17049_),
    .A3(_17052_),
    .ZN(_17053_));
 BUF_X8 _23139_ (.A(_16972_),
    .Z(_17054_));
 BUF_X8 _23140_ (.A(_17054_),
    .Z(_17055_));
 NAND3_X1 _23141_ (.A1(\core.keymem.key_mem[11][77] ),
    .A2(_17048_),
    .A3(_17043_),
    .ZN(_17056_));
 BUF_X4 _23142_ (.A(_16893_),
    .Z(_17057_));
 NAND3_X1 _23143_ (.A1(\core.keymem.key_mem[12][77] ),
    .A2(_17057_),
    .A3(_17051_),
    .ZN(_17058_));
 NAND3_X1 _23144_ (.A1(_17055_),
    .A2(_17056_),
    .A3(_17058_),
    .ZN(_17059_));
 NAND2_X2 _23145_ (.A1(_17053_),
    .A2(_17059_),
    .ZN(_17060_));
 AOI22_X4 _23146_ (.A1(_00220_),
    .A2(_17014_),
    .B1(_17047_),
    .B2(_17060_),
    .ZN(_17061_));
 XNOR2_X2 _23147_ (.A(\core.dec_block.block_w1_reg[13] ),
    .B(_17061_),
    .ZN(_17062_));
 XNOR2_X2 _23148_ (.A(_17012_),
    .B(_17062_),
    .ZN(_17063_));
 XNOR2_X1 _23149_ (.A(_16980_),
    .B(_17063_),
    .ZN(_17064_));
 INV_X1 _23150_ (.A(\core.dec_block.block_w1_reg[29] ),
    .ZN(_17065_));
 AOI22_X1 _23151_ (.A1(\core.keymem.key_mem[2][93] ),
    .A2(_16859_),
    .B1(_16528_),
    .B2(\core.keymem.key_mem[8][93] ),
    .ZN(_17066_));
 NAND2_X4 _23152_ (.A1(_16427_),
    .A2(_16429_),
    .ZN(_17067_));
 AOI22_X2 _23153_ (.A1(\core.keymem.key_mem[14][93] ),
    .A2(_16882_),
    .B1(_17067_),
    .B2(\core.keymem.key_mem[10][93] ),
    .ZN(_17068_));
 OAI21_X1 _23154_ (.A(_17066_),
    .B1(_17068_),
    .B2(_16968_),
    .ZN(_17069_));
 AOI22_X1 _23155_ (.A1(\core.keymem.key_mem[9][93] ),
    .A2(_16535_),
    .B1(_16531_),
    .B2(\core.keymem.key_mem[13][93] ),
    .ZN(_17070_));
 AOI22_X1 _23156_ (.A1(\core.keymem.key_mem[4][93] ),
    .A2(_16456_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][93] ),
    .ZN(_17071_));
 NAND2_X1 _23157_ (.A1(_17070_),
    .A2(_17071_),
    .ZN(_17072_));
 AOI222_X2 _23158_ (.A1(\core.keymem.key_mem[3][93] ),
    .A2(_16385_),
    .B1(_16415_),
    .B2(\core.keymem.key_mem[1][93] ),
    .C1(_16504_),
    .C2(\core.keymem.key_mem[11][93] ),
    .ZN(_17073_));
 BUF_X4 _23159_ (.A(_16481_),
    .Z(_17074_));
 AOI222_X2 _23160_ (.A1(\core.keymem.key_mem[7][93] ),
    .A2(_17074_),
    .B1(_16907_),
    .B2(\core.keymem.key_mem[6][93] ),
    .C1(_16964_),
    .C2(\core.keymem.key_mem[5][93] ),
    .ZN(_17075_));
 OAI21_X1 _23161_ (.A(_17073_),
    .B1(_17075_),
    .B2(_17042_),
    .ZN(_17076_));
 NOR3_X2 _23162_ (.A1(_17069_),
    .A2(_17072_),
    .A3(_17076_),
    .ZN(_17077_));
 MUX2_X2 _23163_ (.A(_00215_),
    .B(_17077_),
    .S(_16488_),
    .Z(_17078_));
 XNOR2_X2 _23164_ (.A(_17065_),
    .B(_17078_),
    .ZN(_17079_));
 NAND2_X1 _23165_ (.A1(_00217_),
    .A2(_16548_),
    .ZN(_17080_));
 AOI222_X2 _23166_ (.A1(\core.keymem.key_mem[14][88] ),
    .A2(_16502_),
    .B1(_16537_),
    .B2(\core.keymem.key_mem[9][88] ),
    .C1(\core.keymem.key_mem[4][88] ),
    .C2(_16458_),
    .ZN(_17081_));
 BUF_X8 _23167_ (.A(_16433_),
    .Z(_17082_));
 AOI22_X2 _23168_ (.A1(\core.keymem.key_mem[10][88] ),
    .A2(_17082_),
    .B1(_16510_),
    .B2(\core.keymem.key_mem[5][88] ),
    .ZN(_17083_));
 BUF_X8 _23169_ (.A(_16955_),
    .Z(_17084_));
 BUF_X8 _23170_ (.A(_17084_),
    .Z(_17085_));
 BUF_X8 _23171_ (.A(_16994_),
    .Z(_17086_));
 AOI22_X2 _23172_ (.A1(\core.keymem.key_mem[7][88] ),
    .A2(_17085_),
    .B1(_17086_),
    .B2(\core.keymem.key_mem[2][88] ),
    .ZN(_17087_));
 NAND3_X2 _23173_ (.A1(_17081_),
    .A2(_17083_),
    .A3(_17087_),
    .ZN(_17088_));
 AOI21_X1 _23174_ (.A(_16852_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][88] ),
    .ZN(_17089_));
 AOI22_X2 _23175_ (.A1(\core.keymem.key_mem[6][88] ),
    .A2(_16522_),
    .B1(_16507_),
    .B2(\core.keymem.key_mem[11][88] ),
    .ZN(_17090_));
 BUF_X8 _23176_ (.A(_16987_),
    .Z(_17091_));
 AOI22_X2 _23177_ (.A1(\core.keymem.key_mem[8][88] ),
    .A2(_16530_),
    .B1(_17091_),
    .B2(\core.keymem.key_mem[3][88] ),
    .ZN(_17092_));
 BUF_X8 _23178_ (.A(_17001_),
    .Z(_17093_));
 AOI22_X2 _23179_ (.A1(\core.keymem.key_mem[12][88] ),
    .A2(_17093_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][88] ),
    .ZN(_17094_));
 NAND4_X2 _23180_ (.A1(_17089_),
    .A2(_17090_),
    .A3(_17092_),
    .A4(_17094_),
    .ZN(_17095_));
 OAI21_X4 _23181_ (.A(_17080_),
    .B1(_17088_),
    .B2(_17095_),
    .ZN(_17096_));
 XOR2_X2 _23182_ (.A(\core.dec_block.block_w1_reg[24] ),
    .B(_17096_),
    .Z(_17097_));
 AND2_X1 _23183_ (.A1(_00219_),
    .A2(_16496_),
    .ZN(_17098_));
 BUF_X4 _23184_ (.A(_16881_),
    .Z(_17099_));
 BUF_X4 _23185_ (.A(_17099_),
    .Z(_17100_));
 BUF_X4 _23186_ (.A(_17026_),
    .Z(_17101_));
 NAND3_X1 _23187_ (.A1(\core.keymem.key_mem[14][80] ),
    .A2(_17100_),
    .A3(_17101_),
    .ZN(_17102_));
 BUF_X4 _23188_ (.A(_17035_),
    .Z(_17103_));
 BUF_X4 _23189_ (.A(_17036_),
    .Z(_17104_));
 OAI211_X2 _23190_ (.A(\core.keymem.key_mem[10][80] ),
    .B(_17101_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_17105_));
 BUF_X4 _23191_ (.A(_17031_),
    .Z(_17106_));
 BUF_X4 _23192_ (.A(_17030_),
    .Z(_17107_));
 OAI211_X2 _23193_ (.A(\core.keymem.key_mem[6][80] ),
    .B(_17101_),
    .C1(_17106_),
    .C2(_17107_),
    .ZN(_17108_));
 NAND3_X1 _23194_ (.A1(\core.keymem.key_mem[12][80] ),
    .A2(_17100_),
    .A3(_17057_),
    .ZN(_17109_));
 NAND4_X2 _23195_ (.A1(_17102_),
    .A2(_17105_),
    .A3(_17108_),
    .A4(_17109_),
    .ZN(_17110_));
 BUF_X4 _23196_ (.A(_16938_),
    .Z(_17111_));
 BUF_X4 _23197_ (.A(_17111_),
    .Z(_17112_));
 OAI211_X2 _23198_ (.A(\core.keymem.key_mem[11][80] ),
    .B(_17112_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_17113_));
 BUF_X4 _23199_ (.A(_16908_),
    .Z(_17114_));
 BUF_X4 _23200_ (.A(_16917_),
    .Z(_17115_));
 BUF_X4 _23201_ (.A(_16913_),
    .Z(_17116_));
 BUF_X4 _23202_ (.A(_16914_),
    .Z(_17117_));
 BUF_X4 _23203_ (.A(_17117_),
    .Z(_17118_));
 OAI221_X2 _23204_ (.A(\core.keymem.key_mem[5][80] ),
    .B1(_17114_),
    .B2(_17115_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_17119_));
 BUF_X4 _23205_ (.A(_16969_),
    .Z(_17120_));
 BUF_X8 _23206_ (.A(_17120_),
    .Z(_17121_));
 OAI211_X2 _23207_ (.A(\core.keymem.key_mem[1][80] ),
    .B(_17121_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_17122_));
 OAI211_X2 _23208_ (.A(\core.keymem.key_mem[13][80] ),
    .B(_17100_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_17123_));
 NAND4_X2 _23209_ (.A1(_17113_),
    .A2(_17119_),
    .A3(_17122_),
    .A4(_17123_),
    .ZN(_17124_));
 OAI211_X2 _23210_ (.A(\core.keymem.key_mem[7][80] ),
    .B(_17112_),
    .C1(_17107_),
    .C2(_17106_),
    .ZN(_17125_));
 NAND3_X1 _23211_ (.A1(\core.keymem.key_mem[2][80] ),
    .A2(_17121_),
    .A3(_17050_),
    .ZN(_17126_));
 NAND3_X1 _23212_ (.A1(\core.keymem.key_mem[3][80] ),
    .A2(_17112_),
    .A3(_16970_),
    .ZN(_17127_));
 BUF_X4 _23213_ (.A(_16922_),
    .Z(_17128_));
 BUF_X4 _23214_ (.A(_16923_),
    .Z(_17129_));
 OAI221_X2 _23215_ (.A(\core.keymem.key_mem[9][80] ),
    .B1(_17128_),
    .B2(_17129_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_17130_));
 NAND4_X2 _23216_ (.A1(_17125_),
    .A2(_17126_),
    .A3(_17127_),
    .A4(_17130_),
    .ZN(_17131_));
 INV_X1 _23217_ (.A(\core.keymem.key_mem[4][80] ),
    .ZN(_17132_));
 OAI21_X1 _23218_ (.A(_17057_),
    .B1(_17107_),
    .B2(_17115_),
    .ZN(_17133_));
 OAI21_X4 _23219_ (.A(_16484_),
    .B1(_16884_),
    .B2(_16888_),
    .ZN(_17134_));
 INV_X1 _23220_ (.A(\core.keymem.key_mem[8][80] ),
    .ZN(_17135_));
 OAI22_X2 _23221_ (.A1(_17132_),
    .A2(_17133_),
    .B1(_17134_),
    .B2(_17135_),
    .ZN(_17136_));
 NOR4_X4 _23222_ (.A1(_17110_),
    .A2(_17124_),
    .A3(_17131_),
    .A4(_17136_),
    .ZN(_17137_));
 AOI21_X4 _23223_ (.A(_17098_),
    .B1(_17137_),
    .B2(_16489_),
    .ZN(_17138_));
 XNOR2_X2 _23224_ (.A(\core.dec_block.block_w1_reg[16] ),
    .B(_17138_),
    .ZN(_17139_));
 XNOR2_X1 _23225_ (.A(_17097_),
    .B(_17139_),
    .ZN(_17140_));
 XNOR2_X2 _23226_ (.A(_17079_),
    .B(_17140_),
    .ZN(_17141_));
 NAND2_X1 _23227_ (.A1(_00228_),
    .A2(_16983_),
    .ZN(_17142_));
 BUF_X4 _23228_ (.A(_17018_),
    .Z(_17143_));
 BUF_X4 _23229_ (.A(_17020_),
    .Z(_17144_));
 OAI211_X2 _23230_ (.A(\core.keymem.key_mem[1][95] ),
    .B(_17120_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_17145_));
 BUF_X4 _23231_ (.A(_16933_),
    .Z(_17146_));
 OAI211_X2 _23232_ (.A(\core.keymem.key_mem[4][95] ),
    .B(_17028_),
    .C1(_17146_),
    .C2(_17031_),
    .ZN(_17147_));
 NAND3_X1 _23233_ (.A1(\core.keymem.key_mem[3][95] ),
    .A2(_17111_),
    .A3(_17120_),
    .ZN(_17148_));
 BUF_X4 _23234_ (.A(_16912_),
    .Z(_17149_));
 OAI221_X1 _23235_ (.A(\core.keymem.key_mem[9][95] ),
    .B1(_16922_),
    .B2(_16923_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_17150_));
 AND4_X1 _23236_ (.A1(_17145_),
    .A2(_17147_),
    .A3(_17148_),
    .A4(_17150_),
    .ZN(_17151_));
 INV_X1 _23237_ (.A(\core.keymem.key_mem[12][95] ),
    .ZN(_17152_));
 INV_X1 _23238_ (.A(\core.keymem.key_mem[2][95] ),
    .ZN(_17153_));
 OAI33_X1 _23239_ (.A1(_17152_),
    .A2(_16390_),
    .A3(_16394_),
    .B1(_16383_),
    .B2(_16421_),
    .B3(_17153_),
    .ZN(_17154_));
 AOI221_X2 _23240_ (.A(_17154_),
    .B1(_16519_),
    .B2(\core.keymem.key_mem[6][95] ),
    .C1(\core.keymem.key_mem[11][95] ),
    .C2(_16441_),
    .ZN(_17155_));
 BUF_X4 _23241_ (.A(_17025_),
    .Z(_17156_));
 AND3_X1 _23242_ (.A1(\core.keymem.key_mem[10][95] ),
    .A2(_17156_),
    .A3(_17043_),
    .ZN(_17157_));
 NAND2_X1 _23243_ (.A1(\core.keymem.key_mem[13][95] ),
    .A2(_16961_),
    .ZN(_17158_));
 AOI21_X1 _23244_ (.A(_17158_),
    .B1(_16413_),
    .B2(_16411_),
    .ZN(_17159_));
 OAI21_X2 _23245_ (.A(_17055_),
    .B1(_17157_),
    .B2(_17159_),
    .ZN(_17160_));
 OAI221_X1 _23246_ (.A(\core.keymem.key_mem[5][95] ),
    .B1(_16908_),
    .B2(_16917_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_17161_));
 OAI211_X2 _23247_ (.A(\core.keymem.key_mem[7][95] ),
    .B(_17074_),
    .C1(_17030_),
    .C2(_16899_),
    .ZN(_17162_));
 BUF_X4 _23248_ (.A(_17025_),
    .Z(_17163_));
 NAND3_X1 _23249_ (.A1(\core.keymem.key_mem[14][95] ),
    .A2(_17099_),
    .A3(_17163_),
    .ZN(_17164_));
 OAI211_X2 _23250_ (.A(\core.keymem.key_mem[8][95] ),
    .B(_16893_),
    .C1(_17035_),
    .C2(_17036_),
    .ZN(_17165_));
 AND4_X1 _23251_ (.A1(_17161_),
    .A2(_17162_),
    .A3(_17164_),
    .A4(_17165_),
    .ZN(_17166_));
 NAND4_X4 _23252_ (.A1(_17151_),
    .A2(_17155_),
    .A3(_17160_),
    .A4(_17166_),
    .ZN(_17167_));
 OAI21_X4 _23253_ (.A(_17142_),
    .B1(_17167_),
    .B2(_16496_),
    .ZN(_17168_));
 XOR2_X2 _23254_ (.A(\core.dec_block.block_w1_reg[31] ),
    .B(_17168_),
    .Z(_17169_));
 INV_X1 _23255_ (.A(\core.dec_block.block_w1_reg[7] ),
    .ZN(_17170_));
 NAND2_X1 _23256_ (.A1(_00224_),
    .A2(_16497_),
    .ZN(_17171_));
 AOI22_X1 _23257_ (.A1(\core.keymem.key_mem[10][71] ),
    .A2(_16515_),
    .B1(_16398_),
    .B2(\core.keymem.key_mem[12][71] ),
    .ZN(_17172_));
 AOI22_X1 _23258_ (.A1(\core.keymem.key_mem[2][71] ),
    .A2(_16424_),
    .B1(_16462_),
    .B2(\core.keymem.key_mem[9][71] ),
    .ZN(_17173_));
 AOI22_X1 _23259_ (.A1(\core.keymem.key_mem[6][71] ),
    .A2(_16448_),
    .B1(_16949_),
    .B2(\core.keymem.key_mem[5][71] ),
    .ZN(_17174_));
 BUF_X8 _23260_ (.A(_16864_),
    .Z(_17175_));
 AOI22_X1 _23261_ (.A1(\core.keymem.key_mem[4][71] ),
    .A2(_16947_),
    .B1(_17175_),
    .B2(\core.keymem.key_mem[3][71] ),
    .ZN(_17176_));
 AND4_X1 _23262_ (.A1(_17172_),
    .A2(_17173_),
    .A3(_17174_),
    .A4(_17176_),
    .ZN(_17177_));
 BUF_X4 _23263_ (.A(_16855_),
    .Z(_17178_));
 AOI22_X2 _23264_ (.A1(\core.keymem.key_mem[11][71] ),
    .A2(_16507_),
    .B1(_17178_),
    .B2(\core.keymem.key_mem[1][71] ),
    .ZN(_17179_));
 AOI22_X4 _23265_ (.A1(\core.keymem.key_mem[7][71] ),
    .A2(_16513_),
    .B1(_16453_),
    .B2(\core.keymem.key_mem[8][71] ),
    .ZN(_17180_));
 AOI22_X2 _23266_ (.A1(\core.keymem.key_mem[14][71] ),
    .A2(_16502_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][71] ),
    .ZN(_17181_));
 NAND4_X4 _23267_ (.A1(_17177_),
    .A2(_17179_),
    .A3(_17180_),
    .A4(_17181_),
    .ZN(_17182_));
 BUF_X8 _23268_ (.A(_17014_),
    .Z(_17183_));
 OAI21_X4 _23269_ (.A(_17171_),
    .B1(_17182_),
    .B2(_17183_),
    .ZN(_17184_));
 XNOR2_X2 _23270_ (.A(_17170_),
    .B(_17184_),
    .ZN(_17185_));
 AOI21_X1 _23271_ (.A(_16494_),
    .B1(_17004_),
    .B2(\core.keymem.key_mem[5][69] ),
    .ZN(_17186_));
 AOI22_X1 _23272_ (.A1(\core.keymem.key_mem[4][69] ),
    .A2(_16456_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][69] ),
    .ZN(_17187_));
 AOI22_X1 _23273_ (.A1(\core.keymem.key_mem[7][69] ),
    .A2(_16955_),
    .B1(_16423_),
    .B2(\core.keymem.key_mem[2][69] ),
    .ZN(_17188_));
 AOI22_X1 _23274_ (.A1(\core.keymem.key_mem[8][69] ),
    .A2(_16528_),
    .B1(_16505_),
    .B2(\core.keymem.key_mem[11][69] ),
    .ZN(_17189_));
 AND4_X2 _23275_ (.A1(_17186_),
    .A2(_17187_),
    .A3(_17188_),
    .A4(_17189_),
    .ZN(_17190_));
 BUF_X8 _23276_ (.A(_16436_),
    .Z(_17191_));
 AOI222_X2 _23277_ (.A1(\core.keymem.key_mem[14][69] ),
    .A2(_17191_),
    .B1(_16447_),
    .B2(\core.keymem.key_mem[6][69] ),
    .C1(_16385_),
    .C2(\core.keymem.key_mem[3][69] ),
    .ZN(_17192_));
 BUF_X4 _23278_ (.A(_16471_),
    .Z(_17193_));
 AOI22_X1 _23279_ (.A1(\core.keymem.key_mem[10][69] ),
    .A2(_16988_),
    .B1(_17193_),
    .B2(\core.keymem.key_mem[13][69] ),
    .ZN(_17194_));
 AOI22_X1 _23280_ (.A1(\core.keymem.key_mem[9][69] ),
    .A2(_16535_),
    .B1(_16524_),
    .B2(\core.keymem.key_mem[1][69] ),
    .ZN(_17195_));
 AND3_X2 _23281_ (.A1(_17192_),
    .A2(_17194_),
    .A3(_17195_),
    .ZN(_17196_));
 AOI22_X4 _23282_ (.A1(_00223_),
    .A2(_17014_),
    .B1(_17190_),
    .B2(_17196_),
    .ZN(_17197_));
 XNOR2_X2 _23283_ (.A(\core.dec_block.block_w1_reg[5] ),
    .B(_17197_),
    .ZN(_17198_));
 XNOR2_X2 _23284_ (.A(_17185_),
    .B(_17198_),
    .ZN(_17199_));
 XNOR2_X1 _23285_ (.A(_17169_),
    .B(_17199_),
    .ZN(_17200_));
 XNOR2_X1 _23286_ (.A(_17141_),
    .B(_17200_),
    .ZN(_17201_));
 XNOR2_X1 _23287_ (.A(_17064_),
    .B(_17201_),
    .ZN(_17202_));
 AOI21_X4 _23288_ (.A(_16276_),
    .B1(_16368_),
    .B2(_16261_),
    .ZN(_17203_));
 BUF_X4 _23289_ (.A(_17203_),
    .Z(_17204_));
 OAI21_X1 _23290_ (.A(_16851_),
    .B1(_17202_),
    .B2(_17204_),
    .ZN(_17205_));
 OAI22_X1 _23291_ (.A1(\core.dec_block.block_w0_reg[0] ),
    .A2(_16366_),
    .B1(_16557_),
    .B2(_17205_),
    .ZN(_17206_));
 INV_X1 _23292_ (.A(_17206_),
    .ZN(_00567_));
 NAND2_X1 _23293_ (.A1(\core.dec_block.block_w0_reg[8] ),
    .A2(_16356_),
    .ZN(_17207_));
 AOI222_X2 _23294_ (.A1(\core.dec_block.block_w2_reg[8] ),
    .A2(_16565_),
    .B1(_16568_),
    .B2(\core.dec_block.block_w1_reg[8] ),
    .C1(_16266_),
    .C2(\core.dec_block.block_w3_reg[8] ),
    .ZN(_17208_));
 OAI21_X4 _23295_ (.A(_17207_),
    .B1(_17208_),
    .B2(_16357_),
    .ZN(_17209_));
 NAND2_X2 _23296_ (.A1(_16576_),
    .A2(_17209_),
    .ZN(_17210_));
 BUF_X4 _23297_ (.A(_17210_),
    .Z(_17211_));
 BUF_X4 _23298_ (.A(_17211_),
    .Z(_17212_));
 CLKBUF_X3 _23299_ (.A(_17212_),
    .Z(_17213_));
 BUF_X4 _23300_ (.A(_17213_),
    .Z(_17214_));
 NAND2_X1 _23301_ (.A1(_16355_),
    .A2(\core.dec_block.block_w0_reg[11] ),
    .ZN(_17215_));
 CLKBUF_X3 _23302_ (.A(\core.dec_block.block_w3_reg[11] ),
    .Z(_17216_));
 AOI222_X2 _23303_ (.A1(\core.dec_block.block_w2_reg[11] ),
    .A2(_16564_),
    .B1(_16567_),
    .B2(\core.dec_block.block_w1_reg[11] ),
    .C1(_16265_),
    .C2(_17216_),
    .ZN(_17217_));
 OAI21_X2 _23304_ (.A(_17215_),
    .B1(_17217_),
    .B2(_16356_),
    .ZN(_17218_));
 NAND2_X4 _23305_ (.A1(_16560_),
    .A2(_17218_),
    .ZN(_17219_));
 BUF_X4 _23306_ (.A(_17219_),
    .Z(_17220_));
 BUF_X4 _23307_ (.A(_17220_),
    .Z(_17221_));
 NAND2_X1 _23308_ (.A1(_16355_),
    .A2(\core.dec_block.block_w0_reg[10] ),
    .ZN(_17222_));
 AOI222_X2 _23309_ (.A1(\core.dec_block.block_w2_reg[10] ),
    .A2(_16564_),
    .B1(_16567_),
    .B2(\core.dec_block.block_w1_reg[10] ),
    .C1(_16265_),
    .C2(\core.dec_block.block_w3_reg[10] ),
    .ZN(_17223_));
 OAI21_X2 _23310_ (.A(_17222_),
    .B1(_17223_),
    .B2(_16355_),
    .ZN(_17224_));
 AND2_X1 _23311_ (.A1(_16559_),
    .A2(_17224_),
    .ZN(_17225_));
 BUF_X4 _23312_ (.A(_17225_),
    .Z(_17226_));
 BUF_X4 _23313_ (.A(_17226_),
    .Z(_17227_));
 BUF_X4 _23314_ (.A(_17227_),
    .Z(_17228_));
 BUF_X4 _23315_ (.A(_17228_),
    .Z(_17229_));
 NAND2_X1 _23316_ (.A1(_22132_),
    .A2(\core.dec_block.block_w0_reg[12] ),
    .ZN(_17230_));
 AOI222_X2 _23317_ (.A1(\core.dec_block.block_w2_reg[12] ),
    .A2(_16564_),
    .B1(_16567_),
    .B2(\core.dec_block.block_w1_reg[12] ),
    .C1(_16265_),
    .C2(\core.dec_block.block_w3_reg[12] ),
    .ZN(_17231_));
 OAI21_X2 _23318_ (.A(_17230_),
    .B1(_17231_),
    .B2(_16355_),
    .ZN(_17232_));
 AND2_X1 _23319_ (.A1(_16558_),
    .A2(_17232_),
    .ZN(_17233_));
 BUF_X4 _23320_ (.A(_17233_),
    .Z(_17234_));
 NAND2_X1 _23321_ (.A1(\core.dec_block.block_w0_reg[13] ),
    .A2(_16355_),
    .ZN(_17235_));
 AOI222_X2 _23322_ (.A1(\core.dec_block.block_w1_reg[13] ),
    .A2(_16567_),
    .B1(_16265_),
    .B2(\core.dec_block.block_w3_reg[13] ),
    .C1(\core.dec_block.block_w2_reg[13] ),
    .C2(_16564_),
    .ZN(_17236_));
 OAI21_X2 _23323_ (.A(_17235_),
    .B1(_17236_),
    .B2(_16355_),
    .ZN(_17237_));
 AND2_X4 _23324_ (.A1(_16559_),
    .A2(_17237_),
    .ZN(_17238_));
 BUF_X4 _23325_ (.A(_17238_),
    .Z(_17239_));
 NAND2_X1 _23326_ (.A1(_17234_),
    .A2(_17239_),
    .ZN(_17240_));
 NAND2_X1 _23327_ (.A1(_16355_),
    .A2(\core.dec_block.block_w0_reg[15] ),
    .ZN(_17241_));
 AOI222_X2 _23328_ (.A1(\core.dec_block.block_w1_reg[15] ),
    .A2(_16567_),
    .B1(_16265_),
    .B2(\core.dec_block.block_w3_reg[15] ),
    .C1(\core.dec_block.block_w2_reg[15] ),
    .C2(_16564_),
    .ZN(_17242_));
 OAI21_X2 _23329_ (.A(_17241_),
    .B1(_17242_),
    .B2(_16355_),
    .ZN(_17243_));
 AND2_X1 _23330_ (.A1(_16558_),
    .A2(_17243_),
    .ZN(_17244_));
 BUF_X4 _23331_ (.A(_17244_),
    .Z(_17245_));
 CLKBUF_X3 _23332_ (.A(\core.dec_block.block_w0_reg[14] ),
    .Z(_17246_));
 NAND2_X1 _23333_ (.A1(_22132_),
    .A2(_17246_),
    .ZN(_17247_));
 CLKBUF_X3 _23334_ (.A(\core.dec_block.block_w3_reg[14] ),
    .Z(_17248_));
 AOI222_X2 _23335_ (.A1(\core.dec_block.block_w1_reg[14] ),
    .A2(_16567_),
    .B1(_16265_),
    .B2(_17248_),
    .C1(\core.dec_block.block_w2_reg[14] ),
    .C2(_16564_),
    .ZN(_17249_));
 OAI21_X2 _23336_ (.A(_17247_),
    .B1(_17249_),
    .B2(_16355_),
    .ZN(_17250_));
 AND2_X1 _23337_ (.A1(_16558_),
    .A2(_17250_),
    .ZN(_17251_));
 BUF_X4 _23338_ (.A(_17251_),
    .Z(_17252_));
 NAND2_X4 _23339_ (.A1(_17245_),
    .A2(_17252_),
    .ZN(_17253_));
 NOR2_X2 _23340_ (.A1(_17240_),
    .A2(_17253_),
    .ZN(_17254_));
 BUF_X4 _23341_ (.A(_17254_),
    .Z(_17255_));
 NAND2_X1 _23342_ (.A1(_17229_),
    .A2(_17255_),
    .ZN(_17256_));
 NOR2_X1 _23343_ (.A1(_17221_),
    .A2(_17256_),
    .ZN(_17257_));
 CLKBUF_X3 _23344_ (.A(_17234_),
    .Z(_17258_));
 NOR2_X4 _23345_ (.A1(_17245_),
    .A2(_17252_),
    .ZN(_17259_));
 NAND2_X1 _23346_ (.A1(_16357_),
    .A2(\core.dec_block.block_w0_reg[9] ),
    .ZN(_17260_));
 AOI222_X2 _23347_ (.A1(\core.dec_block.block_w2_reg[9] ),
    .A2(_16565_),
    .B1(_16569_),
    .B2(\core.dec_block.block_w1_reg[9] ),
    .C1(_16266_),
    .C2(\core.dec_block.block_w3_reg[9] ),
    .ZN(_17261_));
 OAI21_X4 _23348_ (.A(_17260_),
    .B1(_17261_),
    .B2(_16584_),
    .ZN(_17262_));
 NAND2_X2 _23349_ (.A1(_16560_),
    .A2(_17262_),
    .ZN(_17263_));
 BUF_X4 _23350_ (.A(_17263_),
    .Z(_17264_));
 BUF_X4 _23351_ (.A(_17264_),
    .Z(_17265_));
 BUF_X4 _23352_ (.A(_17265_),
    .Z(_17266_));
 BUF_X4 _23353_ (.A(_17266_),
    .Z(_17267_));
 BUF_X4 _23354_ (.A(_17267_),
    .Z(_17268_));
 NAND2_X4 _23355_ (.A1(_16559_),
    .A2(_17224_),
    .ZN(_17269_));
 BUF_X4 _23356_ (.A(_17269_),
    .Z(_17270_));
 CLKBUF_X3 _23357_ (.A(_17270_),
    .Z(_17271_));
 BUF_X4 _23358_ (.A(_17271_),
    .Z(_17272_));
 CLKBUF_X3 _23359_ (.A(_17272_),
    .Z(_17273_));
 OAI21_X1 _23360_ (.A(_17259_),
    .B1(_17268_),
    .B2(_17273_),
    .ZN(_17274_));
 NAND2_X4 _23361_ (.A1(_16559_),
    .A2(_17232_),
    .ZN(_17275_));
 BUF_X4 _23362_ (.A(_17275_),
    .Z(_17276_));
 AND2_X1 _23363_ (.A1(_16561_),
    .A2(_17262_),
    .ZN(_17277_));
 BUF_X4 _23364_ (.A(_17277_),
    .Z(_17278_));
 BUF_X4 _23365_ (.A(_17278_),
    .Z(_17279_));
 BUF_X4 _23366_ (.A(_17279_),
    .Z(_17280_));
 CLKBUF_X3 _23367_ (.A(_17252_),
    .Z(_17281_));
 XNOR2_X1 _23368_ (.A(_17228_),
    .B(_17281_),
    .ZN(_17282_));
 NOR3_X1 _23369_ (.A1(_17276_),
    .A2(_17280_),
    .A3(_17282_),
    .ZN(_17283_));
 NAND2_X4 _23370_ (.A1(_16559_),
    .A2(_17250_),
    .ZN(_17284_));
 NOR2_X2 _23371_ (.A1(_17234_),
    .A2(_17284_),
    .ZN(_17285_));
 AOI21_X1 _23372_ (.A(_17283_),
    .B1(_17285_),
    .B2(_17229_),
    .ZN(_17286_));
 NAND2_X4 _23373_ (.A1(_16559_),
    .A2(_17243_),
    .ZN(_17287_));
 BUF_X4 _23374_ (.A(_17287_),
    .Z(_17288_));
 OAI22_X1 _23375_ (.A1(_17258_),
    .A2(_17274_),
    .B1(_17286_),
    .B2(_17288_),
    .ZN(_17289_));
 AND3_X1 _23376_ (.A1(_17221_),
    .A2(_17239_),
    .A3(_17289_),
    .ZN(_17290_));
 OAI21_X1 _23377_ (.A(_17214_),
    .B1(_17257_),
    .B2(_17290_),
    .ZN(_17291_));
 AND2_X1 _23378_ (.A1(_16560_),
    .A2(_17209_),
    .ZN(_17292_));
 BUF_X4 _23379_ (.A(_17292_),
    .Z(_17293_));
 NOR2_X4 _23380_ (.A1(_17293_),
    .A2(_17264_),
    .ZN(_17294_));
 NAND2_X4 _23381_ (.A1(_16559_),
    .A2(_17237_),
    .ZN(_17295_));
 CLKBUF_X3 _23382_ (.A(_17295_),
    .Z(_17296_));
 NOR2_X4 _23383_ (.A1(_17287_),
    .A2(_17252_),
    .ZN(_17297_));
 NAND2_X2 _23384_ (.A1(_17275_),
    .A2(_17297_),
    .ZN(_17298_));
 NOR2_X1 _23385_ (.A1(_17296_),
    .A2(_17298_),
    .ZN(_17299_));
 BUF_X4 _23386_ (.A(_17299_),
    .Z(_17300_));
 NOR2_X4 _23387_ (.A1(_17219_),
    .A2(_17269_),
    .ZN(_17301_));
 BUF_X4 _23388_ (.A(_17301_),
    .Z(_17302_));
 NAND3_X1 _23389_ (.A1(_17294_),
    .A2(_17300_),
    .A3(_17302_),
    .ZN(_17303_));
 NOR2_X4 _23390_ (.A1(_17219_),
    .A2(_17226_),
    .ZN(_17304_));
 NAND2_X4 _23391_ (.A1(_17294_),
    .A2(_17304_),
    .ZN(_17305_));
 NOR2_X4 _23392_ (.A1(_17275_),
    .A2(_17239_),
    .ZN(_17306_));
 NAND2_X2 _23393_ (.A1(_17297_),
    .A2(_17306_),
    .ZN(_17307_));
 BUF_X4 _23394_ (.A(_17307_),
    .Z(_17308_));
 NOR2_X4 _23395_ (.A1(_17275_),
    .A2(_17295_),
    .ZN(_17309_));
 NAND2_X4 _23396_ (.A1(_17309_),
    .A2(_17297_),
    .ZN(_17310_));
 NOR2_X1 _23397_ (.A1(_17210_),
    .A2(_17278_),
    .ZN(_17311_));
 AND2_X2 _23398_ (.A1(_16559_),
    .A2(_17218_),
    .ZN(_17312_));
 NOR2_X4 _23399_ (.A1(_17312_),
    .A2(_17226_),
    .ZN(_17313_));
 NAND2_X2 _23400_ (.A1(_17311_),
    .A2(_17313_),
    .ZN(_17314_));
 OAI221_X2 _23401_ (.A(_17303_),
    .B1(_17305_),
    .B2(_17308_),
    .C1(_17310_),
    .C2(_17314_),
    .ZN(_17315_));
 BUF_X4 _23402_ (.A(_17212_),
    .Z(_17316_));
 NAND2_X4 _23403_ (.A1(_17309_),
    .A2(_17259_),
    .ZN(_17317_));
 NAND2_X2 _23404_ (.A1(_17212_),
    .A2(_17300_),
    .ZN(_17318_));
 BUF_X4 _23405_ (.A(_17280_),
    .Z(_17319_));
 OAI22_X2 _23406_ (.A1(_17316_),
    .A2(_17317_),
    .B1(_17318_),
    .B2(_17319_),
    .ZN(_17320_));
 BUF_X4 _23407_ (.A(_17313_),
    .Z(_17321_));
 NAND2_X4 _23408_ (.A1(_17288_),
    .A2(_17284_),
    .ZN(_17322_));
 BUF_X4 _23409_ (.A(_17293_),
    .Z(_17323_));
 NAND2_X4 _23410_ (.A1(_17323_),
    .A2(_17265_),
    .ZN(_17324_));
 BUF_X4 _23411_ (.A(_17311_),
    .Z(_17325_));
 NOR2_X4 _23412_ (.A1(_17294_),
    .A2(_17325_),
    .ZN(_17326_));
 XNOR2_X1 _23413_ (.A(_17245_),
    .B(_17326_),
    .ZN(_17327_));
 OAI22_X2 _23414_ (.A1(_17322_),
    .A2(_17324_),
    .B1(_17327_),
    .B2(_17284_),
    .ZN(_17328_));
 BUF_X8 _23415_ (.A(_16562_),
    .Z(_17329_));
 OR2_X1 _23416_ (.A1(\core.dec_block.block_w0_reg[11] ),
    .A2(_17222_),
    .ZN(_17330_));
 AOI22_X1 _23417_ (.A1(\core.dec_block.block_w2_reg[11] ),
    .A2(_16565_),
    .B1(_16265_),
    .B2(_17216_),
    .ZN(_17331_));
 INV_X1 _23418_ (.A(_16568_),
    .ZN(_17332_));
 INV_X1 _23419_ (.A(\core.dec_block.block_w1_reg[11] ),
    .ZN(_17333_));
 OAI21_X1 _23420_ (.A(_17331_),
    .B1(_17332_),
    .B2(_17333_),
    .ZN(_17334_));
 OR3_X2 _23421_ (.A1(_16356_),
    .A2(_17334_),
    .A3(_17223_),
    .ZN(_17335_));
 NAND2_X1 _23422_ (.A1(_17330_),
    .A2(_17335_),
    .ZN(_17336_));
 NAND2_X4 _23423_ (.A1(_17329_),
    .A2(_17336_),
    .ZN(_17337_));
 BUF_X4 _23424_ (.A(_17337_),
    .Z(_17338_));
 NAND2_X4 _23425_ (.A1(_17275_),
    .A2(_17295_),
    .ZN(_17339_));
 NOR2_X1 _23426_ (.A1(_17338_),
    .A2(_17339_),
    .ZN(_17340_));
 AOI221_X2 _23427_ (.A(_17315_),
    .B1(_17320_),
    .B2(_17321_),
    .C1(_17328_),
    .C2(_17340_),
    .ZN(_17341_));
 NAND2_X4 _23428_ (.A1(_17219_),
    .A2(_17269_),
    .ZN(_17342_));
 NOR2_X4 _23429_ (.A1(_17264_),
    .A2(_17342_),
    .ZN(_17343_));
 NAND2_X2 _23430_ (.A1(_17287_),
    .A2(_17252_),
    .ZN(_17344_));
 NOR2_X1 _23431_ (.A1(_17240_),
    .A2(_17344_),
    .ZN(_17345_));
 BUF_X4 _23432_ (.A(_17345_),
    .Z(_17346_));
 NOR2_X4 _23433_ (.A1(_17245_),
    .A2(_17284_),
    .ZN(_17347_));
 NOR2_X4 _23434_ (.A1(_17234_),
    .A2(_17295_),
    .ZN(_17348_));
 AND2_X1 _23435_ (.A1(_17347_),
    .A2(_17348_),
    .ZN(_17349_));
 BUF_X4 _23436_ (.A(_17349_),
    .Z(_17350_));
 NOR2_X4 _23437_ (.A1(_17278_),
    .A2(_17337_),
    .ZN(_17351_));
 NAND2_X4 _23438_ (.A1(_17312_),
    .A2(_17226_),
    .ZN(_17352_));
 NAND2_X4 _23439_ (.A1(_17210_),
    .A2(_17264_),
    .ZN(_17353_));
 NOR2_X2 _23440_ (.A1(_17352_),
    .A2(_17353_),
    .ZN(_17354_));
 NOR4_X4 _23441_ (.A1(_17275_),
    .A2(_17238_),
    .A3(_17287_),
    .A4(_17252_),
    .ZN(_17355_));
 AOI222_X2 _23442_ (.A1(_17343_),
    .A2(_17346_),
    .B1(_17350_),
    .B2(_17351_),
    .C1(_17354_),
    .C2(_17355_),
    .ZN(_17356_));
 BUF_X4 _23443_ (.A(_17312_),
    .Z(_17357_));
 NAND2_X1 _23444_ (.A1(_17357_),
    .A2(_17279_),
    .ZN(_17358_));
 NOR2_X4 _23445_ (.A1(_17238_),
    .A2(_17298_),
    .ZN(_17359_));
 BUF_X4 _23446_ (.A(_17359_),
    .Z(_17360_));
 NOR2_X1 _23447_ (.A1(_17269_),
    .A2(_17288_),
    .ZN(_17361_));
 AOI22_X2 _23448_ (.A1(_17273_),
    .A2(_17360_),
    .B1(_17361_),
    .B2(_17306_),
    .ZN(_17362_));
 OAI21_X2 _23449_ (.A(_17356_),
    .B1(_17358_),
    .B2(_17362_),
    .ZN(_17363_));
 CLKBUF_X3 _23450_ (.A(_17319_),
    .Z(_17364_));
 NAND3_X4 _23451_ (.A1(_17238_),
    .A2(_17287_),
    .A3(_17284_),
    .ZN(_17365_));
 NOR2_X4 _23452_ (.A1(_17234_),
    .A2(_17365_),
    .ZN(_17366_));
 NAND2_X2 _23453_ (.A1(_17309_),
    .A2(_17347_),
    .ZN(_17367_));
 BUF_X4 _23454_ (.A(_17367_),
    .Z(_17368_));
 NOR2_X2 _23455_ (.A1(_17212_),
    .A2(_17368_),
    .ZN(_17369_));
 NOR3_X1 _23456_ (.A1(_17364_),
    .A2(_17366_),
    .A3(_17369_),
    .ZN(_17370_));
 BUF_X4 _23457_ (.A(_17323_),
    .Z(_17371_));
 BUF_X4 _23458_ (.A(_17371_),
    .Z(_17372_));
 NOR2_X1 _23459_ (.A1(_17372_),
    .A2(_17368_),
    .ZN(_17373_));
 CLKBUF_X3 _23460_ (.A(_17372_),
    .Z(_17374_));
 AOI21_X1 _23461_ (.A(_17373_),
    .B1(_17300_),
    .B2(_17374_),
    .ZN(_17375_));
 AOI21_X2 _23462_ (.A(_17370_),
    .B1(_17375_),
    .B2(_17364_),
    .ZN(_17376_));
 BUF_X4 _23463_ (.A(_17304_),
    .Z(_17377_));
 AOI21_X4 _23464_ (.A(_17363_),
    .B1(_17376_),
    .B2(_17377_),
    .ZN(_17378_));
 NAND3_X4 _23465_ (.A1(_16259_),
    .A2(_16351_),
    .A3(_16360_),
    .ZN(_17379_));
 AOI21_X4 _23466_ (.A(_17379_),
    .B1(_17330_),
    .B2(_17335_),
    .ZN(_17380_));
 BUF_X4 _23467_ (.A(_17380_),
    .Z(_17381_));
 NAND2_X4 _23468_ (.A1(_17234_),
    .A2(_17295_),
    .ZN(_17382_));
 NOR2_X1 _23469_ (.A1(_17322_),
    .A2(_17382_),
    .ZN(_17383_));
 BUF_X4 _23470_ (.A(_17383_),
    .Z(_17384_));
 NOR2_X4 _23471_ (.A1(_17288_),
    .A2(_17284_),
    .ZN(_17385_));
 NAND2_X2 _23472_ (.A1(_17385_),
    .A2(_17306_),
    .ZN(_17386_));
 NOR2_X2 _23473_ (.A1(_17212_),
    .A2(_17386_),
    .ZN(_17387_));
 MUX2_X1 _23474_ (.A(_17384_),
    .B(_17387_),
    .S(_17268_),
    .Z(_17388_));
 NOR3_X4 _23475_ (.A1(_17234_),
    .A2(_17287_),
    .A3(_17252_),
    .ZN(_17389_));
 NAND2_X1 _23476_ (.A1(_17296_),
    .A2(_17389_),
    .ZN(_17390_));
 BUF_X4 _23477_ (.A(_17390_),
    .Z(_17391_));
 NAND2_X1 _23478_ (.A1(_17210_),
    .A2(_17278_),
    .ZN(_17392_));
 BUF_X4 _23479_ (.A(_17392_),
    .Z(_17393_));
 OAI22_X1 _23480_ (.A1(_17214_),
    .A2(_17310_),
    .B1(_17391_),
    .B2(_17393_),
    .ZN(_17394_));
 AOI22_X2 _23481_ (.A1(_17381_),
    .A2(_17388_),
    .B1(_17394_),
    .B2(_17302_),
    .ZN(_17395_));
 OR2_X1 _23482_ (.A1(_17234_),
    .A2(_17365_),
    .ZN(_17396_));
 BUF_X4 _23483_ (.A(_17396_),
    .Z(_17397_));
 NOR2_X4 _23484_ (.A1(_17264_),
    .A2(_17337_),
    .ZN(_17398_));
 NAND2_X1 _23485_ (.A1(_17323_),
    .A2(_17398_),
    .ZN(_17399_));
 AOI21_X1 _23486_ (.A(_17397_),
    .B1(_17399_),
    .B2(_17305_),
    .ZN(_17400_));
 BUF_X4 _23487_ (.A(_17357_),
    .Z(_17401_));
 NOR2_X1 _23488_ (.A1(_17371_),
    .A2(_17401_),
    .ZN(_17402_));
 NOR2_X1 _23489_ (.A1(_17322_),
    .A2(_17339_),
    .ZN(_17403_));
 BUF_X4 _23490_ (.A(_17403_),
    .Z(_17404_));
 NOR2_X4 _23491_ (.A1(_17211_),
    .A2(_17219_),
    .ZN(_17405_));
 AOI22_X2 _23492_ (.A1(_17355_),
    .A2(_17402_),
    .B1(_17404_),
    .B2(_17405_),
    .ZN(_17406_));
 NOR3_X2 _23493_ (.A1(_17229_),
    .A2(_17268_),
    .A3(_17406_),
    .ZN(_17407_));
 NAND2_X1 _23494_ (.A1(_17360_),
    .A2(_17398_),
    .ZN(_17408_));
 NOR2_X1 _23495_ (.A1(_17372_),
    .A2(_17408_),
    .ZN(_17409_));
 NAND2_X1 _23496_ (.A1(_17304_),
    .A2(_17403_),
    .ZN(_17410_));
 NAND3_X1 _23497_ (.A1(_17220_),
    .A2(_17228_),
    .A3(_17300_),
    .ZN(_17411_));
 AOI21_X1 _23498_ (.A(_17353_),
    .B1(_17410_),
    .B2(_17411_),
    .ZN(_17412_));
 NOR4_X2 _23499_ (.A1(_17400_),
    .A2(_17407_),
    .A3(_17409_),
    .A4(_17412_),
    .ZN(_17413_));
 NOR2_X4 _23500_ (.A1(_17382_),
    .A2(_17344_),
    .ZN(_17414_));
 NAND2_X1 _23501_ (.A1(_17266_),
    .A2(_17414_),
    .ZN(_17415_));
 OAI21_X1 _23502_ (.A(_17415_),
    .B1(_17318_),
    .B2(_17268_),
    .ZN(_17416_));
 NAND2_X1 _23503_ (.A1(_17385_),
    .A2(_17348_),
    .ZN(_17417_));
 BUF_X4 _23504_ (.A(_17417_),
    .Z(_17418_));
 NOR2_X1 _23505_ (.A1(_17214_),
    .A2(_17418_),
    .ZN(_17419_));
 AOI22_X2 _23506_ (.A1(_17381_),
    .A2(_17416_),
    .B1(_17419_),
    .B2(_17343_),
    .ZN(_17420_));
 NOR2_X1 _23507_ (.A1(_17324_),
    .A2(_17352_),
    .ZN(_17421_));
 NOR3_X2 _23508_ (.A1(_17323_),
    .A2(_17265_),
    .A3(_17338_),
    .ZN(_17422_));
 NOR2_X1 _23509_ (.A1(_17421_),
    .A2(_17422_),
    .ZN(_17423_));
 NOR2_X1 _23510_ (.A1(_17308_),
    .A2(_17423_),
    .ZN(_17424_));
 NOR2_X1 _23511_ (.A1(_17326_),
    .A2(_17368_),
    .ZN(_17425_));
 NAND3_X1 _23512_ (.A1(_17220_),
    .A2(_17280_),
    .A3(_17387_),
    .ZN(_17426_));
 NAND2_X2 _23513_ (.A1(_17357_),
    .A2(_17266_),
    .ZN(_17427_));
 OR2_X1 _23514_ (.A1(_17339_),
    .A2(_17344_),
    .ZN(_17428_));
 BUF_X4 _23515_ (.A(_17428_),
    .Z(_17429_));
 OAI21_X1 _23516_ (.A(_17426_),
    .B1(_17427_),
    .B2(_17429_),
    .ZN(_17430_));
 AOI221_X2 _23517_ (.A(_17424_),
    .B1(_17425_),
    .B2(_17381_),
    .C1(_17430_),
    .C2(_17229_),
    .ZN(_17431_));
 NAND4_X1 _23518_ (.A1(_17395_),
    .A2(_17413_),
    .A3(_17420_),
    .A4(_17431_),
    .ZN(_17432_));
 NOR2_X4 _23519_ (.A1(_17293_),
    .A2(_17279_),
    .ZN(_17433_));
 NOR2_X4 _23520_ (.A1(_17211_),
    .A2(_17266_),
    .ZN(_17434_));
 AOI22_X2 _23521_ (.A1(_17401_),
    .A2(_17433_),
    .B1(_17434_),
    .B2(_17302_),
    .ZN(_17435_));
 NAND2_X4 _23522_ (.A1(_17264_),
    .A2(_17304_),
    .ZN(_17436_));
 NAND2_X4 _23523_ (.A1(_17239_),
    .A2(_17389_),
    .ZN(_17437_));
 OAI22_X2 _23524_ (.A1(_17317_),
    .A2(_17435_),
    .B1(_17436_),
    .B2(_17437_),
    .ZN(_17438_));
 NAND2_X4 _23525_ (.A1(_17279_),
    .A2(_17301_),
    .ZN(_17439_));
 NAND2_X2 _23526_ (.A1(_17263_),
    .A2(_17313_),
    .ZN(_17440_));
 NAND2_X4 _23527_ (.A1(_17306_),
    .A2(_17347_),
    .ZN(_17441_));
 OAI22_X2 _23528_ (.A1(_17429_),
    .A2(_17439_),
    .B1(_17440_),
    .B2(_17441_),
    .ZN(_17442_));
 NOR2_X1 _23529_ (.A1(_17338_),
    .A2(_17324_),
    .ZN(_17443_));
 AOI221_X2 _23530_ (.A(_17438_),
    .B1(_17442_),
    .B2(_17316_),
    .C1(_17384_),
    .C2(_17443_),
    .ZN(_17444_));
 NOR2_X4 _23531_ (.A1(_17278_),
    .A2(_17342_),
    .ZN(_17445_));
 NOR2_X2 _23532_ (.A1(_17253_),
    .A2(_17339_),
    .ZN(_17446_));
 AOI22_X2 _23533_ (.A1(_17357_),
    .A2(_17414_),
    .B1(_17445_),
    .B2(_17446_),
    .ZN(_17447_));
 NAND2_X4 _23534_ (.A1(_17259_),
    .A2(_17306_),
    .ZN(_17448_));
 OAI221_X2 _23535_ (.A(_17447_),
    .B1(_17436_),
    .B2(_17448_),
    .C1(_17314_),
    .C2(_17367_),
    .ZN(_17449_));
 NAND2_X4 _23536_ (.A1(_17293_),
    .A2(_17278_),
    .ZN(_17450_));
 NAND2_X2 _23537_ (.A1(_17347_),
    .A2(_17348_),
    .ZN(_17451_));
 OAI21_X1 _23538_ (.A(_17429_),
    .B1(_17450_),
    .B2(_17451_),
    .ZN(_17452_));
 OAI21_X1 _23539_ (.A(_17305_),
    .B1(_17342_),
    .B2(_17265_),
    .ZN(_17453_));
 AOI221_X2 _23540_ (.A(_17449_),
    .B1(_17452_),
    .B2(_17304_),
    .C1(_17453_),
    .C2(_17254_),
    .ZN(_17454_));
 NOR2_X2 _23541_ (.A1(_17339_),
    .A2(_17344_),
    .ZN(_17455_));
 BUF_X4 _23542_ (.A(_17455_),
    .Z(_17456_));
 MUX2_X1 _23543_ (.A(_17355_),
    .B(_17456_),
    .S(_17280_),
    .Z(_17457_));
 NAND2_X4 _23544_ (.A1(_17357_),
    .A2(_17269_),
    .ZN(_17458_));
 BUF_X4 _23545_ (.A(_17458_),
    .Z(_17459_));
 NOR2_X1 _23546_ (.A1(_17459_),
    .A2(_17450_),
    .ZN(_17460_));
 BUF_X4 _23547_ (.A(_17448_),
    .Z(_17461_));
 NAND3_X1 _23548_ (.A1(_17310_),
    .A2(_17461_),
    .A3(_17418_),
    .ZN(_17462_));
 NAND2_X4 _23549_ (.A1(_17309_),
    .A2(_17385_),
    .ZN(_17463_));
 BUF_X4 _23550_ (.A(_17266_),
    .Z(_17464_));
 OAI22_X1 _23551_ (.A1(_17463_),
    .A2(_17464_),
    .B1(_17461_),
    .B2(_17427_),
    .ZN(_17465_));
 AOI222_X2 _23552_ (.A1(_17321_),
    .A2(_17457_),
    .B1(_17460_),
    .B2(_17462_),
    .C1(_17465_),
    .C2(_17229_),
    .ZN(_17466_));
 BUF_X4 _23553_ (.A(_17451_),
    .Z(_17467_));
 BUF_X4 _23554_ (.A(_17386_),
    .Z(_17468_));
 AOI21_X1 _23555_ (.A(_17280_),
    .B1(_17467_),
    .B2(_17468_),
    .ZN(_17469_));
 OAI21_X1 _23556_ (.A(_17377_),
    .B1(_17387_),
    .B2(_17469_),
    .ZN(_17470_));
 NOR2_X4 _23557_ (.A1(_17276_),
    .A2(_17365_),
    .ZN(_17471_));
 NOR2_X4 _23558_ (.A1(_17279_),
    .A2(_17458_),
    .ZN(_17472_));
 AOI22_X1 _23559_ (.A1(_17471_),
    .A2(_17398_),
    .B1(_17472_),
    .B2(_17360_),
    .ZN(_17473_));
 OR2_X4 _23560_ (.A1(_17253_),
    .A2(_17339_),
    .ZN(_17474_));
 NAND2_X1 _23561_ (.A1(_17467_),
    .A2(_17474_),
    .ZN(_17475_));
 AOI21_X1 _23562_ (.A(_17475_),
    .B1(_17366_),
    .B2(_17372_),
    .ZN(_17476_));
 OAI221_X1 _23563_ (.A(_17470_),
    .B1(_17473_),
    .B2(_17372_),
    .C1(_17476_),
    .C2(_17439_),
    .ZN(_17477_));
 NOR2_X1 _23564_ (.A1(_17357_),
    .A2(_17463_),
    .ZN(_17478_));
 BUF_X4 _23565_ (.A(_17401_),
    .Z(_17479_));
 AOI21_X1 _23566_ (.A(_17478_),
    .B1(_17360_),
    .B2(_17479_),
    .ZN(_17480_));
 NOR3_X1 _23567_ (.A1(_17272_),
    .A2(_17324_),
    .A3(_17480_),
    .ZN(_17481_));
 BUF_X4 _23568_ (.A(_17401_),
    .Z(_17482_));
 NOR2_X2 _23569_ (.A1(_17293_),
    .A2(_17269_),
    .ZN(_17483_));
 NOR2_X1 _23570_ (.A1(_17211_),
    .A2(_17227_),
    .ZN(_17484_));
 OR2_X1 _23571_ (.A1(_17483_),
    .A2(_17484_),
    .ZN(_17485_));
 OR2_X2 _23572_ (.A1(_17322_),
    .A2(_17339_),
    .ZN(_17486_));
 NOR2_X2 _23573_ (.A1(_17267_),
    .A2(_17486_),
    .ZN(_17487_));
 NOR2_X1 _23574_ (.A1(_17271_),
    .A2(_17294_),
    .ZN(_17488_));
 AOI22_X1 _23575_ (.A1(_17485_),
    .A2(_17487_),
    .B1(_17488_),
    .B2(_17355_),
    .ZN(_17489_));
 NOR2_X1 _23576_ (.A1(_17482_),
    .A2(_17489_),
    .ZN(_17490_));
 BUF_X4 _23577_ (.A(_17446_),
    .Z(_17491_));
 NOR2_X4 _23578_ (.A1(_17293_),
    .A2(_17342_),
    .ZN(_17492_));
 AND2_X2 _23579_ (.A1(_17309_),
    .A2(_17297_),
    .ZN(_17493_));
 BUF_X4 _23580_ (.A(_17493_),
    .Z(_17494_));
 AOI22_X1 _23581_ (.A1(_17354_),
    .A2(_17491_),
    .B1(_17492_),
    .B2(_17494_),
    .ZN(_17495_));
 NOR2_X4 _23582_ (.A1(_17253_),
    .A2(_17382_),
    .ZN(_17496_));
 AOI22_X1 _23583_ (.A1(_17313_),
    .A2(_17496_),
    .B1(_17404_),
    .B2(_17302_),
    .ZN(_17497_));
 AOI22_X1 _23584_ (.A1(_17381_),
    .A2(_17360_),
    .B1(_17384_),
    .B2(_17492_),
    .ZN(_17498_));
 OAI221_X1 _23585_ (.A(_17495_),
    .B1(_17497_),
    .B2(_17393_),
    .C1(_17498_),
    .C2(_17319_),
    .ZN(_17499_));
 NOR4_X1 _23586_ (.A1(_17477_),
    .A2(_17481_),
    .A3(_17490_),
    .A4(_17499_),
    .ZN(_17500_));
 NAND4_X1 _23587_ (.A1(_17444_),
    .A2(_17454_),
    .A3(_17466_),
    .A4(_17500_),
    .ZN(_17501_));
 NOR2_X2 _23588_ (.A1(_17432_),
    .A2(_17501_),
    .ZN(_17502_));
 NAND4_X4 _23589_ (.A1(_17291_),
    .A2(_17341_),
    .A3(_17378_),
    .A4(_17502_),
    .ZN(_17503_));
 BUF_X4 _23590_ (.A(_17203_),
    .Z(_17504_));
 INV_X1 _23591_ (.A(\core.dec_block.block_w2_reg[7] ),
    .ZN(_17505_));
 BUF_X4 _23592_ (.A(_16451_),
    .Z(_17506_));
 AOI22_X1 _23593_ (.A1(\core.keymem.key_mem[8][39] ),
    .A2(_17506_),
    .B1(_16865_),
    .B2(\core.keymem.key_mem[3][39] ),
    .ZN(_17507_));
 AOI22_X1 _23594_ (.A1(\core.keymem.key_mem[2][39] ),
    .A2(_16859_),
    .B1(_16505_),
    .B2(\core.keymem.key_mem[11][39] ),
    .ZN(_17508_));
 AOI22_X1 _23595_ (.A1(\core.keymem.key_mem[10][39] ),
    .A2(_16514_),
    .B1(_16854_),
    .B2(\core.keymem.key_mem[1][39] ),
    .ZN(_17509_));
 AOI22_X1 _23596_ (.A1(\core.keymem.key_mem[4][39] ),
    .A2(_16456_),
    .B1(_16437_),
    .B2(\core.keymem.key_mem[14][39] ),
    .ZN(_17510_));
 NAND4_X1 _23597_ (.A1(_17507_),
    .A2(_17508_),
    .A3(_17509_),
    .A4(_17510_),
    .ZN(_17511_));
 AOI222_X2 _23598_ (.A1(\core.keymem.key_mem[7][39] ),
    .A2(_16406_),
    .B1(_16447_),
    .B2(\core.keymem.key_mem[6][39] ),
    .C1(_16397_),
    .C2(\core.keymem.key_mem[12][39] ),
    .ZN(_17512_));
 NAND2_X4 _23599_ (.A1(_16402_),
    .A2(_16404_),
    .ZN(_17513_));
 AOI222_X2 _23600_ (.A1(\core.keymem.key_mem[13][39] ),
    .A2(_17024_),
    .B1(_17513_),
    .B2(\core.keymem.key_mem[5][39] ),
    .C1(_17067_),
    .C2(\core.keymem.key_mem[9][39] ),
    .ZN(_17514_));
 OAI21_X1 _23601_ (.A(_17512_),
    .B1(_17514_),
    .B2(_16880_),
    .ZN(_17515_));
 NOR2_X1 _23602_ (.A1(_17511_),
    .A2(_17515_),
    .ZN(_17516_));
 MUX2_X2 _23603_ (.A(_00272_),
    .B(_17516_),
    .S(_16488_),
    .Z(_17517_));
 XNOR2_X2 _23604_ (.A(_17505_),
    .B(_17517_),
    .ZN(_17518_));
 INV_X1 _23605_ (.A(\core.dec_block.block_w2_reg[2] ),
    .ZN(_17519_));
 AOI22_X1 _23606_ (.A1(\core.keymem.key_mem[7][34] ),
    .A2(_16407_),
    .B1(_16986_),
    .B2(\core.keymem.key_mem[3][34] ),
    .ZN(_17520_));
 AOI22_X1 _23607_ (.A1(\core.keymem.key_mem[2][34] ),
    .A2(_16993_),
    .B1(_17004_),
    .B2(\core.keymem.key_mem[5][34] ),
    .ZN(_17521_));
 BUF_X4 _23608_ (.A(_16460_),
    .Z(_17522_));
 AOI22_X1 _23609_ (.A1(\core.keymem.key_mem[9][34] ),
    .A2(_17522_),
    .B1(_17000_),
    .B2(\core.keymem.key_mem[12][34] ),
    .ZN(_17523_));
 AOI22_X1 _23610_ (.A1(\core.keymem.key_mem[1][34] ),
    .A2(_16416_),
    .B1(_17193_),
    .B2(\core.keymem.key_mem[13][34] ),
    .ZN(_17524_));
 NAND4_X1 _23611_ (.A1(_17520_),
    .A2(_17521_),
    .A3(_17523_),
    .A4(_17524_),
    .ZN(_17525_));
 AOI22_X1 _23612_ (.A1(\core.keymem.key_mem[4][34] ),
    .A2(_16499_),
    .B1(_17007_),
    .B2(\core.keymem.key_mem[11][34] ),
    .ZN(_17526_));
 BUF_X4 _23613_ (.A(_16921_),
    .Z(_17527_));
 AOI22_X1 _23614_ (.A1(\core.keymem.key_mem[8][34] ),
    .A2(_17527_),
    .B1(_17156_),
    .B2(\core.keymem.key_mem[10][34] ),
    .ZN(_17528_));
 NOR2_X4 _23615_ (.A1(_16926_),
    .A2(_16928_),
    .ZN(_17529_));
 AOI22_X1 _23616_ (.A1(\core.keymem.key_mem[14][34] ),
    .A2(_16882_),
    .B1(_17513_),
    .B2(\core.keymem.key_mem[6][34] ),
    .ZN(_17530_));
 OAI221_X1 _23617_ (.A(_17526_),
    .B1(_17528_),
    .B2(_17529_),
    .C1(_16968_),
    .C2(_17530_),
    .ZN(_17531_));
 NOR2_X1 _23618_ (.A1(_17525_),
    .A2(_17531_),
    .ZN(_17532_));
 BUF_X8 _23619_ (.A(_16487_),
    .Z(_17533_));
 MUX2_X2 _23620_ (.A(_00279_),
    .B(_17532_),
    .S(_17533_),
    .Z(_17534_));
 XNOR2_X2 _23621_ (.A(_17519_),
    .B(_17534_),
    .ZN(_17535_));
 XNOR2_X2 _23622_ (.A(_17518_),
    .B(_17535_),
    .ZN(_17536_));
 BUF_X4 _23623_ (.A(\core.dec_block.block_w2_reg[23] ),
    .Z(_17537_));
 NAND3_X1 _23624_ (.A1(\core.keymem.key_mem[1][55] ),
    .A2(_16964_),
    .A3(_16967_),
    .ZN(_17538_));
 NAND3_X1 _23625_ (.A1(\core.keymem.key_mem[10][55] ),
    .A2(_17156_),
    .A3(_17054_),
    .ZN(_17539_));
 AOI21_X2 _23626_ (.A(_17051_),
    .B1(_17538_),
    .B2(_17539_),
    .ZN(_17540_));
 AOI22_X2 _23627_ (.A1(\core.keymem.key_mem[2][55] ),
    .A2(_16423_),
    .B1(_16441_),
    .B2(\core.keymem.key_mem[11][55] ),
    .ZN(_17541_));
 AOI22_X2 _23628_ (.A1(\core.keymem.key_mem[12][55] ),
    .A2(_17024_),
    .B1(_17513_),
    .B2(\core.keymem.key_mem[4][55] ),
    .ZN(_17542_));
 OAI21_X2 _23629_ (.A(_17541_),
    .B1(_17542_),
    .B2(_16394_),
    .ZN(_17543_));
 AOI22_X1 _23630_ (.A1(\core.keymem.key_mem[9][55] ),
    .A2(_16461_),
    .B1(_16471_),
    .B2(\core.keymem.key_mem[13][55] ),
    .ZN(_17544_));
 AOI22_X1 _23631_ (.A1(\core.keymem.key_mem[14][55] ),
    .A2(_16437_),
    .B1(_16948_),
    .B2(\core.keymem.key_mem[5][55] ),
    .ZN(_17545_));
 NAND2_X1 _23632_ (.A1(_17544_),
    .A2(_17545_),
    .ZN(_17546_));
 AOI22_X1 _23633_ (.A1(\core.keymem.key_mem[8][55] ),
    .A2(_16451_),
    .B1(_16864_),
    .B2(\core.keymem.key_mem[3][55] ),
    .ZN(_17547_));
 AOI22_X1 _23634_ (.A1(\core.keymem.key_mem[7][55] ),
    .A2(_16406_),
    .B1(_16447_),
    .B2(\core.keymem.key_mem[6][55] ),
    .ZN(_17548_));
 NAND2_X1 _23635_ (.A1(_17547_),
    .A2(_17548_),
    .ZN(_17549_));
 NOR4_X4 _23636_ (.A1(_17540_),
    .A2(_17543_),
    .A3(_17546_),
    .A4(_17549_),
    .ZN(_17550_));
 MUX2_X2 _23637_ (.A(_00259_),
    .B(_17550_),
    .S(_16487_),
    .Z(_17551_));
 XOR2_X2 _23638_ (.A(_17537_),
    .B(_17551_),
    .Z(_17552_));
 AOI222_X2 _23639_ (.A1(\core.keymem.key_mem[4][50] ),
    .A2(_16455_),
    .B1(_16422_),
    .B2(\core.keymem.key_mem[2][50] ),
    .C1(_16384_),
    .C2(\core.keymem.key_mem[3][50] ),
    .ZN(_17553_));
 AOI22_X1 _23640_ (.A1(\core.keymem.key_mem[14][50] ),
    .A2(_16436_),
    .B1(_16460_),
    .B2(\core.keymem.key_mem[9][50] ),
    .ZN(_17554_));
 AOI22_X1 _23641_ (.A1(\core.keymem.key_mem[11][50] ),
    .A2(_16504_),
    .B1(_16471_),
    .B2(\core.keymem.key_mem[13][50] ),
    .ZN(_17555_));
 AND3_X2 _23642_ (.A1(_17553_),
    .A2(_17554_),
    .A3(_17555_),
    .ZN(_17556_));
 AOI22_X1 _23643_ (.A1(\core.keymem.key_mem[6][50] ),
    .A2(_16519_),
    .B1(_16466_),
    .B2(\core.keymem.key_mem[5][50] ),
    .ZN(_17557_));
 AOI22_X1 _23644_ (.A1(\core.keymem.key_mem[8][50] ),
    .A2(_16450_),
    .B1(_16396_),
    .B2(\core.keymem.key_mem[12][50] ),
    .ZN(_17558_));
 AOI22_X1 _23645_ (.A1(\core.keymem.key_mem[7][50] ),
    .A2(_16954_),
    .B1(_16523_),
    .B2(\core.keymem.key_mem[1][50] ),
    .ZN(_17559_));
 AOI21_X1 _23646_ (.A(_16493_),
    .B1(_16431_),
    .B2(\core.keymem.key_mem[10][50] ),
    .ZN(_17560_));
 AND4_X2 _23647_ (.A1(_17557_),
    .A2(_17558_),
    .A3(_17559_),
    .A4(_17560_),
    .ZN(_17561_));
 AOI22_X4 _23648_ (.A1(_00280_),
    .A2(_17013_),
    .B1(_17556_),
    .B2(_17561_),
    .ZN(_17562_));
 XNOR2_X2 _23649_ (.A(\core.dec_block.block_w2_reg[18] ),
    .B(_17562_),
    .ZN(_17563_));
 AOI22_X1 _23650_ (.A1(\core.keymem.key_mem[3][54] ),
    .A2(_16384_),
    .B1(_16396_),
    .B2(\core.keymem.key_mem[12][54] ),
    .ZN(_17564_));
 AOI21_X1 _23651_ (.A(_16493_),
    .B1(_16405_),
    .B2(\core.keymem.key_mem[7][54] ),
    .ZN(_17565_));
 AOI22_X1 _23652_ (.A1(\core.keymem.key_mem[14][54] ),
    .A2(_16435_),
    .B1(_16440_),
    .B2(\core.keymem.key_mem[11][54] ),
    .ZN(_17566_));
 AOI22_X1 _23653_ (.A1(\core.keymem.key_mem[4][54] ),
    .A2(_16455_),
    .B1(_16430_),
    .B2(\core.keymem.key_mem[10][54] ),
    .ZN(_17567_));
 AND4_X2 _23654_ (.A1(_17564_),
    .A2(_17565_),
    .A3(_17566_),
    .A4(_17567_),
    .ZN(_17568_));
 AOI222_X2 _23655_ (.A1(\core.keymem.key_mem[6][54] ),
    .A2(_16446_),
    .B1(_16422_),
    .B2(\core.keymem.key_mem[2][54] ),
    .C1(_16414_),
    .C2(\core.keymem.key_mem[1][54] ),
    .ZN(_17569_));
 AOI22_X1 _23656_ (.A1(\core.keymem.key_mem[8][54] ),
    .A2(_16450_),
    .B1(_16470_),
    .B2(\core.keymem.key_mem[13][54] ),
    .ZN(_17570_));
 AOI22_X1 _23657_ (.A1(\core.keymem.key_mem[9][54] ),
    .A2(_16460_),
    .B1(_16466_),
    .B2(\core.keymem.key_mem[5][54] ),
    .ZN(_17571_));
 AND3_X2 _23658_ (.A1(_17569_),
    .A2(_17570_),
    .A3(_17571_),
    .ZN(_17572_));
 AOI22_X4 _23659_ (.A1(_00258_),
    .A2(_16545_),
    .B1(_17568_),
    .B2(_17572_),
    .ZN(_17573_));
 XNOR2_X2 _23660_ (.A(\core.dec_block.block_w2_reg[22] ),
    .B(_17573_),
    .ZN(_17574_));
 XOR2_X1 _23661_ (.A(_17563_),
    .B(_17574_),
    .Z(_17575_));
 XNOR2_X1 _23662_ (.A(_17552_),
    .B(_17575_),
    .ZN(_17576_));
 XNOR2_X2 _23663_ (.A(_17536_),
    .B(_17576_),
    .ZN(_17577_));
 BUF_X8 _23664_ (.A(_17183_),
    .Z(_17578_));
 AOI22_X1 _23665_ (.A1(\core.keymem.key_mem[6][58] ),
    .A2(_16522_),
    .B1(_17091_),
    .B2(\core.keymem.key_mem[3][58] ),
    .ZN(_17579_));
 AOI22_X2 _23666_ (.A1(\core.keymem.key_mem[8][58] ),
    .A2(_16530_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][58] ),
    .ZN(_17580_));
 BUF_X8 _23667_ (.A(_16999_),
    .Z(_17581_));
 AOI22_X2 _23668_ (.A1(\core.keymem.key_mem[14][58] ),
    .A2(_17581_),
    .B1(_17093_),
    .B2(\core.keymem.key_mem[12][58] ),
    .ZN(_17582_));
 AOI22_X2 _23669_ (.A1(\core.keymem.key_mem[7][58] ),
    .A2(_17085_),
    .B1(_16507_),
    .B2(\core.keymem.key_mem[11][58] ),
    .ZN(_17583_));
 NAND4_X2 _23670_ (.A1(_17579_),
    .A2(_17580_),
    .A3(_17582_),
    .A4(_17583_),
    .ZN(_17584_));
 BUF_X8 _23671_ (.A(_16463_),
    .Z(_17585_));
 AOI22_X1 _23672_ (.A1(\core.keymem.key_mem[9][58] ),
    .A2(_17585_),
    .B1(_16516_),
    .B2(\core.keymem.key_mem[10][58] ),
    .ZN(_17586_));
 AOI22_X2 _23673_ (.A1(\core.keymem.key_mem[4][58] ),
    .A2(_16501_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][58] ),
    .ZN(_17587_));
 AOI22_X2 _23674_ (.A1(\core.keymem.key_mem[2][58] ),
    .A2(_17086_),
    .B1(_16510_),
    .B2(\core.keymem.key_mem[5][58] ),
    .ZN(_17588_));
 NAND3_X2 _23675_ (.A1(_17586_),
    .A2(_17587_),
    .A3(_17588_),
    .ZN(_17589_));
 NOR3_X4 _23676_ (.A1(_17578_),
    .A2(_17584_),
    .A3(_17589_),
    .ZN(_17590_));
 AOI21_X4 _23677_ (.A(_17590_),
    .B1(_16549_),
    .B2(_00277_),
    .ZN(_17591_));
 XNOR2_X2 _23678_ (.A(\core.dec_block.block_w2_reg[26] ),
    .B(_17591_),
    .ZN(_17592_));
 AOI222_X2 _23679_ (.A1(\core.keymem.key_mem[7][62] ),
    .A2(_16407_),
    .B1(_16993_),
    .B2(\core.keymem.key_mem[2][62] ),
    .C1(_17007_),
    .C2(\core.keymem.key_mem[11][62] ),
    .ZN(_17593_));
 AOI22_X1 _23680_ (.A1(\core.keymem.key_mem[12][62] ),
    .A2(_16539_),
    .B1(_16416_),
    .B2(\core.keymem.key_mem[1][62] ),
    .ZN(_17594_));
 AOI22_X1 _23681_ (.A1(\core.keymem.key_mem[3][62] ),
    .A2(_16386_),
    .B1(_16515_),
    .B2(\core.keymem.key_mem[10][62] ),
    .ZN(_17595_));
 NAND3_X1 _23682_ (.A1(_17593_),
    .A2(_17594_),
    .A3(_17595_),
    .ZN(_17596_));
 AOI22_X1 _23683_ (.A1(\core.keymem.key_mem[5][62] ),
    .A2(_16949_),
    .B1(_16472_),
    .B2(\core.keymem.key_mem[13][62] ),
    .ZN(_17597_));
 AOI22_X1 _23684_ (.A1(\core.keymem.key_mem[4][62] ),
    .A2(_16947_),
    .B1(_16452_),
    .B2(\core.keymem.key_mem[8][62] ),
    .ZN(_17598_));
 AOI22_X1 _23685_ (.A1(\core.keymem.key_mem[14][62] ),
    .A2(_16998_),
    .B1(_16462_),
    .B2(\core.keymem.key_mem[9][62] ),
    .ZN(_17599_));
 AOI21_X1 _23686_ (.A(_16545_),
    .B1(_16448_),
    .B2(\core.keymem.key_mem[6][62] ),
    .ZN(_17600_));
 NAND4_X1 _23687_ (.A1(_17597_),
    .A2(_17598_),
    .A3(_17599_),
    .A4(_17600_),
    .ZN(_17601_));
 NOR2_X2 _23688_ (.A1(_17596_),
    .A2(_17601_),
    .ZN(_17602_));
 AOI21_X4 _23689_ (.A(_17602_),
    .B1(_16984_),
    .B2(_00268_),
    .ZN(_17603_));
 XNOR2_X2 _23690_ (.A(\core.dec_block.block_w2_reg[30] ),
    .B(_17603_),
    .ZN(_17604_));
 XOR2_X1 _23691_ (.A(_17592_),
    .B(_17604_),
    .Z(_17605_));
 INV_X1 _23692_ (.A(\core.dec_block.block_w2_reg[8] ),
    .ZN(_17606_));
 NAND2_X1 _23693_ (.A1(_00262_),
    .A2(_17183_),
    .ZN(_17607_));
 AOI22_X1 _23694_ (.A1(\core.keymem.key_mem[9][40] ),
    .A2(_16536_),
    .B1(_16532_),
    .B2(\core.keymem.key_mem[13][40] ),
    .ZN(_17608_));
 AOI22_X1 _23695_ (.A1(\core.keymem.key_mem[4][40] ),
    .A2(_16457_),
    .B1(_16515_),
    .B2(\core.keymem.key_mem[10][40] ),
    .ZN(_17609_));
 AOI22_X1 _23696_ (.A1(\core.keymem.key_mem[14][40] ),
    .A2(_16438_),
    .B1(_16424_),
    .B2(\core.keymem.key_mem[2][40] ),
    .ZN(_17610_));
 AOI22_X1 _23697_ (.A1(\core.keymem.key_mem[3][40] ),
    .A2(_16386_),
    .B1(_16398_),
    .B2(\core.keymem.key_mem[12][40] ),
    .ZN(_17611_));
 AND4_X1 _23698_ (.A1(_17608_),
    .A2(_17609_),
    .A3(_17610_),
    .A4(_17611_),
    .ZN(_17612_));
 AOI22_X2 _23699_ (.A1(\core.keymem.key_mem[6][40] ),
    .A2(_16449_),
    .B1(_16443_),
    .B2(\core.keymem.key_mem[11][40] ),
    .ZN(_17613_));
 AOI22_X2 _23700_ (.A1(\core.keymem.key_mem[8][40] ),
    .A2(_16530_),
    .B1(_16469_),
    .B2(\core.keymem.key_mem[5][40] ),
    .ZN(_17614_));
 AOI22_X2 _23701_ (.A1(\core.keymem.key_mem[7][40] ),
    .A2(_16513_),
    .B1(_17178_),
    .B2(\core.keymem.key_mem[1][40] ),
    .ZN(_17615_));
 NAND4_X2 _23702_ (.A1(_17612_),
    .A2(_17613_),
    .A3(_17614_),
    .A4(_17615_),
    .ZN(_17616_));
 OAI21_X4 _23703_ (.A(_17607_),
    .B1(_17616_),
    .B2(_16873_),
    .ZN(_17617_));
 XNOR2_X2 _23704_ (.A(_17606_),
    .B(_17617_),
    .ZN(_17618_));
 AND2_X1 _23705_ (.A1(_00256_),
    .A2(_16871_),
    .ZN(_17619_));
 NAND3_X1 _23706_ (.A1(\core.keymem.key_mem[12][56] ),
    .A2(_17100_),
    .A3(_17057_),
    .ZN(_17620_));
 OAI221_X2 _23707_ (.A(\core.keymem.key_mem[9][56] ),
    .B1(_17128_),
    .B2(_17129_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_17621_));
 BUF_X4 _23708_ (.A(_16934_),
    .Z(_17622_));
 OAI221_X2 _23709_ (.A(\core.keymem.key_mem[5][56] ),
    .B1(_17114_),
    .B2(_17622_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_17623_));
 OAI211_X2 _23710_ (.A(\core.keymem.key_mem[6][56] ),
    .B(_17050_),
    .C1(_17115_),
    .C2(_17114_),
    .ZN(_17624_));
 NAND4_X2 _23711_ (.A1(_17620_),
    .A2(_17621_),
    .A3(_17623_),
    .A4(_17624_),
    .ZN(_17625_));
 OAI211_X2 _23712_ (.A(\core.keymem.key_mem[1][56] ),
    .B(_16970_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_17626_));
 OAI211_X2 _23713_ (.A(\core.keymem.key_mem[11][56] ),
    .B(_17048_),
    .C1(_17128_),
    .C2(_17129_),
    .ZN(_17627_));
 NAND3_X1 _23714_ (.A1(\core.keymem.key_mem[2][56] ),
    .A2(_16970_),
    .A3(_17016_),
    .ZN(_17628_));
 OAI211_X2 _23715_ (.A(\core.keymem.key_mem[8][56] ),
    .B(_17527_),
    .C1(_17128_),
    .C2(_17129_),
    .ZN(_17629_));
 NAND4_X2 _23716_ (.A1(_17626_),
    .A2(_17627_),
    .A3(_17628_),
    .A4(_17629_),
    .ZN(_17630_));
 OAI211_X2 _23717_ (.A(\core.keymem.key_mem[10][56] ),
    .B(_17016_),
    .C1(_17128_),
    .C2(_17129_),
    .ZN(_17631_));
 OAI211_X2 _23718_ (.A(\core.keymem.key_mem[4][56] ),
    .B(_17527_),
    .C1(_17114_),
    .C2(_17115_),
    .ZN(_17632_));
 OAI211_X2 _23719_ (.A(\core.keymem.key_mem[7][56] ),
    .B(_17111_),
    .C1(_17114_),
    .C2(_17622_),
    .ZN(_17633_));
 NAND3_X1 _23720_ (.A1(\core.keymem.key_mem[14][56] ),
    .A2(_16882_),
    .A3(_17156_),
    .ZN(_17634_));
 NAND4_X2 _23721_ (.A1(_17631_),
    .A2(_17632_),
    .A3(_17633_),
    .A4(_17634_),
    .ZN(_17635_));
 INV_X1 _23722_ (.A(\core.keymem.key_mem[3][56] ),
    .ZN(_17636_));
 NAND2_X4 _23723_ (.A1(_16481_),
    .A2(_16969_),
    .ZN(_17637_));
 OAI21_X4 _23724_ (.A(_16881_),
    .B1(_16912_),
    .B2(_16914_),
    .ZN(_17638_));
 INV_X1 _23725_ (.A(\core.keymem.key_mem[13][56] ),
    .ZN(_17639_));
 OAI22_X2 _23726_ (.A1(_17636_),
    .A2(_17637_),
    .B1(_17638_),
    .B2(_17639_),
    .ZN(_17640_));
 NOR4_X4 _23727_ (.A1(_17625_),
    .A2(_17630_),
    .A3(_17635_),
    .A4(_17640_),
    .ZN(_17641_));
 AOI21_X4 _23728_ (.A(_17619_),
    .B1(_17641_),
    .B2(_17533_),
    .ZN(_17642_));
 XNOR2_X2 _23729_ (.A(\core.dec_block.block_w2_reg[24] ),
    .B(_17642_),
    .ZN(_17643_));
 XNOR2_X1 _23730_ (.A(_17618_),
    .B(_17643_),
    .ZN(_17644_));
 XNOR2_X1 _23731_ (.A(_17605_),
    .B(_17644_),
    .ZN(_17645_));
 AOI22_X2 _23732_ (.A1(\core.keymem.key_mem[9][38] ),
    .A2(_17522_),
    .B1(_16524_),
    .B2(\core.keymem.key_mem[1][38] ),
    .ZN(_17646_));
 AOI22_X2 _23733_ (.A1(\core.keymem.key_mem[14][38] ),
    .A2(_17191_),
    .B1(_16505_),
    .B2(\core.keymem.key_mem[11][38] ),
    .ZN(_17647_));
 BUF_X8 _23734_ (.A(_16519_),
    .Z(_17648_));
 AOI22_X2 _23735_ (.A1(\core.keymem.key_mem[6][38] ),
    .A2(_17648_),
    .B1(_16423_),
    .B2(\core.keymem.key_mem[2][38] ),
    .ZN(_17649_));
 AOI22_X2 _23736_ (.A1(\core.keymem.key_mem[4][38] ),
    .A2(_16456_),
    .B1(_16955_),
    .B2(\core.keymem.key_mem[7][38] ),
    .ZN(_17650_));
 NAND4_X2 _23737_ (.A1(_17646_),
    .A2(_17647_),
    .A3(_17649_),
    .A4(_17650_),
    .ZN(_17651_));
 AOI22_X2 _23738_ (.A1(\core.keymem.key_mem[3][38] ),
    .A2(_16986_),
    .B1(_16988_),
    .B2(\core.keymem.key_mem[10][38] ),
    .ZN(_17652_));
 AOI22_X2 _23739_ (.A1(\core.keymem.key_mem[8][38] ),
    .A2(_17506_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][38] ),
    .ZN(_17653_));
 AOI22_X2 _23740_ (.A1(\core.keymem.key_mem[5][38] ),
    .A2(_17004_),
    .B1(_17193_),
    .B2(\core.keymem.key_mem[13][38] ),
    .ZN(_17654_));
 NAND3_X2 _23741_ (.A1(_17652_),
    .A2(_17653_),
    .A3(_17654_),
    .ZN(_17655_));
 NOR3_X4 _23742_ (.A1(_16546_),
    .A2(_17651_),
    .A3(_17655_),
    .ZN(_17656_));
 AOI21_X4 _23743_ (.A(_17656_),
    .B1(_16852_),
    .B2(_00264_),
    .ZN(_17657_));
 XNOR2_X2 _23744_ (.A(_16589_),
    .B(_17657_),
    .ZN(_17658_));
 NAND2_X1 _23745_ (.A1(_00273_),
    .A2(_16872_),
    .ZN(_17659_));
 AOI22_X4 _23746_ (.A1(\core.keymem.key_mem[12][33] ),
    .A2(_17001_),
    .B1(_16525_),
    .B2(\core.keymem.key_mem[1][33] ),
    .ZN(_17660_));
 AOI22_X1 _23747_ (.A1(\core.keymem.key_mem[2][33] ),
    .A2(_16859_),
    .B1(_16531_),
    .B2(\core.keymem.key_mem[13][33] ),
    .ZN(_17661_));
 AOI22_X1 _23748_ (.A1(\core.keymem.key_mem[14][33] ),
    .A2(_17191_),
    .B1(_16865_),
    .B2(\core.keymem.key_mem[3][33] ),
    .ZN(_17662_));
 AOI22_X1 _23749_ (.A1(\core.keymem.key_mem[4][33] ),
    .A2(_16456_),
    .B1(_16514_),
    .B2(\core.keymem.key_mem[10][33] ),
    .ZN(_17663_));
 AOI22_X1 _23750_ (.A1(\core.keymem.key_mem[7][33] ),
    .A2(_16955_),
    .B1(_16505_),
    .B2(\core.keymem.key_mem[11][33] ),
    .ZN(_17664_));
 AND4_X1 _23751_ (.A1(_17661_),
    .A2(_17662_),
    .A3(_17663_),
    .A4(_17664_),
    .ZN(_17665_));
 BUF_X8 _23752_ (.A(_17506_),
    .Z(_17666_));
 AOI22_X2 _23753_ (.A1(\core.keymem.key_mem[6][33] ),
    .A2(_16521_),
    .B1(_17666_),
    .B2(\core.keymem.key_mem[8][33] ),
    .ZN(_17667_));
 BUF_X4 _23754_ (.A(_16535_),
    .Z(_17668_));
 AOI22_X2 _23755_ (.A1(\core.keymem.key_mem[9][33] ),
    .A2(_17668_),
    .B1(_16509_),
    .B2(\core.keymem.key_mem[5][33] ),
    .ZN(_17669_));
 NAND4_X4 _23756_ (.A1(_17660_),
    .A2(_17665_),
    .A3(_17667_),
    .A4(_17669_),
    .ZN(_17670_));
 OAI21_X4 _23757_ (.A(_17659_),
    .B1(_17670_),
    .B2(_16547_),
    .ZN(_17671_));
 XOR2_X2 _23758_ (.A(\core.dec_block.block_w2_reg[1] ),
    .B(_17671_),
    .Z(_17672_));
 XNOR2_X2 _23759_ (.A(_17658_),
    .B(_17672_),
    .ZN(_17673_));
 AOI22_X1 _23760_ (.A1(\core.keymem.key_mem[9][41] ),
    .A2(_16537_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][41] ),
    .ZN(_17674_));
 BUF_X8 _23761_ (.A(_16949_),
    .Z(_17675_));
 AOI22_X2 _23762_ (.A1(\core.keymem.key_mem[14][41] ),
    .A2(_16502_),
    .B1(_17675_),
    .B2(\core.keymem.key_mem[5][41] ),
    .ZN(_17676_));
 AOI22_X2 _23763_ (.A1(\core.keymem.key_mem[4][41] ),
    .A2(_16458_),
    .B1(_16443_),
    .B2(\core.keymem.key_mem[11][41] ),
    .ZN(_17677_));
 AOI21_X1 _23764_ (.A(_16546_),
    .B1(_16453_),
    .B2(\core.keymem.key_mem[8][41] ),
    .ZN(_17678_));
 NAND4_X2 _23765_ (.A1(_17674_),
    .A2(_17676_),
    .A3(_17677_),
    .A4(_17678_),
    .ZN(_17679_));
 MUX2_X1 _23766_ (.A(\core.keymem.key_mem[2][41] ),
    .B(\core.keymem.key_mem[10][41] ),
    .S(_17055_),
    .Z(_17680_));
 AOI22_X1 _23767_ (.A1(\core.keymem.key_mem[6][41] ),
    .A2(_17513_),
    .B1(_17043_),
    .B2(_17680_),
    .ZN(_17681_));
 NOR2_X1 _23768_ (.A1(_16968_),
    .A2(_17681_),
    .ZN(_17682_));
 BUF_X4 _23769_ (.A(_17175_),
    .Z(_17683_));
 AOI22_X1 _23770_ (.A1(\core.keymem.key_mem[7][41] ),
    .A2(_16513_),
    .B1(_17683_),
    .B2(\core.keymem.key_mem[3][41] ),
    .ZN(_17684_));
 AOI22_X1 _23771_ (.A1(\core.keymem.key_mem[1][41] ),
    .A2(_17178_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][41] ),
    .ZN(_17685_));
 NAND2_X1 _23772_ (.A1(_17684_),
    .A2(_17685_),
    .ZN(_17686_));
 NOR3_X4 _23773_ (.A1(_17679_),
    .A2(_17682_),
    .A3(_17686_),
    .ZN(_17687_));
 AOI21_X4 _23774_ (.A(_17687_),
    .B1(_16498_),
    .B2(_00271_),
    .ZN(_17688_));
 XNOR2_X2 _23775_ (.A(\core.dec_block.block_w2_reg[9] ),
    .B(_17688_),
    .ZN(_17689_));
 AOI22_X2 _23776_ (.A1(\core.keymem.key_mem[4][46] ),
    .A2(_16457_),
    .B1(_16462_),
    .B2(\core.keymem.key_mem[9][46] ),
    .ZN(_17690_));
 AOI22_X2 _23777_ (.A1(\core.keymem.key_mem[7][46] ),
    .A2(_16512_),
    .B1(_16386_),
    .B2(\core.keymem.key_mem[3][46] ),
    .ZN(_17691_));
 AOI22_X2 _23778_ (.A1(\core.keymem.key_mem[14][46] ),
    .A2(_16438_),
    .B1(_16452_),
    .B2(\core.keymem.key_mem[8][46] ),
    .ZN(_17692_));
 AOI22_X2 _23779_ (.A1(\core.keymem.key_mem[2][46] ),
    .A2(_16424_),
    .B1(_16432_),
    .B2(\core.keymem.key_mem[10][46] ),
    .ZN(_17693_));
 NAND4_X2 _23780_ (.A1(_17690_),
    .A2(_17691_),
    .A3(_17692_),
    .A4(_17693_),
    .ZN(_17694_));
 BUF_X8 _23781_ (.A(_17648_),
    .Z(_17695_));
 AOI22_X2 _23782_ (.A1(\core.keymem.key_mem[6][46] ),
    .A2(_17695_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][46] ),
    .ZN(_17696_));
 AOI22_X2 _23783_ (.A1(\core.keymem.key_mem[11][46] ),
    .A2(_16506_),
    .B1(_16532_),
    .B2(\core.keymem.key_mem[13][46] ),
    .ZN(_17697_));
 AOI22_X2 _23784_ (.A1(\core.keymem.key_mem[12][46] ),
    .A2(_16539_),
    .B1(_16416_),
    .B2(\core.keymem.key_mem[1][46] ),
    .ZN(_17698_));
 NAND3_X2 _23785_ (.A1(_17696_),
    .A2(_17697_),
    .A3(_17698_),
    .ZN(_17699_));
 NOR3_X4 _23786_ (.A1(_16852_),
    .A2(_17694_),
    .A3(_17699_),
    .ZN(_17700_));
 AOI21_X4 _23787_ (.A(_17700_),
    .B1(_17183_),
    .B2(_00270_),
    .ZN(_17701_));
 XNOR2_X2 _23788_ (.A(\core.dec_block.block_w2_reg[14] ),
    .B(_17701_),
    .ZN(_17702_));
 XNOR2_X2 _23789_ (.A(_17689_),
    .B(_17702_),
    .ZN(_17703_));
 XNOR2_X1 _23790_ (.A(_17673_),
    .B(_17703_),
    .ZN(_17704_));
 XNOR2_X1 _23791_ (.A(_17645_),
    .B(_17704_),
    .ZN(_17705_));
 XNOR2_X1 _23792_ (.A(_17577_),
    .B(_17705_),
    .ZN(_17706_));
 NOR2_X1 _23793_ (.A1(_17504_),
    .A2(_17706_),
    .ZN(_17707_));
 NAND2_X1 _23794_ (.A1(_16260_),
    .A2(_16368_),
    .ZN(_17708_));
 BUF_X4 _23795_ (.A(_17708_),
    .Z(_17709_));
 BUF_X4 _23796_ (.A(_17709_),
    .Z(_17710_));
 INV_X1 _23797_ (.A(\block_reg[2][10] ),
    .ZN(_17711_));
 AOI22_X1 _23798_ (.A1(\core.keymem.key_mem[6][42] ),
    .A2(_16521_),
    .B1(_17666_),
    .B2(\core.keymem.key_mem[8][42] ),
    .ZN(_17712_));
 BUF_X8 _23799_ (.A(_16499_),
    .Z(_17713_));
 AOI22_X1 _23800_ (.A1(\core.keymem.key_mem[4][42] ),
    .A2(_17713_),
    .B1(_17084_),
    .B2(\core.keymem.key_mem[7][42] ),
    .ZN(_17714_));
 BUF_X8 _23801_ (.A(_16988_),
    .Z(_17715_));
 AOI22_X1 _23802_ (.A1(\core.keymem.key_mem[2][42] ),
    .A2(_16860_),
    .B1(_17715_),
    .B2(\core.keymem.key_mem[10][42] ),
    .ZN(_17716_));
 AOI22_X1 _23803_ (.A1(\core.keymem.key_mem[9][42] ),
    .A2(_17668_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][42] ),
    .ZN(_17717_));
 NAND4_X1 _23804_ (.A1(_17712_),
    .A2(_17714_),
    .A3(_17716_),
    .A4(_17717_),
    .ZN(_17718_));
 BUF_X8 _23805_ (.A(_17191_),
    .Z(_17719_));
 BUF_X4 _23806_ (.A(_17000_),
    .Z(_17720_));
 AOI22_X1 _23807_ (.A1(\core.keymem.key_mem[14][42] ),
    .A2(_17719_),
    .B1(_17720_),
    .B2(\core.keymem.key_mem[12][42] ),
    .ZN(_17721_));
 BUF_X4 _23808_ (.A(_17193_),
    .Z(_17722_));
 AOI22_X1 _23809_ (.A1(\core.keymem.key_mem[1][42] ),
    .A2(_16525_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][42] ),
    .ZN(_17723_));
 AOI22_X1 _23810_ (.A1(\core.keymem.key_mem[3][42] ),
    .A2(_16866_),
    .B1(_16506_),
    .B2(\core.keymem.key_mem[11][42] ),
    .ZN(_17724_));
 NAND3_X1 _23811_ (.A1(_17721_),
    .A2(_17723_),
    .A3(_17724_),
    .ZN(_17725_));
 NOR2_X2 _23812_ (.A1(_17718_),
    .A2(_17725_),
    .ZN(_17726_));
 MUX2_X2 _23813_ (.A(_00278_),
    .B(_17726_),
    .S(_17533_),
    .Z(_17727_));
 XNOR2_X1 _23814_ (.A(_17711_),
    .B(_17727_),
    .ZN(_17728_));
 AOI22_X1 _23815_ (.A1(\core.keymem.key_mem[4][106] ),
    .A2(_16456_),
    .B1(_16505_),
    .B2(\core.keymem.key_mem[11][106] ),
    .ZN(_17729_));
 AOI21_X1 _23816_ (.A(_16494_),
    .B1(_16986_),
    .B2(\core.keymem.key_mem[3][106] ),
    .ZN(_17730_));
 AOI22_X1 _23817_ (.A1(\core.keymem.key_mem[6][106] ),
    .A2(_17648_),
    .B1(_16423_),
    .B2(\core.keymem.key_mem[2][106] ),
    .ZN(_17731_));
 AOI22_X1 _23818_ (.A1(\core.keymem.key_mem[9][106] ),
    .A2(_16535_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][106] ),
    .ZN(_17732_));
 AND4_X1 _23819_ (.A1(_17729_),
    .A2(_17730_),
    .A3(_17731_),
    .A4(_17732_),
    .ZN(_17733_));
 AOI222_X2 _23820_ (.A1(\core.keymem.key_mem[14][106] ),
    .A2(_16437_),
    .B1(_16431_),
    .B2(\core.keymem.key_mem[10][106] ),
    .C1(_16471_),
    .C2(\core.keymem.key_mem[13][106] ),
    .ZN(_17734_));
 AOI22_X1 _23821_ (.A1(\core.keymem.key_mem[1][106] ),
    .A2(_16524_),
    .B1(_16467_),
    .B2(\core.keymem.key_mem[5][106] ),
    .ZN(_17735_));
 BUF_X8 _23822_ (.A(_16954_),
    .Z(_17736_));
 AOI22_X1 _23823_ (.A1(\core.keymem.key_mem[7][106] ),
    .A2(_17736_),
    .B1(_16528_),
    .B2(\core.keymem.key_mem[8][106] ),
    .ZN(_17737_));
 AND3_X1 _23824_ (.A1(_17734_),
    .A2(_17735_),
    .A3(_17737_),
    .ZN(_17738_));
 AOI22_X4 _23825_ (.A1(_00199_),
    .A2(_16496_),
    .B1(_17733_),
    .B2(_17738_),
    .ZN(_17739_));
 XNOR2_X2 _23826_ (.A(\core.dec_block.block_w0_reg[10] ),
    .B(_17739_),
    .ZN(_17740_));
 BUF_X4 _23827_ (.A(_16554_),
    .Z(_17741_));
 OAI221_X1 _23828_ (.A(_16364_),
    .B1(_17710_),
    .B2(_17728_),
    .C1(_17740_),
    .C2(_17741_),
    .ZN(_17742_));
 NOR3_X1 _23829_ (.A1(_17503_),
    .A2(_17707_),
    .A3(_17742_),
    .ZN(_17743_));
 CLKBUF_X3 _23830_ (.A(_16367_),
    .Z(_17744_));
 INV_X1 _23831_ (.A(\core.dec_block.block_w0_reg[10] ),
    .ZN(_17745_));
 AOI21_X1 _23832_ (.A(_17743_),
    .B1(_17744_),
    .B2(_17745_),
    .ZN(_00568_));
 INV_X1 _23833_ (.A(\core.dec_block.block_w0_reg[11] ),
    .ZN(_17746_));
 OAI22_X4 _23834_ (.A1(_16259_),
    .A2(_16275_),
    .B1(_16369_),
    .B2(_16260_),
    .ZN(_17747_));
 BUF_X4 _23835_ (.A(_17747_),
    .Z(_17748_));
 BUF_X4 _23836_ (.A(_17748_),
    .Z(_17749_));
 AOI22_X1 _23837_ (.A1(\core.keymem.key_mem[14][37] ),
    .A2(_16998_),
    .B1(_16520_),
    .B2(\core.keymem.key_mem[6][37] ),
    .ZN(_17750_));
 AOI22_X1 _23838_ (.A1(\core.keymem.key_mem[5][37] ),
    .A2(_17004_),
    .B1(_17193_),
    .B2(\core.keymem.key_mem[13][37] ),
    .ZN(_17751_));
 AOI22_X1 _23839_ (.A1(\core.keymem.key_mem[2][37] ),
    .A2(_16993_),
    .B1(_16986_),
    .B2(\core.keymem.key_mem[3][37] ),
    .ZN(_17752_));
 AOI22_X1 _23840_ (.A1(\core.keymem.key_mem[12][37] ),
    .A2(_17000_),
    .B1(_16524_),
    .B2(\core.keymem.key_mem[1][37] ),
    .ZN(_17753_));
 NAND4_X1 _23841_ (.A1(_17750_),
    .A2(_17751_),
    .A3(_17752_),
    .A4(_17753_),
    .ZN(_17754_));
 AOI22_X1 _23842_ (.A1(\core.keymem.key_mem[4][37] ),
    .A2(_16947_),
    .B1(_17506_),
    .B2(\core.keymem.key_mem[8][37] ),
    .ZN(_17755_));
 AOI22_X1 _23843_ (.A1(\core.keymem.key_mem[7][37] ),
    .A2(_17736_),
    .B1(_17522_),
    .B2(\core.keymem.key_mem[9][37] ),
    .ZN(_17756_));
 AOI22_X1 _23844_ (.A1(\core.keymem.key_mem[10][37] ),
    .A2(_16432_),
    .B1(_17007_),
    .B2(\core.keymem.key_mem[11][37] ),
    .ZN(_17757_));
 NAND3_X1 _23845_ (.A1(_17755_),
    .A2(_17756_),
    .A3(_17757_),
    .ZN(_17758_));
 NOR3_X2 _23846_ (.A1(_16983_),
    .A2(_17754_),
    .A3(_17758_),
    .ZN(_17759_));
 AOI21_X4 _23847_ (.A(_17759_),
    .B1(_16547_),
    .B2(_00263_),
    .ZN(_17760_));
 XNOR2_X2 _23848_ (.A(\core.dec_block.block_w2_reg[5] ),
    .B(_17760_),
    .ZN(_17761_));
 XNOR2_X2 _23849_ (.A(_17518_),
    .B(_17761_),
    .ZN(_17762_));
 AOI222_X2 _23850_ (.A1(\core.keymem.key_mem[7][32] ),
    .A2(_17085_),
    .B1(_16522_),
    .B2(\core.keymem.key_mem[6][32] ),
    .C1(_17091_),
    .C2(\core.keymem.key_mem[3][32] ),
    .ZN(_17763_));
 AOI22_X2 _23851_ (.A1(\core.keymem.key_mem[10][32] ),
    .A2(_17082_),
    .B1(_17093_),
    .B2(\core.keymem.key_mem[12][32] ),
    .ZN(_17764_));
 BUF_X8 _23852_ (.A(_16453_),
    .Z(_17765_));
 AOI22_X2 _23853_ (.A1(\core.keymem.key_mem[8][32] ),
    .A2(_17765_),
    .B1(_17585_),
    .B2(\core.keymem.key_mem[9][32] ),
    .ZN(_17766_));
 NAND3_X2 _23854_ (.A1(_17763_),
    .A2(_17764_),
    .A3(_17766_),
    .ZN(_17767_));
 BUF_X8 _23855_ (.A(_16442_),
    .Z(_17768_));
 BUF_X8 _23856_ (.A(_17768_),
    .Z(_17769_));
 AOI22_X1 _23857_ (.A1(\core.keymem.key_mem[2][32] ),
    .A2(_17086_),
    .B1(_17769_),
    .B2(\core.keymem.key_mem[11][32] ),
    .ZN(_17770_));
 BUF_X8 _23858_ (.A(_16473_),
    .Z(_17771_));
 AOI22_X2 _23859_ (.A1(\core.keymem.key_mem[1][32] ),
    .A2(_16526_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][32] ),
    .ZN(_17772_));
 AOI22_X2 _23860_ (.A1(\core.keymem.key_mem[4][32] ),
    .A2(_16501_),
    .B1(_16510_),
    .B2(\core.keymem.key_mem[5][32] ),
    .ZN(_17773_));
 AOI21_X1 _23861_ (.A(_16984_),
    .B1(_17581_),
    .B2(\core.keymem.key_mem[14][32] ),
    .ZN(_17774_));
 NAND4_X2 _23862_ (.A1(_17770_),
    .A2(_17772_),
    .A3(_17773_),
    .A4(_17774_),
    .ZN(_17775_));
 NOR2_X4 _23863_ (.A1(_17767_),
    .A2(_17775_),
    .ZN(_17776_));
 AND2_X2 _23864_ (.A1(_00265_),
    .A2(_17578_),
    .ZN(_17777_));
 NOR2_X4 _23865_ (.A1(_17776_),
    .A2(_17777_),
    .ZN(_17778_));
 XNOR2_X2 _23866_ (.A(\core.dec_block.block_w2_reg[0] ),
    .B(_17778_),
    .ZN(_17779_));
 XNOR2_X2 _23867_ (.A(_17762_),
    .B(_17779_),
    .ZN(_17780_));
 BUF_X4 _23868_ (.A(_16452_),
    .Z(_17781_));
 AOI22_X1 _23869_ (.A1(\core.keymem.key_mem[4][57] ),
    .A2(_16500_),
    .B1(_17781_),
    .B2(\core.keymem.key_mem[8][57] ),
    .ZN(_17782_));
 AOI22_X2 _23870_ (.A1(\core.keymem.key_mem[3][57] ),
    .A2(_16987_),
    .B1(_17668_),
    .B2(\core.keymem.key_mem[9][57] ),
    .ZN(_17783_));
 BUF_X4 _23871_ (.A(_17193_),
    .Z(_17784_));
 AOI22_X2 _23872_ (.A1(\core.keymem.key_mem[10][57] ),
    .A2(_16989_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][57] ),
    .ZN(_17785_));
 BUF_X8 _23873_ (.A(_16993_),
    .Z(_17786_));
 AOI22_X2 _23874_ (.A1(\core.keymem.key_mem[2][57] ),
    .A2(_17786_),
    .B1(_17720_),
    .B2(\core.keymem.key_mem[12][57] ),
    .ZN(_17787_));
 NAND4_X2 _23875_ (.A1(_17782_),
    .A2(_17783_),
    .A3(_17785_),
    .A4(_17787_),
    .ZN(_17788_));
 BUF_X4 _23876_ (.A(_16407_),
    .Z(_17789_));
 AOI22_X1 _23877_ (.A1(\core.keymem.key_mem[7][57] ),
    .A2(_17789_),
    .B1(_17008_),
    .B2(\core.keymem.key_mem[11][57] ),
    .ZN(_17790_));
 AOI22_X2 _23878_ (.A1(\core.keymem.key_mem[6][57] ),
    .A2(_16521_),
    .B1(_17003_),
    .B2(\core.keymem.key_mem[1][57] ),
    .ZN(_17791_));
 AOI22_X2 _23879_ (.A1(\core.keymem.key_mem[14][57] ),
    .A2(_16999_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][57] ),
    .ZN(_17792_));
 NAND3_X2 _23880_ (.A1(_17790_),
    .A2(_17791_),
    .A3(_17792_),
    .ZN(_17793_));
 NOR3_X4 _23881_ (.A1(_16984_),
    .A2(_17788_),
    .A3(_17793_),
    .ZN(_17794_));
 AOI21_X4 _23882_ (.A(_17794_),
    .B1(_16548_),
    .B2(_00269_),
    .ZN(_17795_));
 XNOR2_X2 _23883_ (.A(\core.dec_block.block_w2_reg[25] ),
    .B(_17795_),
    .ZN(_17796_));
 XNOR2_X2 _23884_ (.A(_17604_),
    .B(_17796_),
    .ZN(_17797_));
 XNOR2_X2 _23885_ (.A(_17780_),
    .B(_17797_),
    .ZN(_17798_));
 INV_X1 _23886_ (.A(\core.dec_block.block_w2_reg[19] ),
    .ZN(_17799_));
 NAND2_X1 _23887_ (.A1(_00285_),
    .A2(_17014_),
    .ZN(_17800_));
 AOI22_X1 _23888_ (.A1(\core.keymem.key_mem[10][51] ),
    .A2(_16514_),
    .B1(_16854_),
    .B2(\core.keymem.key_mem[1][51] ),
    .ZN(_17801_));
 AOI22_X1 _23889_ (.A1(\core.keymem.key_mem[3][51] ),
    .A2(_16865_),
    .B1(_16461_),
    .B2(\core.keymem.key_mem[9][51] ),
    .ZN(_17802_));
 AOI22_X1 _23890_ (.A1(\core.keymem.key_mem[7][51] ),
    .A2(_16955_),
    .B1(_16948_),
    .B2(\core.keymem.key_mem[5][51] ),
    .ZN(_17803_));
 AOI22_X1 _23891_ (.A1(\core.keymem.key_mem[4][51] ),
    .A2(_16946_),
    .B1(_16397_),
    .B2(\core.keymem.key_mem[12][51] ),
    .ZN(_17804_));
 AND4_X1 _23892_ (.A1(_17801_),
    .A2(_17802_),
    .A3(_17803_),
    .A4(_17804_),
    .ZN(_17805_));
 AOI22_X2 _23893_ (.A1(\core.keymem.key_mem[6][51] ),
    .A2(_17695_),
    .B1(_16442_),
    .B2(\core.keymem.key_mem[11][51] ),
    .ZN(_17806_));
 AOI22_X2 _23894_ (.A1(\core.keymem.key_mem[2][51] ),
    .A2(_16860_),
    .B1(_16529_),
    .B2(\core.keymem.key_mem[8][51] ),
    .ZN(_17807_));
 AOI22_X4 _23895_ (.A1(\core.keymem.key_mem[14][51] ),
    .A2(_16438_),
    .B1(_16532_),
    .B2(\core.keymem.key_mem[13][51] ),
    .ZN(_17808_));
 NAND4_X4 _23896_ (.A1(_17805_),
    .A2(_17806_),
    .A3(_17807_),
    .A4(_17808_),
    .ZN(_17809_));
 OAI21_X4 _23897_ (.A(_17800_),
    .B1(_17809_),
    .B2(_16872_),
    .ZN(_17810_));
 XNOR2_X2 _23898_ (.A(_17799_),
    .B(_17810_),
    .ZN(_17811_));
 XNOR2_X1 _23899_ (.A(_17703_),
    .B(_17811_),
    .ZN(_17812_));
 XNOR2_X2 _23900_ (.A(_17798_),
    .B(_17812_),
    .ZN(_17813_));
 AOI21_X1 _23901_ (.A(_16494_),
    .B1(_16949_),
    .B2(\core.keymem.key_mem[5][45] ),
    .ZN(_17814_));
 AOI22_X1 _23902_ (.A1(\core.keymem.key_mem[14][45] ),
    .A2(_17191_),
    .B1(_17648_),
    .B2(\core.keymem.key_mem[6][45] ),
    .ZN(_17815_));
 AOI22_X1 _23903_ (.A1(\core.keymem.key_mem[9][45] ),
    .A2(_17522_),
    .B1(_17000_),
    .B2(\core.keymem.key_mem[12][45] ),
    .ZN(_17816_));
 AOI22_X1 _23904_ (.A1(\core.keymem.key_mem[11][45] ),
    .A2(_17007_),
    .B1(_17193_),
    .B2(\core.keymem.key_mem[13][45] ),
    .ZN(_17817_));
 AND4_X1 _23905_ (.A1(_17814_),
    .A2(_17815_),
    .A3(_17816_),
    .A4(_17817_),
    .ZN(_17818_));
 AOI222_X2 _23906_ (.A1(\core.keymem.key_mem[7][45] ),
    .A2(_17736_),
    .B1(_16423_),
    .B2(\core.keymem.key_mem[2][45] ),
    .C1(_16385_),
    .C2(\core.keymem.key_mem[3][45] ),
    .ZN(_17819_));
 AOI22_X1 _23907_ (.A1(\core.keymem.key_mem[8][45] ),
    .A2(_17506_),
    .B1(_16988_),
    .B2(\core.keymem.key_mem[10][45] ),
    .ZN(_17820_));
 AOI22_X1 _23908_ (.A1(\core.keymem.key_mem[4][45] ),
    .A2(_16499_),
    .B1(_16524_),
    .B2(\core.keymem.key_mem[1][45] ),
    .ZN(_17821_));
 AND3_X1 _23909_ (.A1(_17819_),
    .A2(_17820_),
    .A3(_17821_),
    .ZN(_17822_));
 AOI22_X4 _23910_ (.A1(_00260_),
    .A2(_17014_),
    .B1(_17818_),
    .B2(_17822_),
    .ZN(_17823_));
 XNOR2_X2 _23911_ (.A(\core.dec_block.block_w2_reg[13] ),
    .B(_17823_),
    .ZN(_17824_));
 AND2_X1 _23912_ (.A1(_00261_),
    .A2(_16982_),
    .ZN(_17825_));
 NAND3_X1 _23913_ (.A1(\core.keymem.key_mem[14][47] ),
    .A2(_16882_),
    .A3(_17156_),
    .ZN(_17826_));
 BUF_X4 _23914_ (.A(_16969_),
    .Z(_17827_));
 OAI211_X2 _23915_ (.A(\core.keymem.key_mem[1][47] ),
    .B(_17827_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_17828_));
 OAI221_X2 _23916_ (.A(\core.keymem.key_mem[5][47] ),
    .B1(_16908_),
    .B2(_16917_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_17829_));
 OAI211_X2 _23917_ (.A(\core.keymem.key_mem[6][47] ),
    .B(_17026_),
    .C1(_17622_),
    .C2(_17030_),
    .ZN(_17830_));
 NAND4_X2 _23918_ (.A1(_17826_),
    .A2(_17828_),
    .A3(_17829_),
    .A4(_17830_),
    .ZN(_17831_));
 NAND3_X1 _23919_ (.A1(\core.keymem.key_mem[3][47] ),
    .A2(_17074_),
    .A3(_17827_),
    .ZN(_17832_));
 NAND3_X1 _23920_ (.A1(\core.keymem.key_mem[2][47] ),
    .A2(_17827_),
    .A3(_17163_),
    .ZN(_17833_));
 OAI211_X2 _23921_ (.A(\core.keymem.key_mem[7][47] ),
    .B(_16901_),
    .C1(_16896_),
    .C2(_16899_),
    .ZN(_17834_));
 OAI211_X2 _23922_ (.A(\core.keymem.key_mem[4][47] ),
    .B(_16893_),
    .C1(_16896_),
    .C2(_16899_),
    .ZN(_17835_));
 NAND4_X2 _23923_ (.A1(_17832_),
    .A2(_17833_),
    .A3(_17834_),
    .A4(_17835_),
    .ZN(_17836_));
 OAI211_X2 _23924_ (.A(\core.keymem.key_mem[8][47] ),
    .B(_16893_),
    .C1(_16927_),
    .C2(_16929_),
    .ZN(_17837_));
 OAI211_X2 _23925_ (.A(\core.keymem.key_mem[11][47] ),
    .B(_16901_),
    .C1(_16927_),
    .C2(_16929_),
    .ZN(_17838_));
 OAI221_X2 _23926_ (.A(\core.keymem.key_mem[9][47] ),
    .B1(_16885_),
    .B2(_16889_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_17839_));
 OAI211_X2 _23927_ (.A(\core.keymem.key_mem[13][47] ),
    .B(_16919_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_17840_));
 NAND4_X2 _23928_ (.A1(_17837_),
    .A2(_17838_),
    .A3(_17839_),
    .A4(_17840_),
    .ZN(_17841_));
 INV_X1 _23929_ (.A(\core.keymem.key_mem[10][47] ),
    .ZN(_17842_));
 NAND2_X4 _23930_ (.A1(_16881_),
    .A2(_16921_),
    .ZN(_17843_));
 INV_X1 _23931_ (.A(\core.keymem.key_mem[12][47] ),
    .ZN(_17844_));
 OAI22_X4 _23932_ (.A1(_17842_),
    .A2(_17038_),
    .B1(_17843_),
    .B2(_17844_),
    .ZN(_17845_));
 NOR4_X4 _23933_ (.A1(_17831_),
    .A2(_17836_),
    .A3(_17841_),
    .A4(_17845_),
    .ZN(_17846_));
 AOI21_X4 _23934_ (.A(_17825_),
    .B1(_17846_),
    .B2(_16488_),
    .ZN(_17847_));
 XNOR2_X2 _23935_ (.A(\core.dec_block.block_w2_reg[15] ),
    .B(_17847_),
    .ZN(_17848_));
 XNOR2_X1 _23936_ (.A(_17824_),
    .B(_17848_),
    .ZN(_17849_));
 XNOR2_X2 _23937_ (.A(_17618_),
    .B(_17849_),
    .ZN(_17850_));
 NAND2_X1 _23938_ (.A1(_00284_),
    .A2(_17014_),
    .ZN(_17851_));
 AOI22_X1 _23939_ (.A1(\core.keymem.key_mem[14][35] ),
    .A2(_17191_),
    .B1(_16415_),
    .B2(\core.keymem.key_mem[1][35] ),
    .ZN(_17852_));
 AOI22_X1 _23940_ (.A1(\core.keymem.key_mem[4][35] ),
    .A2(_16946_),
    .B1(_16423_),
    .B2(\core.keymem.key_mem[2][35] ),
    .ZN(_17853_));
 AOI22_X1 _23941_ (.A1(\core.keymem.key_mem[8][35] ),
    .A2(_16451_),
    .B1(_16385_),
    .B2(\core.keymem.key_mem[3][35] ),
    .ZN(_17854_));
 AOI22_X1 _23942_ (.A1(\core.keymem.key_mem[6][35] ),
    .A2(_16447_),
    .B1(_16441_),
    .B2(\core.keymem.key_mem[11][35] ),
    .ZN(_17855_));
 AND4_X1 _23943_ (.A1(_17852_),
    .A2(_17853_),
    .A3(_17854_),
    .A4(_17855_),
    .ZN(_17856_));
 AOI22_X2 _23944_ (.A1(\core.keymem.key_mem[10][35] ),
    .A2(_17715_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][35] ),
    .ZN(_17857_));
 AOI22_X2 _23945_ (.A1(\core.keymem.key_mem[9][35] ),
    .A2(_16536_),
    .B1(_16532_),
    .B2(\core.keymem.key_mem[13][35] ),
    .ZN(_17858_));
 AOI22_X4 _23946_ (.A1(\core.keymem.key_mem[7][35] ),
    .A2(_16512_),
    .B1(_16398_),
    .B2(\core.keymem.key_mem[12][35] ),
    .ZN(_17859_));
 NAND4_X4 _23947_ (.A1(_17856_),
    .A2(_17857_),
    .A3(_17858_),
    .A4(_17859_),
    .ZN(_17860_));
 OAI21_X4 _23948_ (.A(_17851_),
    .B1(_17860_),
    .B2(_16872_),
    .ZN(_17861_));
 XOR2_X2 _23949_ (.A(\core.dec_block.block_w2_reg[3] ),
    .B(_17861_),
    .Z(_17862_));
 XNOR2_X1 _23950_ (.A(_17850_),
    .B(_17862_),
    .ZN(_17863_));
 INV_X1 _23951_ (.A(\core.dec_block.block_w2_reg[10] ),
    .ZN(_17864_));
 XNOR2_X2 _23952_ (.A(_17864_),
    .B(_17727_),
    .ZN(_17865_));
 XNOR2_X2 _23953_ (.A(_17848_),
    .B(_17865_),
    .ZN(_17866_));
 XOR2_X1 _23954_ (.A(_17536_),
    .B(_17866_),
    .Z(_17867_));
 XNOR2_X1 _23955_ (.A(_17863_),
    .B(_17867_),
    .ZN(_17868_));
 AND2_X1 _23956_ (.A1(_00257_),
    .A2(_16871_),
    .ZN(_17869_));
 OAI211_X2 _23957_ (.A(\core.keymem.key_mem[6][53] ),
    .B(_17016_),
    .C1(_17115_),
    .C2(_17146_),
    .ZN(_17870_));
 NAND3_X1 _23958_ (.A1(\core.keymem.key_mem[3][53] ),
    .A2(_17048_),
    .A3(_16970_),
    .ZN(_17871_));
 OAI211_X2 _23959_ (.A(\core.keymem.key_mem[1][53] ),
    .B(_17120_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_17872_));
 NAND3_X1 _23960_ (.A1(\core.keymem.key_mem[12][53] ),
    .A2(_16882_),
    .A3(_17527_),
    .ZN(_17873_));
 NAND4_X2 _23961_ (.A1(_17870_),
    .A2(_17871_),
    .A3(_17872_),
    .A4(_17873_),
    .ZN(_17874_));
 OAI211_X2 _23962_ (.A(\core.keymem.key_mem[7][53] ),
    .B(_17111_),
    .C1(_17146_),
    .C2(_17622_),
    .ZN(_17875_));
 OAI221_X2 _23963_ (.A(\core.keymem.key_mem[5][53] ),
    .B1(_16896_),
    .B2(_16899_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_17876_));
 NAND3_X1 _23964_ (.A1(\core.keymem.key_mem[14][53] ),
    .A2(_17024_),
    .A3(_17026_),
    .ZN(_17877_));
 OAI211_X2 _23965_ (.A(\core.keymem.key_mem[4][53] ),
    .B(_17028_),
    .C1(_17030_),
    .C2(_17031_),
    .ZN(_17878_));
 NAND4_X2 _23966_ (.A1(_17875_),
    .A2(_17876_),
    .A3(_17877_),
    .A4(_17878_),
    .ZN(_17879_));
 OAI211_X2 _23967_ (.A(\core.keymem.key_mem[8][53] ),
    .B(_17028_),
    .C1(_17035_),
    .C2(_17036_),
    .ZN(_17880_));
 OAI211_X2 _23968_ (.A(\core.keymem.key_mem[13][53] ),
    .B(_17099_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_17881_));
 OAI211_X2 _23969_ (.A(\core.keymem.key_mem[11][53] ),
    .B(_17074_),
    .C1(_17035_),
    .C2(_17036_),
    .ZN(_17882_));
 OAI221_X2 _23970_ (.A(\core.keymem.key_mem[9][53] ),
    .B1(_16922_),
    .B2(_16923_),
    .C1(_16913_),
    .C2(_16915_),
    .ZN(_17883_));
 NAND4_X2 _23971_ (.A1(_17880_),
    .A2(_17881_),
    .A3(_17882_),
    .A4(_17883_),
    .ZN(_17884_));
 INV_X1 _23972_ (.A(\core.keymem.key_mem[2][53] ),
    .ZN(_17885_));
 NAND2_X2 _23973_ (.A1(_16969_),
    .A2(_17015_),
    .ZN(_17886_));
 INV_X1 _23974_ (.A(\core.keymem.key_mem[10][53] ),
    .ZN(_17887_));
 OAI22_X2 _23975_ (.A1(_17885_),
    .A2(_17886_),
    .B1(_17038_),
    .B2(_17887_),
    .ZN(_17888_));
 NOR4_X4 _23976_ (.A1(_17874_),
    .A2(_17879_),
    .A3(_17884_),
    .A4(_17888_),
    .ZN(_17889_));
 AOI21_X4 _23977_ (.A(_17869_),
    .B1(_17889_),
    .B2(_17533_),
    .ZN(_17890_));
 XNOR2_X2 _23978_ (.A(\core.dec_block.block_w2_reg[21] ),
    .B(_17890_),
    .ZN(_17891_));
 INV_X1 _23979_ (.A(\core.dec_block.block_w2_reg[16] ),
    .ZN(_17892_));
 AOI22_X1 _23980_ (.A1(\core.keymem.key_mem[7][48] ),
    .A2(_17084_),
    .B1(_17666_),
    .B2(\core.keymem.key_mem[8][48] ),
    .ZN(_17893_));
 AOI22_X1 _23981_ (.A1(\core.keymem.key_mem[12][48] ),
    .A2(_17720_),
    .B1(_16855_),
    .B2(\core.keymem.key_mem[1][48] ),
    .ZN(_17894_));
 AOI22_X1 _23982_ (.A1(\core.keymem.key_mem[3][48] ),
    .A2(_16866_),
    .B1(_16506_),
    .B2(\core.keymem.key_mem[11][48] ),
    .ZN(_17895_));
 AOI22_X1 _23983_ (.A1(\core.keymem.key_mem[9][48] ),
    .A2(_17668_),
    .B1(_16515_),
    .B2(\core.keymem.key_mem[10][48] ),
    .ZN(_17896_));
 NAND4_X1 _23984_ (.A1(_17893_),
    .A2(_17894_),
    .A3(_17895_),
    .A4(_17896_),
    .ZN(_17897_));
 NAND3_X1 _23985_ (.A1(\core.keymem.key_mem[4][48] ),
    .A2(_17057_),
    .A3(_16967_),
    .ZN(_17898_));
 NAND3_X1 _23986_ (.A1(\core.keymem.key_mem[14][48] ),
    .A2(_17101_),
    .A3(_17055_),
    .ZN(_17899_));
 AOI21_X1 _23987_ (.A(_17043_),
    .B1(_17898_),
    .B2(_17899_),
    .ZN(_17900_));
 AOI22_X1 _23988_ (.A1(\core.keymem.key_mem[6][48] ),
    .A2(_17695_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][48] ),
    .ZN(_17901_));
 AOI22_X1 _23989_ (.A1(\core.keymem.key_mem[2][48] ),
    .A2(_16860_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][48] ),
    .ZN(_17902_));
 NAND2_X1 _23990_ (.A1(_17901_),
    .A2(_17902_),
    .ZN(_17903_));
 NOR3_X1 _23991_ (.A1(_17897_),
    .A2(_17900_),
    .A3(_17903_),
    .ZN(_17904_));
 MUX2_X2 _23992_ (.A(_00266_),
    .B(_17904_),
    .S(_16489_),
    .Z(_17905_));
 XNOR2_X2 _23993_ (.A(_17892_),
    .B(_17905_),
    .ZN(_17906_));
 XNOR2_X2 _23994_ (.A(_17891_),
    .B(_17906_),
    .ZN(_17907_));
 XNOR2_X2 _23995_ (.A(_17552_),
    .B(_17907_),
    .ZN(_17908_));
 INV_X1 _23996_ (.A(\core.dec_block.block_w2_reg[27] ),
    .ZN(_17909_));
 NAND2_X1 _23997_ (.A1(_00282_),
    .A2(_16498_),
    .ZN(_17910_));
 AOI22_X1 _23998_ (.A1(\core.keymem.key_mem[3][59] ),
    .A2(_17683_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][59] ),
    .ZN(_17911_));
 AOI22_X1 _23999_ (.A1(\core.keymem.key_mem[6][59] ),
    .A2(_16991_),
    .B1(_17003_),
    .B2(\core.keymem.key_mem[1][59] ),
    .ZN(_17912_));
 AOI22_X1 _24000_ (.A1(\core.keymem.key_mem[4][59] ),
    .A2(_16500_),
    .B1(_17789_),
    .B2(\core.keymem.key_mem[7][59] ),
    .ZN(_17913_));
 BUF_X4 _24001_ (.A(_17522_),
    .Z(_17914_));
 AOI22_X1 _24002_ (.A1(\core.keymem.key_mem[2][59] ),
    .A2(_16994_),
    .B1(_17914_),
    .B2(\core.keymem.key_mem[9][59] ),
    .ZN(_17915_));
 AND4_X1 _24003_ (.A1(_17911_),
    .A2(_17912_),
    .A3(_17913_),
    .A4(_17915_),
    .ZN(_17916_));
 AOI22_X2 _24004_ (.A1(\core.keymem.key_mem[10][59] ),
    .A2(_17082_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][59] ),
    .ZN(_17917_));
 AOI22_X4 _24005_ (.A1(\core.keymem.key_mem[14][59] ),
    .A2(_17581_),
    .B1(_17769_),
    .B2(\core.keymem.key_mem[11][59] ),
    .ZN(_17918_));
 AOI22_X4 _24006_ (.A1(\core.keymem.key_mem[8][59] ),
    .A2(_17765_),
    .B1(_17093_),
    .B2(\core.keymem.key_mem[12][59] ),
    .ZN(_17919_));
 NAND4_X4 _24007_ (.A1(_17916_),
    .A2(_17917_),
    .A3(_17918_),
    .A4(_17919_),
    .ZN(_17920_));
 OAI21_X4 _24008_ (.A(_17910_),
    .B1(_17920_),
    .B2(_16498_),
    .ZN(_17921_));
 XNOR2_X2 _24009_ (.A(_17909_),
    .B(_17921_),
    .ZN(_17922_));
 INV_X1 _24010_ (.A(\core.dec_block.block_w2_reg[31] ),
    .ZN(_17923_));
 NAND2_X1 _24011_ (.A1(_00276_),
    .A2(_16872_),
    .ZN(_17924_));
 AOI22_X1 _24012_ (.A1(\core.keymem.key_mem[12][63] ),
    .A2(_17000_),
    .B1(_16854_),
    .B2(\core.keymem.key_mem[1][63] ),
    .ZN(_17925_));
 AOI22_X1 _24013_ (.A1(\core.keymem.key_mem[2][63] ),
    .A2(_16859_),
    .B1(_16531_),
    .B2(\core.keymem.key_mem[13][63] ),
    .ZN(_17926_));
 AOI22_X1 _24014_ (.A1(\core.keymem.key_mem[7][63] ),
    .A2(_16955_),
    .B1(_16467_),
    .B2(\core.keymem.key_mem[5][63] ),
    .ZN(_17927_));
 AOI22_X1 _24015_ (.A1(\core.keymem.key_mem[4][63] ),
    .A2(_16456_),
    .B1(_16437_),
    .B2(\core.keymem.key_mem[14][63] ),
    .ZN(_17928_));
 AND4_X1 _24016_ (.A1(_17925_),
    .A2(_17926_),
    .A3(_17927_),
    .A4(_17928_),
    .ZN(_17929_));
 AOI22_X2 _24017_ (.A1(\core.keymem.key_mem[6][63] ),
    .A2(_17695_),
    .B1(_17715_),
    .B2(\core.keymem.key_mem[10][63] ),
    .ZN(_17930_));
 AOI22_X2 _24018_ (.A1(\core.keymem.key_mem[9][63] ),
    .A2(_16536_),
    .B1(_16506_),
    .B2(\core.keymem.key_mem[11][63] ),
    .ZN(_17931_));
 AOI22_X4 _24019_ (.A1(\core.keymem.key_mem[8][63] ),
    .A2(_16529_),
    .B1(_16386_),
    .B2(\core.keymem.key_mem[3][63] ),
    .ZN(_17932_));
 NAND4_X4 _24020_ (.A1(_17929_),
    .A2(_17930_),
    .A3(_17931_),
    .A4(_17932_),
    .ZN(_17933_));
 OAI21_X4 _24021_ (.A(_17924_),
    .B1(_17933_),
    .B2(_16872_),
    .ZN(_17934_));
 XNOR2_X2 _24022_ (.A(_17923_),
    .B(_17934_),
    .ZN(_17935_));
 AOI22_X1 _24023_ (.A1(\core.keymem.key_mem[4][61] ),
    .A2(_16946_),
    .B1(_16514_),
    .B2(\core.keymem.key_mem[10][61] ),
    .ZN(_17936_));
 AOI21_X1 _24024_ (.A(_16544_),
    .B1(_16437_),
    .B2(\core.keymem.key_mem[14][61] ),
    .ZN(_17937_));
 AOI22_X1 _24025_ (.A1(\core.keymem.key_mem[1][61] ),
    .A2(_16415_),
    .B1(_16948_),
    .B2(\core.keymem.key_mem[5][61] ),
    .ZN(_17938_));
 AOI22_X1 _24026_ (.A1(\core.keymem.key_mem[7][61] ),
    .A2(_16406_),
    .B1(_16397_),
    .B2(\core.keymem.key_mem[12][61] ),
    .ZN(_17939_));
 AND4_X1 _24027_ (.A1(_17936_),
    .A2(_17937_),
    .A3(_17938_),
    .A4(_17939_),
    .ZN(_17940_));
 AOI222_X2 _24028_ (.A1(\core.keymem.key_mem[6][61] ),
    .A2(_16447_),
    .B1(_16864_),
    .B2(\core.keymem.key_mem[3][61] ),
    .C1(_16471_),
    .C2(\core.keymem.key_mem[13][61] ),
    .ZN(_17941_));
 AOI22_X1 _24029_ (.A1(\core.keymem.key_mem[8][61] ),
    .A2(_16451_),
    .B1(_16441_),
    .B2(\core.keymem.key_mem[11][61] ),
    .ZN(_17942_));
 AOI22_X1 _24030_ (.A1(\core.keymem.key_mem[2][61] ),
    .A2(_16423_),
    .B1(_16461_),
    .B2(\core.keymem.key_mem[9][61] ),
    .ZN(_17943_));
 AND3_X1 _24031_ (.A1(_17941_),
    .A2(_17942_),
    .A3(_17943_),
    .ZN(_17944_));
 AOI22_X4 _24032_ (.A1(_00255_),
    .A2(_16983_),
    .B1(_17940_),
    .B2(_17944_),
    .ZN(_17945_));
 XNOR2_X2 _24033_ (.A(\core.dec_block.block_w2_reg[29] ),
    .B(_17945_),
    .ZN(_17946_));
 XNOR2_X2 _24034_ (.A(_17643_),
    .B(_17946_),
    .ZN(_17947_));
 XNOR2_X2 _24035_ (.A(_17935_),
    .B(_17947_),
    .ZN(_17948_));
 XNOR2_X1 _24036_ (.A(_17922_),
    .B(_17948_),
    .ZN(_17949_));
 XNOR2_X2 _24037_ (.A(_17908_),
    .B(_17949_),
    .ZN(_17950_));
 XNOR2_X1 _24038_ (.A(_17868_),
    .B(_17950_),
    .ZN(_17951_));
 XNOR2_X1 _24039_ (.A(_17813_),
    .B(_17951_),
    .ZN(_17952_));
 NAND2_X1 _24040_ (.A1(_17749_),
    .A2(_17952_),
    .ZN(_17953_));
 NOR2_X1 _24041_ (.A1(_17467_),
    .A2(_17440_),
    .ZN(_17954_));
 NAND2_X4 _24042_ (.A1(_17263_),
    .A2(_17380_),
    .ZN(_17955_));
 AOI21_X1 _24043_ (.A(_17308_),
    .B1(_17459_),
    .B2(_17955_),
    .ZN(_17956_));
 OAI21_X1 _24044_ (.A(_17374_),
    .B1(_17954_),
    .B2(_17956_),
    .ZN(_17957_));
 AOI22_X2 _24045_ (.A1(_17351_),
    .A2(_17360_),
    .B1(_17404_),
    .B2(_17343_),
    .ZN(_17958_));
 OAI21_X2 _24046_ (.A(_17957_),
    .B1(_17958_),
    .B2(_17374_),
    .ZN(_17959_));
 AOI21_X1 _24047_ (.A(_17280_),
    .B1(_17368_),
    .B2(_17448_),
    .ZN(_17960_));
 OAI21_X1 _24048_ (.A(_17381_),
    .B1(_17373_),
    .B2(_17960_),
    .ZN(_17961_));
 NOR3_X1 _24049_ (.A1(_17213_),
    .A2(_17272_),
    .A3(_17486_),
    .ZN(_17962_));
 NOR2_X2 _24050_ (.A1(_17220_),
    .A2(_17418_),
    .ZN(_17963_));
 AOI21_X1 _24051_ (.A(_17962_),
    .B1(_17963_),
    .B2(_17316_),
    .ZN(_17964_));
 BUF_X4 _24052_ (.A(_17268_),
    .Z(_17965_));
 OAI21_X1 _24053_ (.A(_17961_),
    .B1(_17964_),
    .B2(_17965_),
    .ZN(_17966_));
 AOI21_X1 _24054_ (.A(_17399_),
    .B1(_17397_),
    .B2(_17437_),
    .ZN(_17967_));
 NOR2_X2 _24055_ (.A1(_17211_),
    .A2(_17269_),
    .ZN(_17968_));
 AOI21_X1 _24056_ (.A(_17496_),
    .B1(_17968_),
    .B2(_17350_),
    .ZN(_17969_));
 NOR3_X1 _24057_ (.A1(_17482_),
    .A2(_17268_),
    .A3(_17969_),
    .ZN(_17970_));
 NAND2_X1 _24058_ (.A1(_17445_),
    .A2(_17446_),
    .ZN(_17971_));
 NAND2_X1 _24059_ (.A1(_17471_),
    .A2(_17354_),
    .ZN(_17972_));
 NAND3_X1 _24060_ (.A1(_17408_),
    .A2(_17971_),
    .A3(_17972_),
    .ZN(_17973_));
 NOR4_X2 _24061_ (.A1(_17966_),
    .A2(_17967_),
    .A3(_17970_),
    .A4(_17973_),
    .ZN(_17974_));
 NOR2_X1 _24062_ (.A1(_17270_),
    .A2(_17279_),
    .ZN(_17975_));
 NOR2_X1 _24063_ (.A1(_17479_),
    .A2(_17258_),
    .ZN(_17976_));
 NOR2_X1 _24064_ (.A1(_17276_),
    .A2(_17281_),
    .ZN(_17977_));
 AOI21_X1 _24065_ (.A(_17976_),
    .B1(_17977_),
    .B2(_17482_),
    .ZN(_17978_));
 NOR3_X1 _24066_ (.A1(_17296_),
    .A2(_17288_),
    .A3(_17978_),
    .ZN(_17979_));
 NOR2_X1 _24067_ (.A1(_17372_),
    .A2(_17220_),
    .ZN(_17980_));
 AND4_X1 _24068_ (.A1(_17296_),
    .A2(_17288_),
    .A3(_17285_),
    .A4(_17980_),
    .ZN(_17981_));
 OAI21_X1 _24069_ (.A(_17975_),
    .B1(_17979_),
    .B2(_17981_),
    .ZN(_17982_));
 NAND2_X1 _24070_ (.A1(_17219_),
    .A2(_17264_),
    .ZN(_17983_));
 NOR2_X1 _24071_ (.A1(_17317_),
    .A2(_17983_),
    .ZN(_17984_));
 OAI21_X1 _24072_ (.A(_17437_),
    .B1(_17264_),
    .B2(_17463_),
    .ZN(_17985_));
 AOI221_X2 _24073_ (.A(_17984_),
    .B1(_17492_),
    .B2(_17383_),
    .C1(_17301_),
    .C2(_17985_),
    .ZN(_17986_));
 BUF_X4 _24074_ (.A(_17342_),
    .Z(_17987_));
 OAI33_X1 _24075_ (.A1(_17464_),
    .A2(_17987_),
    .A3(_17418_),
    .B1(_17439_),
    .B2(_17382_),
    .B3(_17322_),
    .ZN(_17988_));
 BUF_X4 _24076_ (.A(_17352_),
    .Z(_17989_));
 NOR2_X1 _24077_ (.A1(_17326_),
    .A2(_17989_),
    .ZN(_17990_));
 NAND3_X1 _24078_ (.A1(_17371_),
    .A2(_17258_),
    .A3(_17377_),
    .ZN(_17991_));
 OAI21_X1 _24079_ (.A(_17991_),
    .B1(_17314_),
    .B2(_17258_),
    .ZN(_17992_));
 NOR2_X2 _24080_ (.A1(_17296_),
    .A2(_17322_),
    .ZN(_17993_));
 AOI221_X2 _24081_ (.A(_17988_),
    .B1(_17990_),
    .B2(_17414_),
    .C1(_17992_),
    .C2(_17993_),
    .ZN(_17994_));
 NAND4_X2 _24082_ (.A1(_17974_),
    .A2(_17982_),
    .A3(_17986_),
    .A4(_17994_),
    .ZN(_17995_));
 NOR2_X2 _24083_ (.A1(_17393_),
    .A2(_17342_),
    .ZN(_17996_));
 OAI21_X1 _24084_ (.A(_17996_),
    .B1(_17350_),
    .B2(_17300_),
    .ZN(_17997_));
 NOR3_X1 _24085_ (.A1(_17276_),
    .A2(_17279_),
    .A3(_17352_),
    .ZN(_17998_));
 NOR3_X1 _24086_ (.A1(_17258_),
    .A2(_17267_),
    .A3(_17458_),
    .ZN(_17999_));
 NOR2_X1 _24087_ (.A1(_17998_),
    .A2(_17999_),
    .ZN(_18000_));
 NOR3_X1 _24088_ (.A1(_17316_),
    .A2(_17365_),
    .A3(_18000_),
    .ZN(_18001_));
 MUX2_X1 _24089_ (.A(_17494_),
    .B(_17496_),
    .S(_17479_),
    .Z(_18002_));
 NOR2_X2 _24090_ (.A1(_17228_),
    .A2(_17267_),
    .ZN(_18003_));
 AOI21_X1 _24091_ (.A(_18001_),
    .B1(_18002_),
    .B2(_18003_),
    .ZN(_18004_));
 NOR2_X4 _24092_ (.A1(_17265_),
    .A2(_17352_),
    .ZN(_18005_));
 NOR2_X1 _24093_ (.A1(_17227_),
    .A2(_17393_),
    .ZN(_18006_));
 OAI33_X1 _24094_ (.A1(_17213_),
    .A2(_17280_),
    .A3(_17448_),
    .B1(_17488_),
    .B2(_18006_),
    .B3(_17310_),
    .ZN(_18007_));
 AOI22_X2 _24095_ (.A1(_17346_),
    .A2(_18005_),
    .B1(_18007_),
    .B2(_17482_),
    .ZN(_18008_));
 NAND3_X2 _24096_ (.A1(_17997_),
    .A2(_18004_),
    .A3(_18008_),
    .ZN(_18009_));
 NAND2_X1 _24097_ (.A1(_17270_),
    .A2(_17456_),
    .ZN(_18010_));
 NAND2_X1 _24098_ (.A1(_17227_),
    .A2(_17491_),
    .ZN(_18011_));
 AOI21_X1 _24099_ (.A(_17358_),
    .B1(_18010_),
    .B2(_18011_),
    .ZN(_18012_));
 OAI22_X1 _24100_ (.A1(_17955_),
    .A2(_17429_),
    .B1(_17474_),
    .B2(_17358_),
    .ZN(_18013_));
 NOR2_X4 _24101_ (.A1(_17323_),
    .A2(_17436_),
    .ZN(_18014_));
 AOI221_X2 _24102_ (.A(_18012_),
    .B1(_18013_),
    .B2(_17371_),
    .C1(_17300_),
    .C2(_18014_),
    .ZN(_18015_));
 OAI21_X1 _24103_ (.A(_17414_),
    .B1(_17492_),
    .B2(_18014_),
    .ZN(_18016_));
 BUF_X4 _24104_ (.A(_17479_),
    .Z(_18017_));
 NAND2_X1 _24105_ (.A1(_17270_),
    .A2(_17255_),
    .ZN(_18018_));
 OAI21_X1 _24106_ (.A(_18018_),
    .B1(_17468_),
    .B2(_17273_),
    .ZN(_18019_));
 NAND3_X1 _24107_ (.A1(_18017_),
    .A2(_17325_),
    .A3(_18019_),
    .ZN(_18020_));
 NOR3_X1 _24108_ (.A1(_17482_),
    .A2(_17324_),
    .A3(_17486_),
    .ZN(_18021_));
 OAI21_X1 _24109_ (.A(_17273_),
    .B1(_17963_),
    .B2(_18021_),
    .ZN(_18022_));
 NAND4_X2 _24110_ (.A1(_18015_),
    .A2(_18016_),
    .A3(_18020_),
    .A4(_18022_),
    .ZN(_18023_));
 NOR4_X4 _24111_ (.A1(_17959_),
    .A2(_17995_),
    .A3(_18009_),
    .A4(_18023_),
    .ZN(_18024_));
 NAND4_X1 _24112_ (.A1(_17258_),
    .A2(_17239_),
    .A3(_17281_),
    .A4(_17325_),
    .ZN(_18025_));
 XNOR2_X1 _24113_ (.A(_17212_),
    .B(_17258_),
    .ZN(_18026_));
 NOR4_X1 _24114_ (.A1(_17239_),
    .A2(_17281_),
    .A3(_17319_),
    .A4(_18026_),
    .ZN(_18027_));
 OAI22_X1 _24115_ (.A1(_17214_),
    .A2(_17240_),
    .B1(_17339_),
    .B2(_17393_),
    .ZN(_18028_));
 AOI21_X1 _24116_ (.A(_18027_),
    .B1(_18028_),
    .B2(_17281_),
    .ZN(_18029_));
 OAI21_X1 _24117_ (.A(_18025_),
    .B1(_18029_),
    .B2(_17288_),
    .ZN(_18030_));
 NAND2_X1 _24118_ (.A1(_17321_),
    .A2(_18030_),
    .ZN(_18031_));
 NAND2_X2 _24119_ (.A1(_17325_),
    .A2(_17301_),
    .ZN(_18032_));
 OAI21_X2 _24120_ (.A(_18031_),
    .B1(_18032_),
    .B2(_17397_),
    .ZN(_18033_));
 INV_X1 _24121_ (.A(_18033_),
    .ZN(_18034_));
 NOR2_X2 _24122_ (.A1(_17270_),
    .A2(_17441_),
    .ZN(_18035_));
 NAND2_X2 _24123_ (.A1(_17211_),
    .A2(_17227_),
    .ZN(_18036_));
 OAI22_X4 _24124_ (.A1(_17228_),
    .A2(_17324_),
    .B1(_18036_),
    .B2(_17266_),
    .ZN(_18037_));
 NAND2_X2 _24125_ (.A1(_17270_),
    .A2(_17494_),
    .ZN(_18038_));
 OAI21_X1 _24126_ (.A(_17228_),
    .B1(_17255_),
    .B2(_17491_),
    .ZN(_18039_));
 NAND2_X1 _24127_ (.A1(_18038_),
    .A2(_18039_),
    .ZN(_18040_));
 AOI221_X2 _24128_ (.A(_18035_),
    .B1(_18037_),
    .B2(_17456_),
    .C1(_18040_),
    .C2(_17433_),
    .ZN(_18041_));
 NOR2_X2 _24129_ (.A1(_18017_),
    .A2(_18041_),
    .ZN(_18042_));
 NAND3_X1 _24130_ (.A1(_17273_),
    .A2(_17326_),
    .A3(_17404_),
    .ZN(_18043_));
 NAND2_X1 _24131_ (.A1(_17229_),
    .A2(_17366_),
    .ZN(_18044_));
 OAI21_X1 _24132_ (.A(_18043_),
    .B1(_18044_),
    .B2(_17450_),
    .ZN(_18045_));
 AOI21_X1 _24133_ (.A(_17464_),
    .B1(_17310_),
    .B2(_17461_),
    .ZN(_18046_));
 OAI21_X1 _24134_ (.A(_17381_),
    .B1(_17496_),
    .B2(_18046_),
    .ZN(_18047_));
 OAI21_X1 _24135_ (.A(_17482_),
    .B1(_17975_),
    .B2(_18003_),
    .ZN(_18048_));
 OAI221_X2 _24136_ (.A(_18047_),
    .B1(_17436_),
    .B2(_17468_),
    .C1(_17467_),
    .C2(_18048_),
    .ZN(_18049_));
 AOI221_X2 _24137_ (.A(_18042_),
    .B1(_18045_),
    .B2(_18017_),
    .C1(_17214_),
    .C2(_18049_),
    .ZN(_18050_));
 NAND4_X4 _24138_ (.A1(_17378_),
    .A2(_18024_),
    .A3(_18034_),
    .A4(_18050_),
    .ZN(_18051_));
 BUF_X4 _24139_ (.A(_16554_),
    .Z(_18052_));
 NAND2_X1 _24140_ (.A1(_00204_),
    .A2(_17578_),
    .ZN(_18053_));
 AOI22_X1 _24141_ (.A1(\core.keymem.key_mem[6][107] ),
    .A2(_16449_),
    .B1(_16387_),
    .B2(\core.keymem.key_mem[3][107] ),
    .ZN(_18054_));
 AOI22_X1 _24142_ (.A1(\core.keymem.key_mem[7][107] ),
    .A2(_16513_),
    .B1(_16540_),
    .B2(\core.keymem.key_mem[12][107] ),
    .ZN(_18055_));
 AOI22_X1 _24143_ (.A1(\core.keymem.key_mem[8][107] ),
    .A2(_16530_),
    .B1(_17178_),
    .B2(\core.keymem.key_mem[1][107] ),
    .ZN(_18056_));
 AOI22_X1 _24144_ (.A1(\core.keymem.key_mem[5][107] ),
    .A2(_16469_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][107] ),
    .ZN(_18057_));
 AND4_X1 _24145_ (.A1(_18054_),
    .A2(_18055_),
    .A3(_18056_),
    .A4(_18057_),
    .ZN(_18058_));
 AOI22_X2 _24146_ (.A1(\core.keymem.key_mem[9][107] ),
    .A2(_17585_),
    .B1(_17769_),
    .B2(\core.keymem.key_mem[11][107] ),
    .ZN(_18059_));
 AOI22_X2 _24147_ (.A1(\core.keymem.key_mem[4][107] ),
    .A2(_16501_),
    .B1(_17086_),
    .B2(\core.keymem.key_mem[2][107] ),
    .ZN(_18060_));
 AOI22_X2 _24148_ (.A1(\core.keymem.key_mem[14][107] ),
    .A2(_17581_),
    .B1(_17082_),
    .B2(\core.keymem.key_mem[10][107] ),
    .ZN(_18061_));
 NAND4_X2 _24149_ (.A1(_18058_),
    .A2(_18059_),
    .A3(_18060_),
    .A4(_18061_),
    .ZN(_18062_));
 OAI21_X4 _24150_ (.A(_18053_),
    .B1(_18062_),
    .B2(_16549_),
    .ZN(_18063_));
 XNOR2_X2 _24151_ (.A(_17746_),
    .B(_18063_),
    .ZN(_18064_));
 INV_X1 _24152_ (.A(\block_reg[2][11] ),
    .ZN(_18065_));
 AOI22_X1 _24153_ (.A1(\core.keymem.key_mem[7][43] ),
    .A2(_17736_),
    .B1(_16988_),
    .B2(\core.keymem.key_mem[10][43] ),
    .ZN(_18066_));
 AOI22_X1 _24154_ (.A1(\core.keymem.key_mem[2][43] ),
    .A2(_16993_),
    .B1(_16524_),
    .B2(\core.keymem.key_mem[1][43] ),
    .ZN(_18067_));
 AOI22_X1 _24155_ (.A1(\core.keymem.key_mem[8][43] ),
    .A2(_17506_),
    .B1(_17007_),
    .B2(\core.keymem.key_mem[11][43] ),
    .ZN(_18068_));
 AOI22_X1 _24156_ (.A1(\core.keymem.key_mem[4][43] ),
    .A2(_16499_),
    .B1(_17193_),
    .B2(\core.keymem.key_mem[13][43] ),
    .ZN(_18069_));
 NAND4_X1 _24157_ (.A1(_18066_),
    .A2(_18067_),
    .A3(_18068_),
    .A4(_18069_),
    .ZN(_18070_));
 AOI22_X1 _24158_ (.A1(\core.keymem.key_mem[9][43] ),
    .A2(_17522_),
    .B1(_17000_),
    .B2(\core.keymem.key_mem[12][43] ),
    .ZN(_18071_));
 AOI22_X1 _24159_ (.A1(\core.keymem.key_mem[6][43] ),
    .A2(_16520_),
    .B1(_17004_),
    .B2(\core.keymem.key_mem[5][43] ),
    .ZN(_18072_));
 AOI22_X1 _24160_ (.A1(\core.keymem.key_mem[14][43] ),
    .A2(_16998_),
    .B1(_16986_),
    .B2(\core.keymem.key_mem[3][43] ),
    .ZN(_18073_));
 NAND3_X1 _24161_ (.A1(_18071_),
    .A2(_18072_),
    .A3(_18073_),
    .ZN(_18074_));
 NOR2_X1 _24162_ (.A1(_18070_),
    .A2(_18074_),
    .ZN(_18075_));
 MUX2_X2 _24163_ (.A(_00283_),
    .B(_18075_),
    .S(_16488_),
    .Z(_18076_));
 XNOR2_X1 _24164_ (.A(_18065_),
    .B(_18076_),
    .ZN(_18077_));
 BUF_X4 _24165_ (.A(_17709_),
    .Z(_18078_));
 OAI22_X1 _24166_ (.A1(_18052_),
    .A2(_18064_),
    .B1(_18077_),
    .B2(_18078_),
    .ZN(_18079_));
 NOR3_X1 _24167_ (.A1(_16367_),
    .A2(_18051_),
    .A3(_18079_),
    .ZN(_18080_));
 AOI22_X1 _24168_ (.A1(_17746_),
    .A2(_17744_),
    .B1(_17953_),
    .B2(_18080_),
    .ZN(_00569_));
 NAND2_X1 _24169_ (.A1(_17371_),
    .A2(_17255_),
    .ZN(_18081_));
 AOI22_X2 _24170_ (.A1(_17397_),
    .A2(_18018_),
    .B1(_18081_),
    .B2(_18003_),
    .ZN(_18082_));
 AOI21_X1 _24171_ (.A(_17384_),
    .B1(_17484_),
    .B2(_17471_),
    .ZN(_18083_));
 AOI21_X1 _24172_ (.A(_18083_),
    .B1(_17268_),
    .B2(_17272_),
    .ZN(_18084_));
 OAI21_X1 _24173_ (.A(_17482_),
    .B1(_18082_),
    .B2(_18084_),
    .ZN(_18085_));
 NAND2_X1 _24174_ (.A1(_17272_),
    .A2(_17429_),
    .ZN(_18086_));
 OAI221_X2 _24175_ (.A(_17221_),
    .B1(_17272_),
    .B2(_17360_),
    .C1(_17487_),
    .C2(_18086_),
    .ZN(_18087_));
 NAND2_X2 _24176_ (.A1(_17293_),
    .A2(_17404_),
    .ZN(_18088_));
 AOI221_X2 _24177_ (.A(_17458_),
    .B1(_17467_),
    .B2(_18088_),
    .C1(_17279_),
    .C2(_17323_),
    .ZN(_18089_));
 MUX2_X1 _24178_ (.A(_17355_),
    .B(_17455_),
    .S(_17266_),
    .Z(_18090_));
 AOI221_X2 _24179_ (.A(_18089_),
    .B1(_18090_),
    .B2(_17302_),
    .C1(_17494_),
    .C2(_17445_),
    .ZN(_18091_));
 NAND3_X2 _24180_ (.A1(_18085_),
    .A2(_18087_),
    .A3(_18091_),
    .ZN(_18092_));
 NAND2_X1 _24181_ (.A1(_17401_),
    .A2(_17993_),
    .ZN(_18093_));
 OAI22_X1 _24182_ (.A1(_17479_),
    .A2(_17391_),
    .B1(_18093_),
    .B2(_17258_),
    .ZN(_18094_));
 NAND2_X1 _24183_ (.A1(_18003_),
    .A2(_18094_),
    .ZN(_18095_));
 NAND3_X1 _24184_ (.A1(_17271_),
    .A2(_17267_),
    .A3(_17404_),
    .ZN(_18096_));
 AOI21_X1 _24185_ (.A(_17212_),
    .B1(_18011_),
    .B2(_18096_),
    .ZN(_18097_));
 AOI21_X1 _24186_ (.A(_17299_),
    .B1(_17491_),
    .B2(_17294_),
    .ZN(_18098_));
 OAI22_X1 _24187_ (.A1(_17280_),
    .A2(_18018_),
    .B1(_18098_),
    .B2(_17271_),
    .ZN(_18099_));
 NOR3_X1 _24188_ (.A1(_17479_),
    .A2(_18097_),
    .A3(_18099_),
    .ZN(_18100_));
 NAND2_X1 _24189_ (.A1(_17271_),
    .A2(_17368_),
    .ZN(_18101_));
 NAND2_X1 _24190_ (.A1(_17254_),
    .A2(_17265_),
    .ZN(_18102_));
 NAND3_X1 _24191_ (.A1(_17228_),
    .A2(_17486_),
    .A3(_18102_),
    .ZN(_18103_));
 AOI21_X1 _24192_ (.A(_17220_),
    .B1(_18101_),
    .B2(_18103_),
    .ZN(_18104_));
 OAI221_X2 _24193_ (.A(_18095_),
    .B1(_18100_),
    .B2(_18104_),
    .C1(_17317_),
    .C2(_17989_),
    .ZN(_18105_));
 NOR2_X2 _24194_ (.A1(_17264_),
    .A2(_17451_),
    .ZN(_18106_));
 OAI21_X1 _24195_ (.A(_17227_),
    .B1(_17345_),
    .B2(_18106_),
    .ZN(_18107_));
 AOI221_X2 _24196_ (.A(_17357_),
    .B1(_17448_),
    .B2(_18107_),
    .C1(_17270_),
    .C2(_17211_),
    .ZN(_18108_));
 OAI21_X1 _24197_ (.A(_17437_),
    .B1(_17317_),
    .B2(_17434_),
    .ZN(_18109_));
 AOI21_X1 _24198_ (.A(_18108_),
    .B1(_18109_),
    .B2(_17377_),
    .ZN(_18110_));
 INV_X1 _24199_ (.A(_18110_),
    .ZN(_18111_));
 MUX2_X1 _24200_ (.A(_17253_),
    .B(_17322_),
    .S(_17296_),
    .Z(_18112_));
 NOR3_X1 _24201_ (.A1(_17258_),
    .A2(_17338_),
    .A3(_18112_),
    .ZN(_18113_));
 AOI221_X2 _24202_ (.A(_18113_),
    .B1(_17472_),
    .B2(_17496_),
    .C1(_17493_),
    .C2(_17398_),
    .ZN(_18114_));
 AOI22_X2 _24203_ (.A1(_17270_),
    .A2(_17355_),
    .B1(_17471_),
    .B2(_17219_),
    .ZN(_18115_));
 MUX2_X1 _24204_ (.A(_17307_),
    .B(_17390_),
    .S(_17227_),
    .Z(_18116_));
 OAI221_X2 _24205_ (.A(_18114_),
    .B1(_18115_),
    .B2(_17267_),
    .C1(_18116_),
    .C2(_17220_),
    .ZN(_18117_));
 NOR3_X1 _24206_ (.A1(_17269_),
    .A2(_17265_),
    .A3(_17429_),
    .ZN(_18118_));
 OAI21_X1 _24207_ (.A(_17397_),
    .B1(_17353_),
    .B2(_17367_),
    .ZN(_18119_));
 NOR2_X2 _24208_ (.A1(_17219_),
    .A2(_17474_),
    .ZN(_18120_));
 AOI221_X2 _24209_ (.A(_18118_),
    .B1(_18119_),
    .B2(_17313_),
    .C1(_17270_),
    .C2(_18120_),
    .ZN(_18121_));
 AOI22_X2 _24210_ (.A1(_17301_),
    .A2(_17350_),
    .B1(_17359_),
    .B2(_17313_),
    .ZN(_18122_));
 OAI221_X2 _24211_ (.A(_18121_),
    .B1(_17423_),
    .B2(_17308_),
    .C1(_17280_),
    .C2(_18122_),
    .ZN(_18123_));
 AOI21_X1 _24212_ (.A(_17281_),
    .B1(_17392_),
    .B2(_17361_),
    .ZN(_18124_));
 OR3_X1 _24213_ (.A1(_17357_),
    .A2(_17382_),
    .A3(_18124_),
    .ZN(_18125_));
 NOR2_X1 _24214_ (.A1(_17325_),
    .A2(_17410_),
    .ZN(_18126_));
 AOI21_X1 _24215_ (.A(_18126_),
    .B1(_17351_),
    .B2(_17493_),
    .ZN(_18127_));
 OAI21_X1 _24216_ (.A(_17417_),
    .B1(_17467_),
    .B2(_17211_),
    .ZN(_18128_));
 NAND2_X1 _24217_ (.A1(_17343_),
    .A2(_18128_),
    .ZN(_18129_));
 AND4_X1 _24218_ (.A1(_17356_),
    .A2(_18125_),
    .A3(_18127_),
    .A4(_18129_),
    .ZN(_18130_));
 AOI21_X1 _24219_ (.A(_17245_),
    .B1(_17278_),
    .B2(_17226_),
    .ZN(_18131_));
 OAI22_X1 _24220_ (.A1(_17269_),
    .A2(_17288_),
    .B1(_18131_),
    .B2(_17296_),
    .ZN(_18132_));
 AOI21_X1 _24221_ (.A(_17493_),
    .B1(_18132_),
    .B2(_17285_),
    .ZN(_18133_));
 OR2_X1 _24222_ (.A1(_17219_),
    .A2(_18133_),
    .ZN(_18134_));
 OAI21_X1 _24223_ (.A(_17386_),
    .B1(_17368_),
    .B2(_17219_),
    .ZN(_18135_));
 OAI21_X1 _24224_ (.A(_17227_),
    .B1(_17478_),
    .B2(_18135_),
    .ZN(_18136_));
 AND3_X1 _24225_ (.A1(_17986_),
    .A2(_18134_),
    .A3(_18136_),
    .ZN(_18137_));
 NOR4_X4 _24226_ (.A1(_17234_),
    .A2(_17295_),
    .A3(_17287_),
    .A4(_17284_),
    .ZN(_18138_));
 NOR2_X1 _24227_ (.A1(_17355_),
    .A2(_18138_),
    .ZN(_18139_));
 OAI22_X2 _24228_ (.A1(_17955_),
    .A2(_17396_),
    .B1(_17440_),
    .B2(_18139_),
    .ZN(_18140_));
 AOI221_X2 _24229_ (.A(_18140_),
    .B1(_17492_),
    .B2(_17350_),
    .C1(_17304_),
    .C2(_17359_),
    .ZN(_18141_));
 AOI22_X1 _24230_ (.A1(_17269_),
    .A2(_17350_),
    .B1(_17455_),
    .B2(_17483_),
    .ZN(_18142_));
 OAI21_X2 _24231_ (.A(_18141_),
    .B1(_18142_),
    .B2(_17983_),
    .ZN(_18143_));
 MUX2_X1 _24232_ (.A(_17455_),
    .B(_17446_),
    .S(_17210_),
    .Z(_18144_));
 MUX2_X1 _24233_ (.A(_17366_),
    .B(_18144_),
    .S(_17264_),
    .Z(_18145_));
 XNOR2_X1 _24234_ (.A(_17295_),
    .B(_17252_),
    .ZN(_18146_));
 AOI22_X1 _24235_ (.A1(_17284_),
    .A2(_17348_),
    .B1(_18146_),
    .B2(_17278_),
    .ZN(_18147_));
 OAI33_X1 _24236_ (.A1(_17284_),
    .A2(_17265_),
    .A3(_17382_),
    .B1(_18147_),
    .B2(_17357_),
    .B3(_17226_),
    .ZN(_18148_));
 AOI221_X2 _24237_ (.A(_18143_),
    .B1(_18145_),
    .B2(_17380_),
    .C1(_17245_),
    .C2(_18148_),
    .ZN(_18149_));
 NAND4_X1 _24238_ (.A1(_17454_),
    .A2(_18130_),
    .A3(_18137_),
    .A4(_18149_),
    .ZN(_18150_));
 OR4_X1 _24239_ (.A1(_18111_),
    .A2(_18117_),
    .A3(_18123_),
    .A4(_18150_),
    .ZN(_18151_));
 OAI33_X1 _24240_ (.A1(_17463_),
    .A2(_17987_),
    .A3(_17450_),
    .B1(_18092_),
    .B2(_18105_),
    .B3(_18151_),
    .ZN(_18152_));
 AOI21_X1 _24241_ (.A(_18032_),
    .B1(_17418_),
    .B2(_17368_),
    .ZN(_18153_));
 MUX2_X1 _24242_ (.A(_17355_),
    .B(_18138_),
    .S(_17280_),
    .Z(_18154_));
 AOI221_X2 _24243_ (.A(_18153_),
    .B1(_18154_),
    .B2(_17492_),
    .C1(_17996_),
    .C2(_17456_),
    .ZN(_18155_));
 MUX2_X1 _24244_ (.A(_17468_),
    .B(_17486_),
    .S(_17353_),
    .Z(_18156_));
 OAI21_X1 _24245_ (.A(_18155_),
    .B1(_18156_),
    .B2(_17989_),
    .ZN(_18157_));
 NOR2_X2 _24246_ (.A1(net15),
    .A2(_18157_),
    .ZN(_18158_));
 INV_X1 _24247_ (.A(_18123_),
    .ZN(_18159_));
 NAND2_X1 _24248_ (.A1(_17213_),
    .A2(_17255_),
    .ZN(_18160_));
 NAND2_X1 _24249_ (.A1(_17213_),
    .A2(_17471_),
    .ZN(_18161_));
 AOI21_X1 _24250_ (.A(_17464_),
    .B1(_17255_),
    .B2(_17371_),
    .ZN(_18162_));
 AOI221_X2 _24251_ (.A(_17272_),
    .B1(_17464_),
    .B2(_18160_),
    .C1(_18161_),
    .C2(_18162_),
    .ZN(_18163_));
 CLKBUF_X3 _24252_ (.A(_17229_),
    .Z(_18164_));
 NOR3_X1 _24253_ (.A1(_18164_),
    .A2(_17364_),
    .A3(_17317_),
    .ZN(_18165_));
 OAI21_X2 _24254_ (.A(_18017_),
    .B1(_18163_),
    .B2(_18165_),
    .ZN(_18166_));
 AOI21_X1 _24255_ (.A(_17377_),
    .B1(_17968_),
    .B2(_17220_),
    .ZN(_18167_));
 OAI22_X1 _24256_ (.A1(_17316_),
    .A2(_17459_),
    .B1(_18167_),
    .B2(_17319_),
    .ZN(_18168_));
 AND2_X1 _24257_ (.A1(_17494_),
    .A2(_18168_),
    .ZN(_18169_));
 NOR2_X2 _24258_ (.A1(_17323_),
    .A2(_17468_),
    .ZN(_18170_));
 OAI22_X2 _24259_ (.A1(_18005_),
    .A2(_18169_),
    .B1(_18170_),
    .B2(_17494_),
    .ZN(_18171_));
 NAND4_X2 _24260_ (.A1(_17413_),
    .A2(_18159_),
    .A3(_18166_),
    .A4(_18171_),
    .ZN(_18172_));
 NAND3_X1 _24261_ (.A1(_17211_),
    .A2(_17494_),
    .A3(_17398_),
    .ZN(_18173_));
 NAND3_X1 _24262_ (.A1(_17323_),
    .A2(_18005_),
    .A3(_17491_),
    .ZN(_18174_));
 NAND2_X1 _24263_ (.A1(_18173_),
    .A2(_18174_),
    .ZN(_18175_));
 OAI21_X1 _24264_ (.A(_17415_),
    .B1(_17468_),
    .B2(_17266_),
    .ZN(_18176_));
 NAND3_X1 _24265_ (.A1(_17239_),
    .A2(_17302_),
    .A3(_17353_),
    .ZN(_18177_));
 OAI21_X1 _24266_ (.A(_18177_),
    .B1(_17436_),
    .B2(_17239_),
    .ZN(_18178_));
 AOI221_X2 _24267_ (.A(_18175_),
    .B1(_18176_),
    .B2(_17304_),
    .C1(_17389_),
    .C2(_18178_),
    .ZN(_18179_));
 OAI21_X1 _24268_ (.A(_17422_),
    .B1(_17384_),
    .B2(_17255_),
    .ZN(_18180_));
 OAI21_X1 _24269_ (.A(_18180_),
    .B1(_18032_),
    .B2(_17397_),
    .ZN(_18181_));
 OAI21_X1 _24270_ (.A(_17305_),
    .B1(_17484_),
    .B2(_17983_),
    .ZN(_18182_));
 NAND2_X1 _24271_ (.A1(_17308_),
    .A2(_17429_),
    .ZN(_18183_));
 AOI221_X1 _24272_ (.A(_18181_),
    .B1(_18182_),
    .B2(_17255_),
    .C1(_18183_),
    .C2(_17354_),
    .ZN(_18184_));
 OAI33_X1 _24273_ (.A1(_17296_),
    .A2(_17305_),
    .A3(_17344_),
    .B1(_17353_),
    .B2(_17441_),
    .B3(_17338_),
    .ZN(_18185_));
 NOR2_X2 _24274_ (.A1(_17323_),
    .A2(_17458_),
    .ZN(_18186_));
 OAI21_X1 _24275_ (.A(_17468_),
    .B1(_17467_),
    .B2(_17212_),
    .ZN(_18187_));
 AOI221_X2 _24276_ (.A(_18185_),
    .B1(_18186_),
    .B2(_17456_),
    .C1(_17351_),
    .C2(_18187_),
    .ZN(_18188_));
 NAND3_X1 _24277_ (.A1(_18179_),
    .A2(_18184_),
    .A3(_18188_),
    .ZN(_18189_));
 OAI21_X1 _24278_ (.A(_17971_),
    .B1(_17468_),
    .B2(_17314_),
    .ZN(_18190_));
 NOR2_X1 _24279_ (.A1(_17393_),
    .A2(_17307_),
    .ZN(_18191_));
 OAI22_X2 _24280_ (.A1(_17308_),
    .A2(_17436_),
    .B1(_17439_),
    .B2(_17391_),
    .ZN(_18192_));
 AOI221_X2 _24281_ (.A(_18190_),
    .B1(_18191_),
    .B2(_17401_),
    .C1(_18192_),
    .C2(_17371_),
    .ZN(_18193_));
 AOI221_X2 _24282_ (.A(_17211_),
    .B1(_17265_),
    .B2(_17493_),
    .C1(_17306_),
    .C2(_17347_),
    .ZN(_18194_));
 NOR3_X1 _24283_ (.A1(_17213_),
    .A2(_17987_),
    .A3(_18194_),
    .ZN(_18195_));
 NAND3_X1 _24284_ (.A1(_17276_),
    .A2(_17267_),
    .A3(_17347_),
    .ZN(_18196_));
 OAI21_X1 _24285_ (.A(_18196_),
    .B1(_18088_),
    .B2(_17464_),
    .ZN(_18197_));
 AOI21_X1 _24286_ (.A(_18195_),
    .B1(_18197_),
    .B2(_17321_),
    .ZN(_18198_));
 NAND2_X1 _24287_ (.A1(_18193_),
    .A2(_18198_),
    .ZN(_18199_));
 OAI33_X1 _24288_ (.A1(_17228_),
    .A2(_17324_),
    .A3(_17437_),
    .B1(_17989_),
    .B2(_17391_),
    .B3(_17279_),
    .ZN(_18200_));
 AOI21_X1 _24289_ (.A(_18200_),
    .B1(_18138_),
    .B2(_17398_),
    .ZN(_18201_));
 NOR2_X1 _24290_ (.A1(_17212_),
    .A2(_17317_),
    .ZN(_18202_));
 MUX2_X1 _24291_ (.A(_17350_),
    .B(_17384_),
    .S(_17267_),
    .Z(_18203_));
 AOI21_X1 _24292_ (.A(_18202_),
    .B1(_18203_),
    .B2(_17213_),
    .ZN(_18204_));
 OAI21_X1 _24293_ (.A(_18201_),
    .B1(_18204_),
    .B2(_17338_),
    .ZN(_18205_));
 MUX2_X1 _24294_ (.A(_17310_),
    .B(_17448_),
    .S(_17270_),
    .Z(_18206_));
 OAI22_X1 _24295_ (.A1(_17479_),
    .A2(_18038_),
    .B1(_18206_),
    .B2(_17427_),
    .ZN(_18207_));
 NAND2_X1 _24296_ (.A1(_17316_),
    .A2(_18207_),
    .ZN(_18208_));
 NOR2_X1 _24297_ (.A1(_17459_),
    .A2(_17418_),
    .ZN(_18209_));
 NOR2_X1 _24298_ (.A1(_17213_),
    .A2(_17401_),
    .ZN(_18210_));
 AOI21_X1 _24299_ (.A(_18209_),
    .B1(_18210_),
    .B2(_17491_),
    .ZN(_18211_));
 OAI21_X2 _24300_ (.A(_18208_),
    .B1(_18211_),
    .B2(_17268_),
    .ZN(_18212_));
 OR4_X1 _24301_ (.A1(_18189_),
    .A2(_18199_),
    .A3(_18205_),
    .A4(_18212_),
    .ZN(_18213_));
 NAND2_X2 _24302_ (.A1(_17401_),
    .A2(_18138_),
    .ZN(_18214_));
 NAND2_X1 _24303_ (.A1(_17441_),
    .A2(_18214_),
    .ZN(_18215_));
 AOI221_X2 _24304_ (.A(_17272_),
    .B1(_17414_),
    .B2(_17221_),
    .C1(_18215_),
    .C2(_17316_),
    .ZN(_18216_));
 AOI221_X2 _24305_ (.A(_17229_),
    .B1(_17405_),
    .B2(_17414_),
    .C1(_17300_),
    .C2(_17221_),
    .ZN(_18217_));
 NOR3_X2 _24306_ (.A1(_17965_),
    .A2(_18216_),
    .A3(_18217_),
    .ZN(_18218_));
 OAI21_X1 _24307_ (.A(_17464_),
    .B1(_17369_),
    .B2(_17404_),
    .ZN(_18219_));
 AOI21_X1 _24308_ (.A(_17338_),
    .B1(_18088_),
    .B2(_18219_),
    .ZN(_18220_));
 OAI21_X1 _24309_ (.A(_18032_),
    .B1(_18194_),
    .B2(_17987_),
    .ZN(_18221_));
 NOR4_X1 _24310_ (.A1(_17239_),
    .A2(_17288_),
    .A3(_17285_),
    .A4(_17977_),
    .ZN(_18222_));
 OAI21_X1 _24311_ (.A(_17343_),
    .B1(_17346_),
    .B2(_18222_),
    .ZN(_18223_));
 OAI21_X1 _24312_ (.A(_18223_),
    .B1(_17436_),
    .B2(_17467_),
    .ZN(_18224_));
 AOI221_X2 _24313_ (.A(_18220_),
    .B1(_18221_),
    .B2(_17384_),
    .C1(_18224_),
    .C2(_17214_),
    .ZN(_18225_));
 INV_X1 _24314_ (.A(_18225_),
    .ZN(_18226_));
 NOR4_X4 _24315_ (.A1(_18172_),
    .A2(_18213_),
    .A3(_18218_),
    .A4(_18226_),
    .ZN(_18227_));
 AOI21_X4 _24316_ (.A(_17379_),
    .B1(_18158_),
    .B2(_18227_),
    .ZN(_18228_));
 NAND2_X1 _24317_ (.A1(_00288_),
    .A2(_16984_),
    .ZN(_18229_));
 AOI222_X2 _24318_ (.A1(\core.keymem.key_mem[2][44] ),
    .A2(_16994_),
    .B1(_16525_),
    .B2(\core.keymem.key_mem[1][44] ),
    .C1(_17715_),
    .C2(\core.keymem.key_mem[10][44] ),
    .ZN(_18230_));
 AOI22_X2 _24319_ (.A1(\core.keymem.key_mem[8][44] ),
    .A2(_16453_),
    .B1(_17683_),
    .B2(\core.keymem.key_mem[3][44] ),
    .ZN(_18231_));
 BUF_X8 _24320_ (.A(_16947_),
    .Z(_18232_));
 AOI22_X2 _24321_ (.A1(\core.keymem.key_mem[4][44] ),
    .A2(_18232_),
    .B1(_16443_),
    .B2(\core.keymem.key_mem[11][44] ),
    .ZN(_18233_));
 NAND3_X2 _24322_ (.A1(_18230_),
    .A2(_18231_),
    .A3(_18233_),
    .ZN(_18234_));
 AOI21_X1 _24323_ (.A(_16546_),
    .B1(_16537_),
    .B2(\core.keymem.key_mem[9][44] ),
    .ZN(_18235_));
 AOI22_X2 _24324_ (.A1(\core.keymem.key_mem[14][44] ),
    .A2(_16439_),
    .B1(_17789_),
    .B2(\core.keymem.key_mem[7][44] ),
    .ZN(_18236_));
 AOI22_X2 _24325_ (.A1(\core.keymem.key_mem[6][44] ),
    .A2(_16991_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][44] ),
    .ZN(_18237_));
 AOI22_X2 _24326_ (.A1(\core.keymem.key_mem[12][44] ),
    .A2(_17001_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][44] ),
    .ZN(_18238_));
 NAND4_X2 _24327_ (.A1(_18235_),
    .A2(_18236_),
    .A3(_18237_),
    .A4(_18238_),
    .ZN(_18239_));
 OAI21_X4 _24328_ (.A(_18229_),
    .B1(_18234_),
    .B2(_18239_),
    .ZN(_18240_));
 XNOR2_X1 _24329_ (.A(\block_reg[2][12] ),
    .B(_18240_),
    .ZN(_18241_));
 AOI21_X1 _24330_ (.A(_16367_),
    .B1(_16371_),
    .B2(_18241_),
    .ZN(_18242_));
 XNOR2_X2 _24331_ (.A(_17604_),
    .B(_17935_),
    .ZN(_18243_));
 XNOR2_X1 _24332_ (.A(_17866_),
    .B(_18243_),
    .ZN(_18244_));
 XNOR2_X2 _24333_ (.A(_17592_),
    .B(_18244_),
    .ZN(_18245_));
 XNOR2_X1 _24334_ (.A(_17689_),
    .B(_17946_),
    .ZN(_18246_));
 XNOR2_X2 _24335_ (.A(_17797_),
    .B(_18246_),
    .ZN(_18247_));
 AOI222_X2 _24336_ (.A1(\core.keymem.key_mem[14][49] ),
    .A2(_16999_),
    .B1(_17715_),
    .B2(\core.keymem.key_mem[10][49] ),
    .C1(_16949_),
    .C2(\core.keymem.key_mem[5][49] ),
    .ZN(_18248_));
 AOI22_X1 _24337_ (.A1(\core.keymem.key_mem[4][49] ),
    .A2(_16500_),
    .B1(_17781_),
    .B2(\core.keymem.key_mem[8][49] ),
    .ZN(_18249_));
 AOI22_X1 _24338_ (.A1(\core.keymem.key_mem[2][49] ),
    .A2(_16994_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][49] ),
    .ZN(_18250_));
 NAND3_X1 _24339_ (.A1(_18248_),
    .A2(_18249_),
    .A3(_18250_),
    .ZN(_18251_));
 AOI22_X1 _24340_ (.A1(\core.keymem.key_mem[6][49] ),
    .A2(_16521_),
    .B1(_17008_),
    .B2(\core.keymem.key_mem[11][49] ),
    .ZN(_18252_));
 AOI22_X1 _24341_ (.A1(\core.keymem.key_mem[12][49] ),
    .A2(_17001_),
    .B1(_16525_),
    .B2(\core.keymem.key_mem[1][49] ),
    .ZN(_18253_));
 AOI22_X1 _24342_ (.A1(\core.keymem.key_mem[3][49] ),
    .A2(_16987_),
    .B1(_17668_),
    .B2(\core.keymem.key_mem[9][49] ),
    .ZN(_18254_));
 AOI21_X1 _24343_ (.A(_16495_),
    .B1(_17789_),
    .B2(\core.keymem.key_mem[7][49] ),
    .ZN(_18255_));
 NAND4_X1 _24344_ (.A1(_18252_),
    .A2(_18253_),
    .A3(_18254_),
    .A4(_18255_),
    .ZN(_18256_));
 NOR2_X2 _24345_ (.A1(_18251_),
    .A2(_18256_),
    .ZN(_18257_));
 AOI21_X4 _24346_ (.A(_18257_),
    .B1(_16873_),
    .B2(_00274_),
    .ZN(_18258_));
 XNOR2_X2 _24347_ (.A(\core.dec_block.block_w2_reg[17] ),
    .B(_18258_),
    .ZN(_18259_));
 XNOR2_X2 _24348_ (.A(_17574_),
    .B(_18259_),
    .ZN(_18260_));
 XNOR2_X2 _24349_ (.A(_17824_),
    .B(_17891_),
    .ZN(_18261_));
 XNOR2_X2 _24350_ (.A(_18260_),
    .B(_18261_),
    .ZN(_18262_));
 XNOR2_X2 _24351_ (.A(_18247_),
    .B(_18262_),
    .ZN(_18263_));
 XNOR2_X2 _24352_ (.A(_18245_),
    .B(_18263_),
    .ZN(_18264_));
 XNOR2_X2 _24353_ (.A(_17673_),
    .B(_17761_),
    .ZN(_18265_));
 INV_X1 _24354_ (.A(\core.dec_block.block_w2_reg[11] ),
    .ZN(_18266_));
 XNOR2_X2 _24355_ (.A(_18266_),
    .B(_18076_),
    .ZN(_18267_));
 XNOR2_X2 _24356_ (.A(_17848_),
    .B(_18267_),
    .ZN(_18268_));
 XOR2_X2 _24357_ (.A(_18265_),
    .B(_18268_),
    .Z(_18269_));
 INV_X1 _24358_ (.A(\core.dec_block.block_w2_reg[4] ),
    .ZN(_18270_));
 NAND2_X1 _24359_ (.A1(_00289_),
    .A2(_16498_),
    .ZN(_18271_));
 AOI22_X1 _24360_ (.A1(\core.keymem.key_mem[2][36] ),
    .A2(_16425_),
    .B1(_16417_),
    .B2(\core.keymem.key_mem[1][36] ),
    .ZN(_18272_));
 AOI22_X1 _24361_ (.A1(\core.keymem.key_mem[7][36] ),
    .A2(_16408_),
    .B1(_16991_),
    .B2(\core.keymem.key_mem[6][36] ),
    .ZN(_18273_));
 AOI22_X1 _24362_ (.A1(\core.keymem.key_mem[9][36] ),
    .A2(_16463_),
    .B1(_17768_),
    .B2(\core.keymem.key_mem[11][36] ),
    .ZN(_18274_));
 AOI22_X1 _24363_ (.A1(\core.keymem.key_mem[4][36] ),
    .A2(_18232_),
    .B1(_17683_),
    .B2(\core.keymem.key_mem[3][36] ),
    .ZN(_18275_));
 AND4_X1 _24364_ (.A1(_18272_),
    .A2(_18273_),
    .A3(_18274_),
    .A4(_18275_),
    .ZN(_18276_));
 AOI22_X2 _24365_ (.A1(\core.keymem.key_mem[12][36] ),
    .A2(_17093_),
    .B1(_16510_),
    .B2(\core.keymem.key_mem[5][36] ),
    .ZN(_18277_));
 AOI22_X2 _24366_ (.A1(\core.keymem.key_mem[14][36] ),
    .A2(_17581_),
    .B1(_17082_),
    .B2(\core.keymem.key_mem[10][36] ),
    .ZN(_18278_));
 AOI22_X2 _24367_ (.A1(\core.keymem.key_mem[8][36] ),
    .A2(_17765_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][36] ),
    .ZN(_18279_));
 NAND4_X2 _24368_ (.A1(_18276_),
    .A2(_18277_),
    .A3(_18278_),
    .A4(_18279_),
    .ZN(_18280_));
 OAI21_X4 _24369_ (.A(_18271_),
    .B1(_18280_),
    .B2(_17578_),
    .ZN(_18281_));
 XNOR2_X2 _24370_ (.A(_18270_),
    .B(_18281_),
    .ZN(_18282_));
 XNOR2_X2 _24371_ (.A(_17518_),
    .B(_17862_),
    .ZN(_18283_));
 XNOR2_X2 _24372_ (.A(_18282_),
    .B(_18283_),
    .ZN(_18284_));
 INV_X1 _24373_ (.A(\core.dec_block.block_w2_reg[20] ),
    .ZN(_18285_));
 NAND2_X1 _24374_ (.A1(_00290_),
    .A2(_17578_),
    .ZN(_18286_));
 AOI22_X1 _24375_ (.A1(\core.keymem.key_mem[5][52] ),
    .A2(_16510_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][52] ),
    .ZN(_18287_));
 AOI22_X1 _24376_ (.A1(\core.keymem.key_mem[4][52] ),
    .A2(_16458_),
    .B1(_16449_),
    .B2(\core.keymem.key_mem[6][52] ),
    .ZN(_18288_));
 AOI22_X1 _24377_ (.A1(\core.keymem.key_mem[3][52] ),
    .A2(_16387_),
    .B1(_17178_),
    .B2(\core.keymem.key_mem[1][52] ),
    .ZN(_18289_));
 AOI22_X1 _24378_ (.A1(\core.keymem.key_mem[14][52] ),
    .A2(_16502_),
    .B1(_16408_),
    .B2(\core.keymem.key_mem[7][52] ),
    .ZN(_18290_));
 AND4_X1 _24379_ (.A1(_18287_),
    .A2(_18288_),
    .A3(_18289_),
    .A4(_18290_),
    .ZN(_18291_));
 AOI22_X2 _24380_ (.A1(\core.keymem.key_mem[10][52] ),
    .A2(_17082_),
    .B1(_17769_),
    .B2(\core.keymem.key_mem[11][52] ),
    .ZN(_18292_));
 AOI22_X2 _24381_ (.A1(\core.keymem.key_mem[2][52] ),
    .A2(_17086_),
    .B1(_17585_),
    .B2(\core.keymem.key_mem[9][52] ),
    .ZN(_18293_));
 AOI22_X2 _24382_ (.A1(\core.keymem.key_mem[8][52] ),
    .A2(_17765_),
    .B1(_17093_),
    .B2(\core.keymem.key_mem[12][52] ),
    .ZN(_18294_));
 NAND4_X2 _24383_ (.A1(_18291_),
    .A2(_18292_),
    .A3(_18293_),
    .A4(_18294_),
    .ZN(_18295_));
 OAI21_X4 _24384_ (.A(_18286_),
    .B1(_18295_),
    .B2(_16549_),
    .ZN(_18296_));
 XNOR2_X2 _24385_ (.A(_18285_),
    .B(_18296_),
    .ZN(_18297_));
 AOI22_X1 _24386_ (.A1(\core.keymem.key_mem[9][60] ),
    .A2(_16463_),
    .B1(_16417_),
    .B2(\core.keymem.key_mem[1][60] ),
    .ZN(_18298_));
 AOI22_X1 _24387_ (.A1(\core.keymem.key_mem[14][60] ),
    .A2(_16439_),
    .B1(_17768_),
    .B2(\core.keymem.key_mem[11][60] ),
    .ZN(_18299_));
 AOI22_X1 _24388_ (.A1(\core.keymem.key_mem[6][60] ),
    .A2(_16991_),
    .B1(_17786_),
    .B2(\core.keymem.key_mem[2][60] ),
    .ZN(_18300_));
 AOI22_X1 _24389_ (.A1(\core.keymem.key_mem[4][60] ),
    .A2(_16500_),
    .B1(_17789_),
    .B2(\core.keymem.key_mem[7][60] ),
    .ZN(_18301_));
 NAND4_X1 _24390_ (.A1(_18298_),
    .A2(_18299_),
    .A3(_18300_),
    .A4(_18301_),
    .ZN(_18302_));
 AOI22_X1 _24391_ (.A1(\core.keymem.key_mem[3][60] ),
    .A2(_17683_),
    .B1(_16433_),
    .B2(\core.keymem.key_mem[10][60] ),
    .ZN(_18303_));
 AOI22_X1 _24392_ (.A1(\core.keymem.key_mem[8][60] ),
    .A2(_16453_),
    .B1(_17001_),
    .B2(\core.keymem.key_mem[12][60] ),
    .ZN(_18304_));
 AOI22_X1 _24393_ (.A1(\core.keymem.key_mem[5][60] ),
    .A2(_17675_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][60] ),
    .ZN(_18305_));
 NAND3_X1 _24394_ (.A1(_18303_),
    .A2(_18304_),
    .A3(_18305_),
    .ZN(_18306_));
 OR3_X1 _24395_ (.A1(_16497_),
    .A2(_18302_),
    .A3(_18306_),
    .ZN(_18307_));
 NAND2_X1 _24396_ (.A1(_00287_),
    .A2(_16548_),
    .ZN(_18308_));
 AND2_X4 _24397_ (.A1(_18307_),
    .A2(_18308_),
    .ZN(_18309_));
 XNOR2_X2 _24398_ (.A(\core.dec_block.block_w2_reg[28] ),
    .B(_18309_),
    .ZN(_18310_));
 XNOR2_X2 _24399_ (.A(_18297_),
    .B(_18310_),
    .ZN(_18311_));
 XOR2_X1 _24400_ (.A(_18284_),
    .B(_18311_),
    .Z(_18312_));
 XNOR2_X1 _24401_ (.A(_18269_),
    .B(_18312_),
    .ZN(_18313_));
 XNOR2_X1 _24402_ (.A(_18264_),
    .B(_18313_),
    .ZN(_18314_));
 AOI22_X1 _24403_ (.A1(\core.keymem.key_mem[12][108] ),
    .A2(_17001_),
    .B1(_16509_),
    .B2(\core.keymem.key_mem[5][108] ),
    .ZN(_18315_));
 AOI22_X1 _24404_ (.A1(\core.keymem.key_mem[14][108] ),
    .A2(_16999_),
    .B1(_17084_),
    .B2(\core.keymem.key_mem[7][108] ),
    .ZN(_18316_));
 AOI22_X1 _24405_ (.A1(\core.keymem.key_mem[8][108] ),
    .A2(_17666_),
    .B1(_17008_),
    .B2(\core.keymem.key_mem[11][108] ),
    .ZN(_18317_));
 AOI22_X1 _24406_ (.A1(\core.keymem.key_mem[2][108] ),
    .A2(_17786_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][108] ),
    .ZN(_18318_));
 NAND4_X1 _24407_ (.A1(_18315_),
    .A2(_18316_),
    .A3(_18317_),
    .A4(_18318_),
    .ZN(_18319_));
 AOI22_X1 _24408_ (.A1(\core.keymem.key_mem[10][108] ),
    .A2(_16989_),
    .B1(_17003_),
    .B2(\core.keymem.key_mem[1][108] ),
    .ZN(_18320_));
 AOI22_X1 _24409_ (.A1(\core.keymem.key_mem[6][108] ),
    .A2(_16521_),
    .B1(_17668_),
    .B2(\core.keymem.key_mem[9][108] ),
    .ZN(_18321_));
 AOI22_X1 _24410_ (.A1(\core.keymem.key_mem[4][108] ),
    .A2(_16500_),
    .B1(_16866_),
    .B2(\core.keymem.key_mem[3][108] ),
    .ZN(_18322_));
 NAND3_X1 _24411_ (.A1(_18320_),
    .A2(_18321_),
    .A3(_18322_),
    .ZN(_18323_));
 NOR3_X2 _24412_ (.A1(_16984_),
    .A2(_18319_),
    .A3(_18323_),
    .ZN(_18324_));
 AOI21_X4 _24413_ (.A(_18324_),
    .B1(_16548_),
    .B2(_00209_),
    .ZN(_18325_));
 XNOR2_X2 _24414_ (.A(\core.dec_block.block_w0_reg[12] ),
    .B(_18325_),
    .ZN(_18326_));
 OAI221_X1 _24415_ (.A(_18242_),
    .B1(_18314_),
    .B2(_17203_),
    .C1(_16556_),
    .C2(_18326_),
    .ZN(_18327_));
 OAI22_X1 _24416_ (.A1(\core.dec_block.block_w0_reg[12] ),
    .A2(_16366_),
    .B1(_18228_),
    .B2(_18327_),
    .ZN(_18328_));
 INV_X1 _24417_ (.A(_18328_),
    .ZN(_00570_));
 BUF_X4 _24418_ (.A(_16364_),
    .Z(_18329_));
 BUF_X4 _24419_ (.A(_18329_),
    .Z(_18330_));
 NOR2_X1 _24420_ (.A1(\core.dec_block.block_w0_reg[13] ),
    .A2(_18330_),
    .ZN(_18331_));
 BUF_X4 _24421_ (.A(_17748_),
    .Z(_18332_));
 BUF_X4 _24422_ (.A(_18332_),
    .Z(_18333_));
 XNOR2_X2 _24423_ (.A(_17577_),
    .B(_17658_),
    .ZN(_18334_));
 XOR2_X2 _24424_ (.A(_17702_),
    .B(_18334_),
    .Z(_18335_));
 XNOR2_X2 _24425_ (.A(_18245_),
    .B(_18335_),
    .ZN(_18336_));
 XOR2_X2 _24426_ (.A(\core.dec_block.block_w2_reg[12] ),
    .B(_18240_),
    .Z(_18337_));
 XNOR2_X2 _24427_ (.A(_17935_),
    .B(_18337_),
    .ZN(_18338_));
 XNOR2_X1 _24428_ (.A(_17891_),
    .B(_18282_),
    .ZN(_18339_));
 XNOR2_X2 _24429_ (.A(_18338_),
    .B(_18339_),
    .ZN(_18340_));
 XNOR2_X2 _24430_ (.A(_17922_),
    .B(_18268_),
    .ZN(_18341_));
 XOR2_X1 _24431_ (.A(_18340_),
    .B(_18341_),
    .Z(_18342_));
 XNOR2_X1 _24432_ (.A(_17761_),
    .B(_17946_),
    .ZN(_18343_));
 XNOR2_X1 _24433_ (.A(_18342_),
    .B(_18343_),
    .ZN(_18344_));
 XNOR2_X1 _24434_ (.A(_18336_),
    .B(_18344_),
    .ZN(_18345_));
 NAND2_X1 _24435_ (.A1(_18333_),
    .A2(_18345_),
    .ZN(_18346_));
 AOI21_X1 _24436_ (.A(_18035_),
    .B1(_18106_),
    .B2(_17271_),
    .ZN(_18347_));
 OR3_X1 _24437_ (.A1(_17479_),
    .A2(_17434_),
    .A3(_18347_),
    .ZN(_18348_));
 AOI222_X2 _24438_ (.A1(_17381_),
    .A2(_17366_),
    .B1(_17496_),
    .B2(_17321_),
    .C1(_17405_),
    .C2(_17255_),
    .ZN(_18349_));
 NAND2_X1 _24439_ (.A1(_17393_),
    .A2(_17377_),
    .ZN(_18350_));
 OAI221_X2 _24440_ (.A(_18348_),
    .B1(_18349_),
    .B2(_17965_),
    .C1(_17463_),
    .C2(_18350_),
    .ZN(_18351_));
 MUX2_X1 _24441_ (.A(_17306_),
    .B(_17348_),
    .S(_17220_),
    .Z(_18352_));
 AOI22_X1 _24442_ (.A1(_17482_),
    .A2(_17471_),
    .B1(_18352_),
    .B2(_17385_),
    .ZN(_18353_));
 OAI22_X1 _24443_ (.A1(_17989_),
    .A2(_17461_),
    .B1(_18353_),
    .B2(_18164_),
    .ZN(_18354_));
 AOI21_X1 _24444_ (.A(_17456_),
    .B1(_17300_),
    .B2(_18164_),
    .ZN(_18355_));
 OAI22_X1 _24445_ (.A1(_17459_),
    .A2(_17368_),
    .B1(_18355_),
    .B2(_18017_),
    .ZN(_18356_));
 AOI221_X2 _24446_ (.A(_18351_),
    .B1(_18354_),
    .B2(_17294_),
    .C1(_18356_),
    .C2(_17325_),
    .ZN(_18357_));
 OAI22_X1 _24447_ (.A1(_17450_),
    .A2(_18214_),
    .B1(_17980_),
    .B2(_18102_),
    .ZN(_18358_));
 NAND2_X1 _24448_ (.A1(_18164_),
    .A2(_18358_),
    .ZN(_18359_));
 NOR2_X1 _24449_ (.A1(_17468_),
    .A2(_17450_),
    .ZN(_18360_));
 NOR3_X1 _24450_ (.A1(_17372_),
    .A2(_17319_),
    .A3(_17441_),
    .ZN(_18361_));
 OAI21_X1 _24451_ (.A(_17302_),
    .B1(_18360_),
    .B2(_18361_),
    .ZN(_18362_));
 OAI21_X1 _24452_ (.A(_17443_),
    .B1(_17496_),
    .B2(_17346_),
    .ZN(_18363_));
 NOR2_X1 _24453_ (.A1(_17213_),
    .A2(_17989_),
    .ZN(_18364_));
 AOI21_X1 _24454_ (.A(_18364_),
    .B1(_17450_),
    .B2(_17381_),
    .ZN(_18365_));
 NAND2_X1 _24455_ (.A1(_17302_),
    .A2(_17491_),
    .ZN(_18366_));
 OAI221_X1 _24456_ (.A(_18363_),
    .B1(_18365_),
    .B2(_17308_),
    .C1(_18366_),
    .C2(_17374_),
    .ZN(_18367_));
 OAI22_X1 _24457_ (.A1(_17256_),
    .A2(_17965_),
    .B1(_17437_),
    .B2(_18164_),
    .ZN(_18368_));
 AOI21_X1 _24458_ (.A(_18367_),
    .B1(_18368_),
    .B2(_18210_),
    .ZN(_18369_));
 AOI21_X1 _24459_ (.A(_17381_),
    .B1(_17377_),
    .B2(_17276_),
    .ZN(_18370_));
 OAI22_X1 _24460_ (.A1(_17276_),
    .A2(_17314_),
    .B1(_17353_),
    .B2(_18370_),
    .ZN(_18371_));
 NAND2_X1 _24461_ (.A1(_17993_),
    .A2(_18371_),
    .ZN(_18372_));
 AOI221_X1 _24462_ (.A(_18170_),
    .B1(_17348_),
    .B2(_17385_),
    .C1(_17371_),
    .C2(_17414_),
    .ZN(_18373_));
 OAI21_X1 _24463_ (.A(_18372_),
    .B1(_18373_),
    .B2(_17440_),
    .ZN(_18374_));
 MUX2_X1 _24464_ (.A(_17393_),
    .B(_17324_),
    .S(_17296_),
    .Z(_18375_));
 NOR2_X1 _24465_ (.A1(_17422_),
    .A2(_17445_),
    .ZN(_18376_));
 OAI33_X1 _24466_ (.A1(_17459_),
    .A2(_17298_),
    .A3(_18375_),
    .B1(_18376_),
    .B2(_17322_),
    .B3(_17382_),
    .ZN(_18377_));
 NAND3_X1 _24467_ (.A1(_17273_),
    .A2(_17384_),
    .A3(_17402_),
    .ZN(_18378_));
 AOI22_X1 _24468_ (.A1(_17494_),
    .A2(_17405_),
    .B1(_18364_),
    .B2(_17346_),
    .ZN(_18379_));
 AOI21_X1 _24469_ (.A(_17965_),
    .B1(_18378_),
    .B2(_18379_),
    .ZN(_18380_));
 NOR3_X1 _24470_ (.A1(_18374_),
    .A2(_18377_),
    .A3(_18380_),
    .ZN(_18381_));
 NAND4_X1 _24471_ (.A1(_18359_),
    .A2(_18362_),
    .A3(_18369_),
    .A4(_18381_),
    .ZN(_18382_));
 NOR3_X2 _24472_ (.A1(_18117_),
    .A2(_18212_),
    .A3(_18382_),
    .ZN(_18383_));
 AOI21_X1 _24473_ (.A(_17404_),
    .B1(_17346_),
    .B2(_17319_),
    .ZN(_18384_));
 OAI21_X1 _24474_ (.A(_17214_),
    .B1(_18164_),
    .B2(_18384_),
    .ZN(_18385_));
 OAI221_X1 _24475_ (.A(_17374_),
    .B1(_17273_),
    .B2(_17486_),
    .C1(_17429_),
    .C2(_17364_),
    .ZN(_18386_));
 NAND3_X1 _24476_ (.A1(_18017_),
    .A2(_18385_),
    .A3(_18386_),
    .ZN(_18387_));
 OAI21_X1 _24477_ (.A(_18387_),
    .B1(_18010_),
    .B2(_18017_),
    .ZN(_18388_));
 AOI21_X1 _24478_ (.A(_17338_),
    .B1(_17467_),
    .B2(_17391_),
    .ZN(_18389_));
 OAI21_X1 _24479_ (.A(_17325_),
    .B1(_18209_),
    .B2(_18389_),
    .ZN(_18390_));
 OAI21_X2 _24480_ (.A(_17408_),
    .B1(_17397_),
    .B2(_17987_),
    .ZN(_18391_));
 AOI22_X4 _24481_ (.A1(_17487_),
    .A2(_17492_),
    .B1(_18391_),
    .B2(_17372_),
    .ZN(_18392_));
 NAND2_X1 _24482_ (.A1(_17267_),
    .A2(_17350_),
    .ZN(_18393_));
 AOI21_X1 _24483_ (.A(_17989_),
    .B1(_17318_),
    .B2(_18393_),
    .ZN(_18394_));
 AOI221_X2 _24484_ (.A(_18394_),
    .B1(_18014_),
    .B2(_17491_),
    .C1(_17350_),
    .C2(_17472_),
    .ZN(_18395_));
 NAND4_X2 _24485_ (.A1(_17444_),
    .A2(_18390_),
    .A3(_18392_),
    .A4(_18395_),
    .ZN(_18396_));
 NOR3_X2 _24486_ (.A1(_18033_),
    .A2(_18388_),
    .A3(_18396_),
    .ZN(_18397_));
 NAND3_X4 _24487_ (.A1(_18357_),
    .A2(_18383_),
    .A3(_18397_),
    .ZN(_18398_));
 BUF_X4 _24488_ (.A(_16555_),
    .Z(_18399_));
 AOI222_X2 _24489_ (.A1(\core.keymem.key_mem[14][109] ),
    .A2(_16437_),
    .B1(_16858_),
    .B2(\core.keymem.key_mem[2][109] ),
    .C1(_16504_),
    .C2(\core.keymem.key_mem[11][109] ),
    .ZN(_18400_));
 AOI22_X1 _24490_ (.A1(\core.keymem.key_mem[6][109] ),
    .A2(_16447_),
    .B1(_16397_),
    .B2(\core.keymem.key_mem[12][109] ),
    .ZN(_18401_));
 AOI22_X1 _24491_ (.A1(\core.keymem.key_mem[1][109] ),
    .A2(_16415_),
    .B1(_16531_),
    .B2(\core.keymem.key_mem[13][109] ),
    .ZN(_18402_));
 AND3_X1 _24492_ (.A1(_18400_),
    .A2(_18401_),
    .A3(_18402_),
    .ZN(_18403_));
 AOI22_X1 _24493_ (.A1(\core.keymem.key_mem[3][109] ),
    .A2(_16385_),
    .B1(_16431_),
    .B2(\core.keymem.key_mem[10][109] ),
    .ZN(_18404_));
 AOI22_X1 _24494_ (.A1(\core.keymem.key_mem[8][109] ),
    .A2(_16451_),
    .B1(_16948_),
    .B2(\core.keymem.key_mem[5][109] ),
    .ZN(_18405_));
 AOI22_X1 _24495_ (.A1(\core.keymem.key_mem[7][109] ),
    .A2(_16406_),
    .B1(_16461_),
    .B2(\core.keymem.key_mem[9][109] ),
    .ZN(_18406_));
 AOI21_X1 _24496_ (.A(_16544_),
    .B1(_16946_),
    .B2(\core.keymem.key_mem[4][109] ),
    .ZN(_18407_));
 AND4_X1 _24497_ (.A1(_18404_),
    .A2(_18405_),
    .A3(_18406_),
    .A4(_18407_),
    .ZN(_18408_));
 AOI22_X4 _24498_ (.A1(_00181_),
    .A2(_16546_),
    .B1(_18403_),
    .B2(_18408_),
    .ZN(_18409_));
 XNOR2_X2 _24499_ (.A(\core.dec_block.block_w0_reg[13] ),
    .B(_18409_),
    .ZN(_18410_));
 XNOR2_X1 _24500_ (.A(\block_reg[2][13] ),
    .B(_17823_),
    .ZN(_18411_));
 BUF_X4 _24501_ (.A(_17709_),
    .Z(_18412_));
 OAI22_X1 _24502_ (.A1(_18399_),
    .A2(_18410_),
    .B1(_18411_),
    .B2(_18412_),
    .ZN(_18413_));
 NOR3_X1 _24503_ (.A1(_17744_),
    .A2(_18398_),
    .A3(_18413_),
    .ZN(_18414_));
 AOI21_X1 _24504_ (.A(_18331_),
    .B1(_18346_),
    .B2(_18414_),
    .ZN(_00571_));
 NOR2_X1 _24505_ (.A1(_17246_),
    .A2(_18330_),
    .ZN(_18415_));
 BUF_X8 _24506_ (.A(_17329_),
    .Z(_18416_));
 INV_X1 _24507_ (.A(_18166_),
    .ZN(_18417_));
 NOR3_X1 _24508_ (.A1(_17272_),
    .A2(_17393_),
    .A3(_17467_),
    .ZN(_18418_));
 MUX2_X1 _24509_ (.A(_17437_),
    .B(_18102_),
    .S(_17227_),
    .Z(_18419_));
 OAI222_X2 _24510_ (.A1(_17368_),
    .A2(_17439_),
    .B1(_18038_),
    .B2(_17427_),
    .C1(_18419_),
    .C2(_17401_),
    .ZN(_18420_));
 AOI221_X2 _24511_ (.A(_17266_),
    .B1(_18138_),
    .B2(_17483_),
    .C1(_17485_),
    .C2(_17494_),
    .ZN(_18421_));
 AOI22_X1 _24512_ (.A1(_17271_),
    .A2(_17300_),
    .B1(_17471_),
    .B2(_17968_),
    .ZN(_18422_));
 AOI21_X1 _24513_ (.A(_18421_),
    .B1(_18422_),
    .B2(_17464_),
    .ZN(_18423_));
 AOI221_X2 _24514_ (.A(_18418_),
    .B1(_18420_),
    .B2(_17372_),
    .C1(_17221_),
    .C2(_18423_),
    .ZN(_18424_));
 OAI21_X1 _24515_ (.A(_17364_),
    .B1(_17391_),
    .B2(_18164_),
    .ZN(_18425_));
 OAI21_X1 _24516_ (.A(_18044_),
    .B1(_17418_),
    .B2(_17229_),
    .ZN(_18426_));
 OAI21_X1 _24517_ (.A(_18425_),
    .B1(_18426_),
    .B2(_17364_),
    .ZN(_18427_));
 NAND2_X1 _24518_ (.A1(_17374_),
    .A2(_17221_),
    .ZN(_18428_));
 NAND3_X1 _24519_ (.A1(_17316_),
    .A2(_17268_),
    .A3(_17456_),
    .ZN(_18429_));
 OAI21_X1 _24520_ (.A(_18429_),
    .B1(_17310_),
    .B2(_17965_),
    .ZN(_18430_));
 AOI22_X1 _24521_ (.A1(_18138_),
    .A2(_17968_),
    .B1(_18430_),
    .B2(_17273_),
    .ZN(_18431_));
 OAI221_X1 _24522_ (.A(_18424_),
    .B1(_18427_),
    .B2(_18428_),
    .C1(_18431_),
    .C2(_17221_),
    .ZN(_18432_));
 OAI21_X1 _24523_ (.A(_18088_),
    .B1(_17353_),
    .B2(_17317_),
    .ZN(_18433_));
 NAND4_X1 _24524_ (.A1(_17258_),
    .A2(_17296_),
    .A3(_17281_),
    .A4(_17267_),
    .ZN(_18434_));
 AOI22_X1 _24525_ (.A1(_17281_),
    .A2(_17306_),
    .B1(_17348_),
    .B2(_17325_),
    .ZN(_18435_));
 OAI21_X1 _24526_ (.A(_18434_),
    .B1(_18435_),
    .B2(_17245_),
    .ZN(_18436_));
 AOI22_X1 _24527_ (.A1(_17302_),
    .A2(_18433_),
    .B1(_18436_),
    .B2(_17321_),
    .ZN(_18437_));
 OAI22_X1 _24528_ (.A1(_17989_),
    .A2(_17391_),
    .B1(_17397_),
    .B2(_17987_),
    .ZN(_18438_));
 AOI21_X1 _24529_ (.A(_18377_),
    .B1(_18438_),
    .B2(_17433_),
    .ZN(_18439_));
 NAND2_X1 _24530_ (.A1(_17975_),
    .A2(_17494_),
    .ZN(_18440_));
 OAI21_X1 _24531_ (.A(_17355_),
    .B1(_17421_),
    .B2(_17996_),
    .ZN(_18441_));
 NAND2_X1 _24532_ (.A1(_18440_),
    .A2(_18441_),
    .ZN(_18442_));
 OAI21_X1 _24533_ (.A(_17496_),
    .B1(_17968_),
    .B2(_18006_),
    .ZN(_18443_));
 OAI21_X1 _24534_ (.A(_18443_),
    .B1(_17310_),
    .B2(_17271_),
    .ZN(_18444_));
 AOI221_X2 _24535_ (.A(_18442_),
    .B1(_18014_),
    .B2(_17346_),
    .C1(_17479_),
    .C2(_18444_),
    .ZN(_18445_));
 NAND4_X1 _24536_ (.A1(_18015_),
    .A2(_18437_),
    .A3(_18439_),
    .A4(_18445_),
    .ZN(_18446_));
 MUX2_X1 _24537_ (.A(_17359_),
    .B(_17404_),
    .S(_17228_),
    .Z(_18447_));
 AOI22_X1 _24538_ (.A1(_17321_),
    .A2(_18202_),
    .B1(_18447_),
    .B2(_17482_),
    .ZN(_18448_));
 NOR2_X1 _24539_ (.A1(_17965_),
    .A2(_18448_),
    .ZN(_18449_));
 OAI22_X1 _24540_ (.A1(_17316_),
    .A2(_17308_),
    .B1(_18139_),
    .B2(_17319_),
    .ZN(_18450_));
 NAND2_X1 _24541_ (.A1(_17377_),
    .A2(_18450_),
    .ZN(_18451_));
 NOR2_X1 _24542_ (.A1(_17463_),
    .A2(_17265_),
    .ZN(_18452_));
 AOI22_X2 _24543_ (.A1(_17266_),
    .A2(_17346_),
    .B1(_18452_),
    .B2(_17227_),
    .ZN(_18453_));
 NOR3_X2 _24544_ (.A1(_17323_),
    .A2(_17357_),
    .A3(_18453_),
    .ZN(_18454_));
 NOR2_X1 _24545_ (.A1(_17401_),
    .A2(_17474_),
    .ZN(_18455_));
 AOI221_X2 _24546_ (.A(_18454_),
    .B1(_18455_),
    .B2(_18037_),
    .C1(_17387_),
    .C2(_17472_),
    .ZN(_18456_));
 NAND2_X1 _24547_ (.A1(_18451_),
    .A2(_18456_),
    .ZN(_18457_));
 NOR3_X1 _24548_ (.A1(_18446_),
    .A2(_18449_),
    .A3(_18457_),
    .ZN(_18458_));
 OAI22_X1 _24549_ (.A1(_17308_),
    .A2(_17955_),
    .B1(_17441_),
    .B2(_17459_),
    .ZN(_18459_));
 AOI21_X1 _24550_ (.A(_18170_),
    .B1(_18035_),
    .B2(_17371_),
    .ZN(_18460_));
 OAI22_X2 _24551_ (.A1(_17459_),
    .A2(_17441_),
    .B1(_18460_),
    .B2(_17479_),
    .ZN(_18461_));
 AOI222_X2 _24552_ (.A1(_17214_),
    .A2(_18459_),
    .B1(_18461_),
    .B2(_17319_),
    .C1(_17360_),
    .C2(_18005_),
    .ZN(_18462_));
 NAND3_X1 _24553_ (.A1(_17420_),
    .A2(_18458_),
    .A3(_18462_),
    .ZN(_18463_));
 OR4_X2 _24554_ (.A1(_18092_),
    .A2(_18417_),
    .A3(_18432_),
    .A4(_18463_),
    .ZN(_18464_));
 OAI21_X2 _24555_ (.A(_18416_),
    .B1(_18152_),
    .B2(_18464_),
    .ZN(_18465_));
 BUF_X4 _24556_ (.A(_17709_),
    .Z(_18466_));
 XNOR2_X1 _24557_ (.A(\block_reg[2][14] ),
    .B(_17701_),
    .ZN(_18467_));
 AOI22_X1 _24558_ (.A1(\core.keymem.key_mem[3][110] ),
    .A2(_16384_),
    .B1(_16466_),
    .B2(\core.keymem.key_mem[5][110] ),
    .ZN(_18468_));
 AOI21_X1 _24559_ (.A(_16493_),
    .B1(_16523_),
    .B2(\core.keymem.key_mem[1][110] ),
    .ZN(_18469_));
 AOI22_X1 _24560_ (.A1(\core.keymem.key_mem[6][110] ),
    .A2(_16519_),
    .B1(_16440_),
    .B2(\core.keymem.key_mem[11][110] ),
    .ZN(_18470_));
 AOI22_X1 _24561_ (.A1(\core.keymem.key_mem[8][110] ),
    .A2(_16450_),
    .B1(_16430_),
    .B2(\core.keymem.key_mem[10][110] ),
    .ZN(_18471_));
 AND4_X1 _24562_ (.A1(_18468_),
    .A2(_18469_),
    .A3(_18470_),
    .A4(_18471_),
    .ZN(_18472_));
 AOI222_X2 _24563_ (.A1(\core.keymem.key_mem[14][110] ),
    .A2(_16436_),
    .B1(_16459_),
    .B2(\core.keymem.key_mem[9][110] ),
    .C1(_16395_),
    .C2(\core.keymem.key_mem[12][110] ),
    .ZN(_18473_));
 AOI22_X1 _24564_ (.A1(\core.keymem.key_mem[4][110] ),
    .A2(_16455_),
    .B1(_16470_),
    .B2(\core.keymem.key_mem[13][110] ),
    .ZN(_18474_));
 AOI22_X1 _24565_ (.A1(\core.keymem.key_mem[7][110] ),
    .A2(_16954_),
    .B1(_16422_),
    .B2(\core.keymem.key_mem[2][110] ),
    .ZN(_18475_));
 AND3_X1 _24566_ (.A1(_18473_),
    .A2(_18474_),
    .A3(_18475_),
    .ZN(_18476_));
 AOI22_X4 _24567_ (.A1(_00192_),
    .A2(_16982_),
    .B1(_18472_),
    .B2(_18476_),
    .ZN(_18477_));
 XNOR2_X2 _24568_ (.A(_17246_),
    .B(_18477_),
    .ZN(_18478_));
 BUF_X4 _24569_ (.A(_16554_),
    .Z(_18479_));
 OAI221_X2 _24570_ (.A(_18329_),
    .B1(_18466_),
    .B2(_18467_),
    .C1(_18478_),
    .C2(_18479_),
    .ZN(_18480_));
 XNOR2_X2 _24571_ (.A(_17935_),
    .B(_18341_),
    .ZN(_18481_));
 XNOR2_X2 _24572_ (.A(_17552_),
    .B(_17811_),
    .ZN(_18482_));
 XOR2_X1 _24573_ (.A(_18283_),
    .B(_18482_),
    .Z(_18483_));
 XNOR2_X1 _24574_ (.A(_17658_),
    .B(_18483_),
    .ZN(_18484_));
 XNOR2_X2 _24575_ (.A(_18481_),
    .B(_18484_),
    .ZN(_18485_));
 XOR2_X2 _24576_ (.A(_17604_),
    .B(_18485_),
    .Z(_18486_));
 XNOR2_X2 _24577_ (.A(_17824_),
    .B(_18337_),
    .ZN(_18487_));
 XNOR2_X2 _24578_ (.A(_17574_),
    .B(_18487_),
    .ZN(_18488_));
 XNOR2_X2 _24579_ (.A(_17761_),
    .B(_18310_),
    .ZN(_18489_));
 XOR2_X2 _24580_ (.A(_18488_),
    .B(_18489_),
    .Z(_18490_));
 XNOR2_X1 _24581_ (.A(_18486_),
    .B(_18490_),
    .ZN(_18491_));
 AOI21_X1 _24582_ (.A(_18480_),
    .B1(_18491_),
    .B2(_17749_),
    .ZN(_18492_));
 AOI21_X1 _24583_ (.A(_18415_),
    .B1(_18465_),
    .B2(_18492_),
    .ZN(_00572_));
 NOR2_X1 _24584_ (.A1(\core.dec_block.block_w0_reg[15] ),
    .A2(_18330_),
    .ZN(_18493_));
 INV_X1 _24585_ (.A(_18143_),
    .ZN(_18494_));
 NAND2_X1 _24586_ (.A1(_17279_),
    .A2(_17346_),
    .ZN(_18495_));
 AOI21_X1 _24587_ (.A(_18036_),
    .B1(_18495_),
    .B2(_17418_),
    .ZN(_18496_));
 AOI21_X1 _24588_ (.A(_17404_),
    .B1(_17306_),
    .B2(_17281_),
    .ZN(_18497_));
 OAI21_X1 _24589_ (.A(_18038_),
    .B1(_18497_),
    .B2(_17273_),
    .ZN(_18498_));
 OAI21_X1 _24590_ (.A(_18017_),
    .B1(_18496_),
    .B2(_18498_),
    .ZN(_18499_));
 NAND2_X1 _24591_ (.A1(_17212_),
    .A2(_17276_),
    .ZN(_18500_));
 MUX2_X1 _24592_ (.A(_17326_),
    .B(_18500_),
    .S(_17271_),
    .Z(_18501_));
 AOI22_X1 _24593_ (.A1(_17294_),
    .A2(_17456_),
    .B1(_17434_),
    .B2(_17496_),
    .ZN(_18502_));
 OAI22_X2 _24594_ (.A1(_18093_),
    .A2(_18501_),
    .B1(_18502_),
    .B2(_17987_),
    .ZN(_18503_));
 MUX2_X1 _24595_ (.A(_17346_),
    .B(_17496_),
    .S(_17434_),
    .Z(_18504_));
 OAI21_X1 _24596_ (.A(_18393_),
    .B1(_17298_),
    .B2(_17965_),
    .ZN(_18505_));
 AOI221_X2 _24597_ (.A(_18503_),
    .B1(_18504_),
    .B2(_17377_),
    .C1(_17381_),
    .C2(_18505_),
    .ZN(_18506_));
 NAND4_X1 _24598_ (.A1(_18494_),
    .A2(_18395_),
    .A3(_18499_),
    .A4(_18506_),
    .ZN(_18507_));
 OAI21_X1 _24599_ (.A(_18127_),
    .B1(_17439_),
    .B2(_17429_),
    .ZN(_18508_));
 OAI21_X1 _24600_ (.A(_17418_),
    .B1(_17317_),
    .B2(_17305_),
    .ZN(_18509_));
 OAI21_X1 _24601_ (.A(_17305_),
    .B1(_17353_),
    .B2(_17338_),
    .ZN(_18510_));
 OAI221_X2 _24602_ (.A(_17461_),
    .B1(_17474_),
    .B2(_17326_),
    .C1(_17308_),
    .C2(_17393_),
    .ZN(_18511_));
 AOI222_X2 _24603_ (.A1(_17255_),
    .A2(_18014_),
    .B1(_18509_),
    .B2(_18510_),
    .C1(_18511_),
    .C2(_17302_),
    .ZN(_18512_));
 INV_X1 _24604_ (.A(_18512_),
    .ZN(_18513_));
 OAI21_X1 _24605_ (.A(_17429_),
    .B1(_17461_),
    .B2(_17316_),
    .ZN(_18514_));
 AOI221_X1 _24606_ (.A(_17221_),
    .B1(_17965_),
    .B2(_18514_),
    .C1(_17456_),
    .C2(_17374_),
    .ZN(_18515_));
 NAND2_X1 _24607_ (.A1(_17397_),
    .A2(_17474_),
    .ZN(_18516_));
 AOI221_X1 _24608_ (.A(_18017_),
    .B1(_17294_),
    .B2(_18516_),
    .C1(_17384_),
    .C2(_17374_),
    .ZN(_18517_));
 NOR3_X1 _24609_ (.A1(_18164_),
    .A2(_18515_),
    .A3(_18517_),
    .ZN(_18518_));
 NOR4_X1 _24610_ (.A1(_18507_),
    .A2(_18508_),
    .A3(_18513_),
    .A4(_18518_),
    .ZN(_18519_));
 AOI21_X1 _24611_ (.A(_17364_),
    .B1(_17360_),
    .B2(_17374_),
    .ZN(_18520_));
 NOR2_X1 _24612_ (.A1(_17965_),
    .A2(_17369_),
    .ZN(_18521_));
 AOI21_X1 _24613_ (.A(_18520_),
    .B1(_18521_),
    .B2(_18161_),
    .ZN(_18522_));
 AOI21_X2 _24614_ (.A(_17490_),
    .B1(_18522_),
    .B2(_17321_),
    .ZN(_18523_));
 NOR2_X1 _24615_ (.A1(_18042_),
    .A2(_18205_),
    .ZN(_18524_));
 AND4_X1 _24616_ (.A1(_17395_),
    .A2(_18451_),
    .A3(_18456_),
    .A4(_18524_),
    .ZN(_18525_));
 AND3_X2 _24617_ (.A1(_18519_),
    .A2(_18523_),
    .A3(_18525_),
    .ZN(_18526_));
 AND2_X1 _24618_ (.A1(_00198_),
    .A2(_16495_),
    .ZN(_18527_));
 NAND3_X1 _24619_ (.A1(\core.keymem.key_mem[12][111] ),
    .A2(_17024_),
    .A3(_17527_),
    .ZN(_18528_));
 OAI211_X2 _24620_ (.A(\core.keymem.key_mem[6][111] ),
    .B(_17163_),
    .C1(_17031_),
    .C2(_16896_),
    .ZN(_18529_));
 NAND3_X1 _24621_ (.A1(\core.keymem.key_mem[3][111] ),
    .A2(_17074_),
    .A3(_17827_),
    .ZN(_18530_));
 NAND3_X1 _24622_ (.A1(\core.keymem.key_mem[2][111] ),
    .A2(_17827_),
    .A3(_17163_),
    .ZN(_18531_));
 NAND4_X2 _24623_ (.A1(_18528_),
    .A2(_18529_),
    .A3(_18530_),
    .A4(_18531_),
    .ZN(_18532_));
 OAI221_X2 _24624_ (.A(\core.keymem.key_mem[5][111] ),
    .B1(_16933_),
    .B2(_16934_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_18533_));
 OAI211_X2 _24625_ (.A(\core.keymem.key_mem[13][111] ),
    .B(_16919_),
    .C1(_16913_),
    .C2(_16915_),
    .ZN(_18534_));
 OAI211_X2 _24626_ (.A(\core.keymem.key_mem[8][111] ),
    .B(_16931_),
    .C1(_16927_),
    .C2(_16929_),
    .ZN(_18535_));
 OAI211_X2 _24627_ (.A(\core.keymem.key_mem[10][111] ),
    .B(_17015_),
    .C1(_16922_),
    .C2(_16923_),
    .ZN(_18536_));
 NAND4_X2 _24628_ (.A1(_18533_),
    .A2(_18534_),
    .A3(_18535_),
    .A4(_18536_),
    .ZN(_18537_));
 OAI211_X2 _24629_ (.A(\core.keymem.key_mem[4][111] ),
    .B(_16931_),
    .C1(_16908_),
    .C2(_16917_),
    .ZN(_18538_));
 OAI211_X2 _24630_ (.A(\core.keymem.key_mem[11][111] ),
    .B(_16901_),
    .C1(_16922_),
    .C2(_16923_),
    .ZN(_18539_));
 NAND3_X1 _24631_ (.A1(\core.keymem.key_mem[14][111] ),
    .A2(_16881_),
    .A3(_17015_),
    .ZN(_18540_));
 OAI221_X2 _24632_ (.A(\core.keymem.key_mem[9][111] ),
    .B1(_16926_),
    .B2(_16928_),
    .C1(_17018_),
    .C2(_17020_),
    .ZN(_18541_));
 NAND4_X2 _24633_ (.A1(_18538_),
    .A2(_18539_),
    .A3(_18540_),
    .A4(_18541_),
    .ZN(_18542_));
 INV_X1 _24634_ (.A(\core.keymem.key_mem[7][111] ),
    .ZN(_18543_));
 OAI21_X4 _24635_ (.A(_16481_),
    .B1(_16895_),
    .B2(_16898_),
    .ZN(_18544_));
 OAI21_X4 _24636_ (.A(_16969_),
    .B1(_17018_),
    .B2(_17020_),
    .ZN(_18545_));
 INV_X1 _24637_ (.A(\core.keymem.key_mem[1][111] ),
    .ZN(_18546_));
 OAI22_X4 _24638_ (.A1(_18543_),
    .A2(_18544_),
    .B1(_18545_),
    .B2(_18546_),
    .ZN(_18547_));
 NOR4_X4 _24639_ (.A1(_18532_),
    .A2(_18537_),
    .A3(_18542_),
    .A4(_18547_),
    .ZN(_18548_));
 AOI21_X4 _24640_ (.A(_18527_),
    .B1(_18548_),
    .B2(_16488_),
    .ZN(_18549_));
 XNOR2_X2 _24641_ (.A(\core.dec_block.block_w0_reg[15] ),
    .B(_18549_),
    .ZN(_18550_));
 XNOR2_X2 _24642_ (.A(\block_reg[2][15] ),
    .B(_17847_),
    .ZN(_18551_));
 BUF_X4 _24643_ (.A(_17709_),
    .Z(_18552_));
 BUF_X4 _24644_ (.A(_18552_),
    .Z(_18553_));
 OAI221_X2 _24645_ (.A(_18329_),
    .B1(_17741_),
    .B2(_18550_),
    .C1(_18551_),
    .C2(_18553_),
    .ZN(_18554_));
 XNOR2_X2 _24646_ (.A(_17552_),
    .B(_18297_),
    .ZN(_18555_));
 XNOR2_X1 _24647_ (.A(_17518_),
    .B(_18282_),
    .ZN(_18556_));
 XNOR2_X2 _24648_ (.A(_17946_),
    .B(_18310_),
    .ZN(_18557_));
 XNOR2_X1 _24649_ (.A(_18556_),
    .B(_18557_),
    .ZN(_18558_));
 XNOR2_X2 _24650_ (.A(_18555_),
    .B(_18558_),
    .ZN(_18559_));
 XNOR2_X2 _24651_ (.A(_17702_),
    .B(_17824_),
    .ZN(_18560_));
 XOR2_X1 _24652_ (.A(_18338_),
    .B(_18560_),
    .Z(_18561_));
 XNOR2_X1 _24653_ (.A(_17658_),
    .B(_18561_),
    .ZN(_18562_));
 XNOR2_X1 _24654_ (.A(_18559_),
    .B(_18562_),
    .ZN(_18563_));
 AOI21_X1 _24655_ (.A(_18554_),
    .B1(_18563_),
    .B2(_17749_),
    .ZN(_18564_));
 AOI21_X1 _24656_ (.A(_18493_),
    .B1(_18526_),
    .B2(_18564_),
    .ZN(_00573_));
 NOR2_X1 _24657_ (.A1(\core.dec_block.block_w0_reg[16] ),
    .A2(_18330_),
    .ZN(_18565_));
 BUF_X4 _24658_ (.A(_16358_),
    .Z(_18566_));
 NAND2_X1 _24659_ (.A1(_18566_),
    .A2(\core.dec_block.block_w0_reg[18] ),
    .ZN(_18567_));
 BUF_X4 _24660_ (.A(_16569_),
    .Z(_18568_));
 BUF_X4 _24661_ (.A(_16566_),
    .Z(_18569_));
 AOI222_X2 _24662_ (.A1(\core.dec_block.block_w1_reg[18] ),
    .A2(_18568_),
    .B1(_16268_),
    .B2(\core.dec_block.block_w3_reg[18] ),
    .C1(\core.dec_block.block_w2_reg[18] ),
    .C2(_18569_),
    .ZN(_18570_));
 OAI21_X2 _24663_ (.A(_18567_),
    .B1(_18570_),
    .B2(_16359_),
    .ZN(_18571_));
 NAND2_X4 _24664_ (.A1(_17329_),
    .A2(_18571_),
    .ZN(_18572_));
 BUF_X4 _24665_ (.A(_18572_),
    .Z(_18573_));
 CLKBUF_X3 _24666_ (.A(\core.dec_block.block_w0_reg[23] ),
    .Z(_18574_));
 NAND2_X1 _24667_ (.A1(_18566_),
    .A2(_18574_),
    .ZN(_18575_));
 BUF_X2 _24668_ (.A(\core.dec_block.block_w3_reg[23] ),
    .Z(_18576_));
 BUF_X2 _24669_ (.A(\core.dec_block.block_w1_reg[23] ),
    .Z(_18577_));
 AOI222_X2 _24670_ (.A1(_17537_),
    .A2(_18569_),
    .B1(_16268_),
    .B2(_18576_),
    .C1(_18568_),
    .C2(_18577_),
    .ZN(_18578_));
 OAI21_X2 _24671_ (.A(_18575_),
    .B1(_18578_),
    .B2(_16359_),
    .ZN(_18579_));
 NAND2_X2 _24672_ (.A1(_17329_),
    .A2(_18579_),
    .ZN(_18580_));
 BUF_X4 _24673_ (.A(_18580_),
    .Z(_18581_));
 NAND2_X1 _24674_ (.A1(\core.dec_block.block_w0_reg[22] ),
    .A2(_18566_),
    .ZN(_18582_));
 AOI222_X2 _24675_ (.A1(\core.dec_block.block_w2_reg[22] ),
    .A2(_18569_),
    .B1(_16268_),
    .B2(\core.dec_block.block_w3_reg[22] ),
    .C1(_18568_),
    .C2(\core.dec_block.block_w1_reg[22] ),
    .ZN(_18583_));
 OAI21_X2 _24676_ (.A(_18582_),
    .B1(_18583_),
    .B2(_16359_),
    .ZN(_18584_));
 NAND2_X4 _24677_ (.A1(_17329_),
    .A2(_18584_),
    .ZN(_18585_));
 NOR2_X4 _24678_ (.A1(_18581_),
    .A2(_18585_),
    .ZN(_18586_));
 NAND2_X1 _24679_ (.A1(_18566_),
    .A2(\core.dec_block.block_w0_reg[20] ),
    .ZN(_18587_));
 AOI222_X2 _24680_ (.A1(\core.dec_block.block_w1_reg[20] ),
    .A2(_18568_),
    .B1(_16267_),
    .B2(\core.dec_block.block_w3_reg[20] ),
    .C1(\core.dec_block.block_w2_reg[20] ),
    .C2(_18569_),
    .ZN(_18588_));
 OAI21_X2 _24681_ (.A(_18587_),
    .B1(_18588_),
    .B2(_16359_),
    .ZN(_18589_));
 AND2_X1 _24682_ (.A1(_16562_),
    .A2(_18589_),
    .ZN(_18590_));
 BUF_X4 _24683_ (.A(_18590_),
    .Z(_18591_));
 NAND2_X1 _24684_ (.A1(\core.dec_block.block_w0_reg[21] ),
    .A2(_18566_),
    .ZN(_18592_));
 AOI222_X2 _24685_ (.A1(\core.dec_block.block_w2_reg[21] ),
    .A2(_18569_),
    .B1(_16267_),
    .B2(\core.dec_block.block_w3_reg[21] ),
    .C1(_18568_),
    .C2(\core.dec_block.block_w1_reg[21] ),
    .ZN(_18593_));
 OAI21_X2 _24686_ (.A(_18592_),
    .B1(_18593_),
    .B2(_18566_),
    .ZN(_18594_));
 AND2_X1 _24687_ (.A1(_16562_),
    .A2(_18594_),
    .ZN(_18595_));
 BUF_X4 _24688_ (.A(_18595_),
    .Z(_18596_));
 NOR2_X4 _24689_ (.A1(_18591_),
    .A2(_18596_),
    .ZN(_18597_));
 NAND2_X4 _24690_ (.A1(_18586_),
    .A2(_18597_),
    .ZN(_18598_));
 NOR2_X1 _24691_ (.A1(_18573_),
    .A2(_18598_),
    .ZN(_18599_));
 NAND2_X1 _24692_ (.A1(_16359_),
    .A2(\core.dec_block.block_w0_reg[17] ),
    .ZN(_18600_));
 AOI222_X2 _24693_ (.A1(\core.dec_block.block_w1_reg[17] ),
    .A2(_18568_),
    .B1(_16268_),
    .B2(\core.dec_block.block_w3_reg[17] ),
    .C1(\core.dec_block.block_w2_reg[17] ),
    .C2(_18569_),
    .ZN(_18601_));
 OAI21_X2 _24694_ (.A(_18600_),
    .B1(_18601_),
    .B2(_16359_),
    .ZN(_18602_));
 AND2_X2 _24695_ (.A1(_17329_),
    .A2(_18602_),
    .ZN(_18603_));
 NAND2_X1 _24696_ (.A1(\core.dec_block.block_w0_reg[16] ),
    .A2(_18566_),
    .ZN(_18604_));
 AOI222_X2 _24697_ (.A1(\core.dec_block.block_w1_reg[16] ),
    .A2(_18568_),
    .B1(_16268_),
    .B2(\core.dec_block.block_w3_reg[16] ),
    .C1(\core.dec_block.block_w2_reg[16] ),
    .C2(_18569_),
    .ZN(_18605_));
 OAI21_X2 _24698_ (.A(_18604_),
    .B1(_18605_),
    .B2(_16359_),
    .ZN(_18606_));
 NAND2_X4 _24699_ (.A1(_17329_),
    .A2(_18606_),
    .ZN(_18607_));
 NOR2_X2 _24700_ (.A1(_18603_),
    .A2(_18607_),
    .ZN(_18608_));
 BUF_X4 _24701_ (.A(_18608_),
    .Z(_18609_));
 NAND2_X2 _24702_ (.A1(_17329_),
    .A2(_18602_),
    .ZN(_18610_));
 AND2_X1 _24703_ (.A1(_16622_),
    .A2(_18606_),
    .ZN(_18611_));
 BUF_X8 _24704_ (.A(_18611_),
    .Z(_18612_));
 NOR2_X4 _24705_ (.A1(_18610_),
    .A2(_18612_),
    .ZN(_18613_));
 NOR2_X2 _24706_ (.A1(_18613_),
    .A2(_18608_),
    .ZN(_18614_));
 NAND2_X1 _24707_ (.A1(_18566_),
    .A2(\core.dec_block.block_w0_reg[19] ),
    .ZN(_18615_));
 AOI222_X2 _24708_ (.A1(\core.dec_block.block_w1_reg[19] ),
    .A2(_18568_),
    .B1(_16268_),
    .B2(\core.dec_block.block_w3_reg[19] ),
    .C1(\core.dec_block.block_w2_reg[19] ),
    .C2(_18569_),
    .ZN(_18616_));
 OAI21_X2 _24709_ (.A(_18615_),
    .B1(_18616_),
    .B2(_16359_),
    .ZN(_18617_));
 AND2_X1 _24710_ (.A1(_16622_),
    .A2(_18617_),
    .ZN(_18618_));
 BUF_X4 _24711_ (.A(_18618_),
    .Z(_18619_));
 BUF_X4 _24712_ (.A(_18619_),
    .Z(_18620_));
 BUF_X4 _24713_ (.A(_18620_),
    .Z(_18621_));
 MUX2_X1 _24714_ (.A(_18609_),
    .B(_18614_),
    .S(_18621_),
    .Z(_18622_));
 BUF_X4 _24715_ (.A(_18603_),
    .Z(_18623_));
 NAND2_X4 _24716_ (.A1(_18416_),
    .A2(_18617_),
    .ZN(_18624_));
 AND2_X1 _24717_ (.A1(_16622_),
    .A2(_18571_),
    .ZN(_18625_));
 BUF_X4 _24718_ (.A(_18625_),
    .Z(_18626_));
 NAND2_X2 _24719_ (.A1(_18624_),
    .A2(_18626_),
    .ZN(_18627_));
 NOR2_X4 _24720_ (.A1(_18623_),
    .A2(_18627_),
    .ZN(_18628_));
 BUF_X4 _24721_ (.A(_18591_),
    .Z(_18629_));
 NAND2_X2 _24722_ (.A1(_16622_),
    .A2(_18594_),
    .ZN(_18630_));
 BUF_X4 _24723_ (.A(_18630_),
    .Z(_18631_));
 AND2_X2 _24724_ (.A1(_16622_),
    .A2(_18584_),
    .ZN(_18632_));
 BUF_X4 _24725_ (.A(_18632_),
    .Z(_18633_));
 NOR2_X4 _24726_ (.A1(_18581_),
    .A2(_18633_),
    .ZN(_18634_));
 NAND2_X4 _24727_ (.A1(_18631_),
    .A2(_18634_),
    .ZN(_18635_));
 NOR2_X2 _24728_ (.A1(_18629_),
    .A2(_18635_),
    .ZN(_18636_));
 AOI22_X1 _24729_ (.A1(_18599_),
    .A2(_18622_),
    .B1(_18628_),
    .B2(_18636_),
    .ZN(_18637_));
 NAND2_X2 _24730_ (.A1(_18619_),
    .A2(_18572_),
    .ZN(_18638_));
 BUF_X4 _24731_ (.A(_18638_),
    .Z(_18639_));
 CLKBUF_X3 _24732_ (.A(_18639_),
    .Z(_18640_));
 NAND2_X2 _24733_ (.A1(_17329_),
    .A2(_18589_),
    .ZN(_18641_));
 BUF_X4 _24734_ (.A(_18641_),
    .Z(_18642_));
 NAND2_X4 _24735_ (.A1(_18642_),
    .A2(_18596_),
    .ZN(_18643_));
 AND2_X1 _24736_ (.A1(_16622_),
    .A2(_18579_),
    .ZN(_18644_));
 BUF_X4 _24737_ (.A(_18644_),
    .Z(_18645_));
 NAND2_X4 _24738_ (.A1(_18645_),
    .A2(_18632_),
    .ZN(_18646_));
 NOR2_X4 _24739_ (.A1(_18643_),
    .A2(_18646_),
    .ZN(_18647_));
 BUF_X4 _24740_ (.A(_18612_),
    .Z(_18648_));
 NOR2_X4 _24741_ (.A1(_18642_),
    .A2(_18596_),
    .ZN(_18649_));
 NOR2_X4 _24742_ (.A1(_18645_),
    .A2(_18632_),
    .ZN(_18650_));
 NAND2_X4 _24743_ (.A1(_18649_),
    .A2(_18650_),
    .ZN(_18651_));
 NOR2_X2 _24744_ (.A1(_18648_),
    .A2(_18651_),
    .ZN(_18652_));
 BUF_X4 _24745_ (.A(_18623_),
    .Z(_18653_));
 BUF_X4 _24746_ (.A(_18653_),
    .Z(_18654_));
 BUF_X4 _24747_ (.A(_18654_),
    .Z(_18655_));
 AOI22_X1 _24748_ (.A1(_18647_),
    .A2(_18609_),
    .B1(_18652_),
    .B2(_18655_),
    .ZN(_18656_));
 OAI21_X1 _24749_ (.A(_18637_),
    .B1(_18640_),
    .B2(_18656_),
    .ZN(_18657_));
 BUF_X4 _24750_ (.A(_18624_),
    .Z(_18658_));
 BUF_X4 _24751_ (.A(_18658_),
    .Z(_18659_));
 NAND2_X4 _24752_ (.A1(_18580_),
    .A2(_18632_),
    .ZN(_18660_));
 NOR2_X1 _24753_ (.A1(_18643_),
    .A2(_18660_),
    .ZN(_18661_));
 BUF_X4 _24754_ (.A(_18661_),
    .Z(_18662_));
 OAI21_X1 _24755_ (.A(_18659_),
    .B1(_18662_),
    .B2(_18599_),
    .ZN(_18663_));
 NOR2_X4 _24756_ (.A1(_18591_),
    .A2(_18631_),
    .ZN(_18664_));
 NAND2_X2 _24757_ (.A1(_18664_),
    .A2(_18586_),
    .ZN(_18665_));
 BUF_X4 _24758_ (.A(_18665_),
    .Z(_18666_));
 OAI21_X1 _24759_ (.A(_18663_),
    .B1(_18640_),
    .B2(_18666_),
    .ZN(_18667_));
 BUF_X4 _24760_ (.A(_18613_),
    .Z(_18668_));
 AOI21_X2 _24761_ (.A(_18657_),
    .B1(_18667_),
    .B2(_18668_),
    .ZN(_18669_));
 BUF_X4 _24762_ (.A(_18627_),
    .Z(_18670_));
 NAND2_X1 _24763_ (.A1(_18664_),
    .A2(_18634_),
    .ZN(_18671_));
 BUF_X4 _24764_ (.A(_18671_),
    .Z(_18672_));
 AOI21_X2 _24765_ (.A(_18670_),
    .B1(_18651_),
    .B2(_18672_),
    .ZN(_18673_));
 NAND2_X4 _24766_ (.A1(_18619_),
    .A2(_18626_),
    .ZN(_18674_));
 BUF_X4 _24767_ (.A(_18610_),
    .Z(_18675_));
 NAND2_X4 _24768_ (.A1(_18675_),
    .A2(_18612_),
    .ZN(_18676_));
 NOR2_X4 _24769_ (.A1(_18674_),
    .A2(_18676_),
    .ZN(_18677_));
 NAND2_X4 _24770_ (.A1(_18645_),
    .A2(_18585_),
    .ZN(_18678_));
 NAND2_X4 _24771_ (.A1(_18591_),
    .A2(_18596_),
    .ZN(_18679_));
 NOR2_X4 _24772_ (.A1(_18678_),
    .A2(_18679_),
    .ZN(_18680_));
 NAND2_X4 _24773_ (.A1(_18610_),
    .A2(_18607_),
    .ZN(_18681_));
 NOR2_X4 _24774_ (.A1(_18638_),
    .A2(_18681_),
    .ZN(_18682_));
 AOI221_X1 _24775_ (.A(_18673_),
    .B1(_18677_),
    .B2(_18680_),
    .C1(_18662_),
    .C2(_18682_),
    .ZN(_18683_));
 NAND2_X4 _24776_ (.A1(_18591_),
    .A2(_18630_),
    .ZN(_18684_));
 NOR2_X2 _24777_ (.A1(_18646_),
    .A2(_18684_),
    .ZN(_18685_));
 BUF_X4 _24778_ (.A(_18685_),
    .Z(_18686_));
 NOR2_X1 _24779_ (.A1(_18686_),
    .A2(_18652_),
    .ZN(_18687_));
 NOR2_X4 _24780_ (.A1(_18619_),
    .A2(_18626_),
    .ZN(_18688_));
 NAND2_X4 _24781_ (.A1(_18623_),
    .A2(_18688_),
    .ZN(_18689_));
 OAI21_X1 _24782_ (.A(_18683_),
    .B1(_18687_),
    .B2(_18689_),
    .ZN(_18690_));
 NOR2_X4 _24783_ (.A1(_18596_),
    .A2(_18678_),
    .ZN(_18691_));
 NAND2_X4 _24784_ (.A1(_18642_),
    .A2(_18691_),
    .ZN(_18692_));
 BUF_X4 _24785_ (.A(_18692_),
    .Z(_18693_));
 NAND2_X4 _24786_ (.A1(_18623_),
    .A2(_18607_),
    .ZN(_18694_));
 NOR2_X4 _24787_ (.A1(_18645_),
    .A2(_18585_),
    .ZN(_18695_));
 NAND2_X4 _24788_ (.A1(_18695_),
    .A2(_18649_),
    .ZN(_18696_));
 BUF_X4 _24789_ (.A(_18607_),
    .Z(_18697_));
 BUF_X4 _24790_ (.A(_18697_),
    .Z(_18698_));
 BUF_X4 _24791_ (.A(_18698_),
    .Z(_18699_));
 BUF_X4 _24792_ (.A(_18699_),
    .Z(_18700_));
 OAI22_X1 _24793_ (.A1(_18693_),
    .A2(_18694_),
    .B1(_18696_),
    .B2(_18700_),
    .ZN(_18701_));
 NOR2_X4 _24794_ (.A1(_18624_),
    .A2(_18626_),
    .ZN(_18702_));
 BUF_X4 _24795_ (.A(_18702_),
    .Z(_18703_));
 AOI21_X1 _24796_ (.A(_18690_),
    .B1(_18701_),
    .B2(_18703_),
    .ZN(_18704_));
 NAND2_X2 _24797_ (.A1(_18675_),
    .A2(_18688_),
    .ZN(_18705_));
 NAND2_X4 _24798_ (.A1(_18580_),
    .A2(_18585_),
    .ZN(_18706_));
 NOR2_X2 _24799_ (.A1(_18684_),
    .A2(_18706_),
    .ZN(_18707_));
 BUF_X4 _24800_ (.A(_18707_),
    .Z(_18708_));
 NAND2_X1 _24801_ (.A1(_18648_),
    .A2(_18708_),
    .ZN(_18709_));
 NAND2_X4 _24802_ (.A1(_18642_),
    .A2(_18631_),
    .ZN(_18710_));
 NOR2_X4 _24803_ (.A1(_18646_),
    .A2(_18710_),
    .ZN(_18711_));
 NOR2_X4 _24804_ (.A1(_18646_),
    .A2(_18679_),
    .ZN(_18712_));
 NOR2_X1 _24805_ (.A1(_18711_),
    .A2(_18712_),
    .ZN(_18713_));
 AOI21_X1 _24806_ (.A(_18705_),
    .B1(_18709_),
    .B2(_18713_),
    .ZN(_18714_));
 CLKBUF_X3 _24807_ (.A(_18573_),
    .Z(_18715_));
 CLKBUF_X3 _24808_ (.A(_18715_),
    .Z(_18716_));
 NOR2_X4 _24809_ (.A1(_18603_),
    .A2(_18612_),
    .ZN(_18717_));
 NAND2_X4 _24810_ (.A1(_18603_),
    .A2(_18612_),
    .ZN(_18718_));
 BUF_X4 _24811_ (.A(_18718_),
    .Z(_18719_));
 AOI21_X1 _24812_ (.A(_18717_),
    .B1(_18719_),
    .B2(_18658_),
    .ZN(_18720_));
 NAND2_X2 _24813_ (.A1(_18597_),
    .A2(_18650_),
    .ZN(_18721_));
 BUF_X4 _24814_ (.A(_18721_),
    .Z(_18722_));
 BUF_X4 _24815_ (.A(_18648_),
    .Z(_18723_));
 OAI33_X1 _24816_ (.A1(_18716_),
    .A2(_18696_),
    .A3(_18720_),
    .B1(_18722_),
    .B2(_18640_),
    .B3(_18723_),
    .ZN(_18724_));
 NAND2_X2 _24817_ (.A1(_18612_),
    .A2(_18688_),
    .ZN(_18725_));
 NOR2_X4 _24818_ (.A1(_18643_),
    .A2(_18706_),
    .ZN(_18726_));
 NAND2_X2 _24819_ (.A1(_18675_),
    .A2(_18726_),
    .ZN(_18727_));
 NOR2_X2 _24820_ (.A1(_18675_),
    .A2(_18607_),
    .ZN(_18728_));
 NAND2_X2 _24821_ (.A1(_18702_),
    .A2(_18728_),
    .ZN(_18729_));
 OAI22_X4 _24822_ (.A1(_18725_),
    .A2(_18727_),
    .B1(_18729_),
    .B2(_18598_),
    .ZN(_18730_));
 NOR2_X4 _24823_ (.A1(_18641_),
    .A2(_18631_),
    .ZN(_18731_));
 NAND2_X2 _24824_ (.A1(_18731_),
    .A2(_18650_),
    .ZN(_18732_));
 BUF_X4 _24825_ (.A(_18732_),
    .Z(_18733_));
 OAI33_X1 _24826_ (.A1(_18598_),
    .A2(_18640_),
    .A3(_18681_),
    .B1(_18733_),
    .B2(_18689_),
    .B3(_18723_),
    .ZN(_18734_));
 NOR4_X2 _24827_ (.A1(_18714_),
    .A2(_18724_),
    .A3(_18730_),
    .A4(_18734_),
    .ZN(_18735_));
 BUF_X4 _24828_ (.A(_18728_),
    .Z(_18736_));
 NAND3_X1 _24829_ (.A1(_18658_),
    .A2(_18711_),
    .A3(_18736_),
    .ZN(_18737_));
 CLKBUF_X3 _24830_ (.A(_18624_),
    .Z(_18738_));
 NOR3_X1 _24831_ (.A1(_18738_),
    .A2(_18642_),
    .A3(_18614_),
    .ZN(_18739_));
 NOR2_X4 _24832_ (.A1(_18648_),
    .A2(_18689_),
    .ZN(_18740_));
 CLKBUF_X3 _24833_ (.A(_18642_),
    .Z(_18741_));
 AOI21_X1 _24834_ (.A(_18739_),
    .B1(_18740_),
    .B2(_18741_),
    .ZN(_18742_));
 NAND2_X2 _24835_ (.A1(_18586_),
    .A2(_18649_),
    .ZN(_18743_));
 BUF_X4 _24836_ (.A(_18743_),
    .Z(_18744_));
 BUF_X4 _24837_ (.A(_18675_),
    .Z(_18745_));
 NOR2_X4 _24838_ (.A1(_18619_),
    .A2(_18572_),
    .ZN(_18746_));
 NAND2_X2 _24839_ (.A1(_18745_),
    .A2(_18746_),
    .ZN(_18747_));
 OAI221_X2 _24840_ (.A(_18737_),
    .B1(_18742_),
    .B2(_18635_),
    .C1(_18744_),
    .C2(_18747_),
    .ZN(_18748_));
 NAND2_X4 _24841_ (.A1(_18609_),
    .A2(_18688_),
    .ZN(_18749_));
 CLKBUF_X3 _24842_ (.A(_18596_),
    .Z(_18750_));
 OAI22_X1 _24843_ (.A1(_18674_),
    .A2(_18719_),
    .B1(_18749_),
    .B2(_18750_),
    .ZN(_18751_));
 NOR2_X1 _24844_ (.A1(_18642_),
    .A2(_18585_),
    .ZN(_18752_));
 NOR2_X2 _24845_ (.A1(_18674_),
    .A2(_18718_),
    .ZN(_18753_));
 MUX2_X1 _24846_ (.A(_18682_),
    .B(_18753_),
    .S(_18750_),
    .Z(_18754_));
 NOR2_X1 _24847_ (.A1(_18591_),
    .A2(_18633_),
    .ZN(_18755_));
 AOI22_X1 _24848_ (.A1(_18751_),
    .A2(_18752_),
    .B1(_18754_),
    .B2(_18755_),
    .ZN(_18756_));
 NOR2_X1 _24849_ (.A1(_18581_),
    .A2(_18756_),
    .ZN(_18757_));
 NAND2_X2 _24850_ (.A1(_18695_),
    .A2(_18731_),
    .ZN(_18758_));
 NOR3_X1 _24851_ (.A1(_18758_),
    .A2(_18614_),
    .A3(_18670_),
    .ZN(_18759_));
 NOR2_X2 _24852_ (.A1(_18694_),
    .A2(_18627_),
    .ZN(_18760_));
 NOR2_X4 _24853_ (.A1(_18639_),
    .A2(_18718_),
    .ZN(_18761_));
 AOI221_X2 _24854_ (.A(_18759_),
    .B1(_18760_),
    .B2(_18647_),
    .C1(_18662_),
    .C2(_18761_),
    .ZN(_18762_));
 BUF_X4 _24855_ (.A(_18626_),
    .Z(_18763_));
 NOR2_X1 _24856_ (.A1(_18660_),
    .A2(_18710_),
    .ZN(_18764_));
 BUF_X4 _24857_ (.A(_18764_),
    .Z(_18765_));
 NAND2_X2 _24858_ (.A1(_18763_),
    .A2(_18765_),
    .ZN(_18766_));
 INV_X1 _24859_ (.A(_18766_),
    .ZN(_18767_));
 NOR2_X4 _24860_ (.A1(_18643_),
    .A2(_18678_),
    .ZN(_18768_));
 AOI21_X2 _24861_ (.A(_18767_),
    .B1(_18768_),
    .B2(_18715_),
    .ZN(_18769_));
 NAND2_X4 _24862_ (.A1(_18620_),
    .A2(_18745_),
    .ZN(_18770_));
 AOI22_X1 _24863_ (.A1(_18694_),
    .A2(_18703_),
    .B1(_18736_),
    .B2(_18746_),
    .ZN(_18771_));
 OAI221_X2 _24864_ (.A(_18762_),
    .B1(_18769_),
    .B2(_18770_),
    .C1(_18771_),
    .C2(_18744_),
    .ZN(_18772_));
 NAND2_X2 _24865_ (.A1(_18624_),
    .A2(_18572_),
    .ZN(_18773_));
 NOR2_X4 _24866_ (.A1(_18607_),
    .A2(_18773_),
    .ZN(_18774_));
 NAND2_X1 _24867_ (.A1(_18653_),
    .A2(_18774_),
    .ZN(_18775_));
 NAND2_X2 _24868_ (.A1(_18613_),
    .A2(_18746_),
    .ZN(_18776_));
 OAI21_X1 _24869_ (.A(_18775_),
    .B1(_18776_),
    .B2(_18722_),
    .ZN(_18777_));
 NOR2_X4 _24870_ (.A1(_18710_),
    .A2(_18706_),
    .ZN(_18778_));
 NOR2_X4 _24871_ (.A1(_18660_),
    .A2(_18679_),
    .ZN(_18779_));
 CLKBUF_X3 _24872_ (.A(_18779_),
    .Z(_18780_));
 OAI21_X1 _24873_ (.A(_18777_),
    .B1(_18778_),
    .B2(_18780_),
    .ZN(_18781_));
 BUF_X4 _24874_ (.A(_18674_),
    .Z(_18782_));
 BUF_X4 _24875_ (.A(_18726_),
    .Z(_18783_));
 AOI21_X1 _24876_ (.A(_18778_),
    .B1(_18783_),
    .B2(_18668_),
    .ZN(_18784_));
 OAI221_X2 _24877_ (.A(_18781_),
    .B1(_18749_),
    .B2(_18693_),
    .C1(_18782_),
    .C2(_18784_),
    .ZN(_18785_));
 NOR4_X2 _24878_ (.A1(_18748_),
    .A2(_18757_),
    .A3(_18772_),
    .A4(_18785_),
    .ZN(_18786_));
 NAND4_X2 _24879_ (.A1(_18669_),
    .A2(_18704_),
    .A3(_18735_),
    .A4(_18786_),
    .ZN(_18787_));
 BUF_X4 _24880_ (.A(_18621_),
    .Z(_18788_));
 BUF_X4 _24881_ (.A(_18788_),
    .Z(_18789_));
 NAND3_X1 _24882_ (.A1(_18623_),
    .A2(_18697_),
    .A3(_18680_),
    .ZN(_18790_));
 NAND3_X1 _24883_ (.A1(_18675_),
    .A2(_18612_),
    .A3(_18712_),
    .ZN(_18791_));
 AOI21_X1 _24884_ (.A(_18573_),
    .B1(_18790_),
    .B2(_18791_),
    .ZN(_18792_));
 NOR2_X4 _24885_ (.A1(_18626_),
    .A2(_18607_),
    .ZN(_18793_));
 NAND2_X2 _24886_ (.A1(_18634_),
    .A2(_18731_),
    .ZN(_18794_));
 OAI21_X1 _24887_ (.A(_18671_),
    .B1(_18794_),
    .B2(_18745_),
    .ZN(_18795_));
 BUF_X4 _24888_ (.A(_18745_),
    .Z(_18796_));
 NAND2_X1 _24889_ (.A1(_18626_),
    .A2(_18612_),
    .ZN(_18797_));
 OAI22_X1 _24890_ (.A1(_18763_),
    .A2(_18672_),
    .B1(_18733_),
    .B2(_18797_),
    .ZN(_18798_));
 AOI221_X1 _24891_ (.A(_18792_),
    .B1(_18793_),
    .B2(_18795_),
    .C1(_18796_),
    .C2(_18798_),
    .ZN(_18799_));
 OR2_X1 _24892_ (.A1(_18789_),
    .A2(_18799_),
    .ZN(_18800_));
 NAND2_X4 _24893_ (.A1(_18586_),
    .A2(_18731_),
    .ZN(_18801_));
 NOR2_X2 _24894_ (.A1(_18668_),
    .A2(_18801_),
    .ZN(_18802_));
 NOR2_X1 _24895_ (.A1(_18621_),
    .A2(_18693_),
    .ZN(_18803_));
 AOI22_X2 _24896_ (.A1(_18788_),
    .A2(_18802_),
    .B1(_18803_),
    .B2(_18736_),
    .ZN(_18804_));
 BUF_X4 _24897_ (.A(_18763_),
    .Z(_18805_));
 BUF_X4 _24898_ (.A(_18805_),
    .Z(_18806_));
 BUF_X4 _24899_ (.A(_18723_),
    .Z(_18807_));
 CLKBUF_X3 _24900_ (.A(_18796_),
    .Z(_18808_));
 NOR3_X1 _24901_ (.A1(_18715_),
    .A2(_18808_),
    .A3(_18758_),
    .ZN(_18809_));
 BUF_X4 _24902_ (.A(_18794_),
    .Z(_18810_));
 NOR3_X1 _24903_ (.A1(_18805_),
    .A2(_18655_),
    .A3(_18810_),
    .ZN(_18811_));
 OAI21_X1 _24904_ (.A(_18807_),
    .B1(_18809_),
    .B2(_18811_),
    .ZN(_18812_));
 OAI221_X2 _24905_ (.A(_18800_),
    .B1(_18804_),
    .B2(_18806_),
    .C1(_18659_),
    .C2(_18812_),
    .ZN(_18813_));
 NOR2_X1 _24906_ (.A1(_18624_),
    .A2(_18573_),
    .ZN(_18814_));
 BUF_X4 _24907_ (.A(_18814_),
    .Z(_18815_));
 BUF_X4 _24908_ (.A(_18745_),
    .Z(_18816_));
 CLKBUF_X3 _24909_ (.A(_18816_),
    .Z(_18817_));
 NOR2_X1 _24910_ (.A1(_18697_),
    .A2(_18692_),
    .ZN(_18818_));
 NAND2_X2 _24911_ (.A1(_18664_),
    .A2(_18695_),
    .ZN(_18819_));
 BUF_X4 _24912_ (.A(_18819_),
    .Z(_18820_));
 NOR2_X1 _24913_ (.A1(_18807_),
    .A2(_18820_),
    .ZN(_18821_));
 NOR3_X1 _24914_ (.A1(_18817_),
    .A2(_18818_),
    .A3(_18821_),
    .ZN(_18822_));
 BUF_X4 _24915_ (.A(_18654_),
    .Z(_18823_));
 NOR2_X1 _24916_ (.A1(_18698_),
    .A2(_18820_),
    .ZN(_18824_));
 NOR4_X1 _24917_ (.A1(_18823_),
    .A2(_18780_),
    .A3(_18686_),
    .A4(_18824_),
    .ZN(_18825_));
 OAI21_X1 _24918_ (.A(_18666_),
    .B1(_18822_),
    .B2(_18825_),
    .ZN(_18826_));
 NAND2_X1 _24919_ (.A1(_18815_),
    .A2(_18826_),
    .ZN(_18827_));
 AOI21_X1 _24920_ (.A(_18650_),
    .B1(_18745_),
    .B2(_18586_),
    .ZN(_18828_));
 NOR3_X1 _24921_ (.A1(_18738_),
    .A2(_18631_),
    .A3(_18828_),
    .ZN(_18829_));
 AOI21_X1 _24922_ (.A(_18829_),
    .B1(_18691_),
    .B2(_18658_),
    .ZN(_18830_));
 NAND3_X1 _24923_ (.A1(_18581_),
    .A2(_18585_),
    .A3(_18655_),
    .ZN(_18831_));
 CLKBUF_X3 _24924_ (.A(_18738_),
    .Z(_18832_));
 NAND2_X1 _24925_ (.A1(_18832_),
    .A2(_18664_),
    .ZN(_18833_));
 OAI221_X2 _24926_ (.A(_18806_),
    .B1(_18741_),
    .B2(_18830_),
    .C1(_18831_),
    .C2(_18833_),
    .ZN(_18834_));
 NAND3_X1 _24927_ (.A1(_18832_),
    .A2(_18609_),
    .A3(_18778_),
    .ZN(_18835_));
 AOI21_X1 _24928_ (.A(_18780_),
    .B1(_18783_),
    .B2(_18655_),
    .ZN(_18836_));
 OAI21_X1 _24929_ (.A(_18835_),
    .B1(_18836_),
    .B2(_18659_),
    .ZN(_18837_));
 OAI21_X1 _24930_ (.A(_18834_),
    .B1(_18837_),
    .B2(_18806_),
    .ZN(_18838_));
 NAND2_X1 _24931_ (.A1(_18827_),
    .A2(_18838_),
    .ZN(_18839_));
 NOR2_X2 _24932_ (.A1(_18648_),
    .A2(_18696_),
    .ZN(_18840_));
 OAI21_X1 _24933_ (.A(_18655_),
    .B1(_18708_),
    .B2(_18840_),
    .ZN(_18841_));
 NOR2_X4 _24934_ (.A1(_18660_),
    .A2(_18684_),
    .ZN(_18842_));
 NAND3_X1 _24935_ (.A1(_18808_),
    .A2(_18807_),
    .A3(_18842_),
    .ZN(_18843_));
 NAND3_X1 _24936_ (.A1(_18806_),
    .A2(_18841_),
    .A3(_18843_),
    .ZN(_18844_));
 NOR2_X1 _24937_ (.A1(_18697_),
    .A2(_18733_),
    .ZN(_18845_));
 OAI21_X2 _24938_ (.A(_18844_),
    .B1(_18845_),
    .B2(_18806_),
    .ZN(_18846_));
 OAI22_X4 _24939_ (.A1(_18666_),
    .A2(_18689_),
    .B1(_18846_),
    .B2(_18659_),
    .ZN(_18847_));
 NOR4_X4 _24940_ (.A1(_18787_),
    .A2(_18813_),
    .A3(_18839_),
    .A4(_18847_),
    .ZN(_18848_));
 AOI22_X2 _24941_ (.A1(\core.keymem.key_mem[14][16] ),
    .A2(_16439_),
    .B1(_16991_),
    .B2(\core.keymem.key_mem[6][16] ),
    .ZN(_18849_));
 AOI22_X2 _24942_ (.A1(\core.keymem.key_mem[4][16] ),
    .A2(_18232_),
    .B1(_17003_),
    .B2(\core.keymem.key_mem[1][16] ),
    .ZN(_18850_));
 AOI22_X2 _24943_ (.A1(\core.keymem.key_mem[7][16] ),
    .A2(_16408_),
    .B1(_17914_),
    .B2(\core.keymem.key_mem[9][16] ),
    .ZN(_18851_));
 AOI22_X2 _24944_ (.A1(\core.keymem.key_mem[2][16] ),
    .A2(_16994_),
    .B1(_17768_),
    .B2(\core.keymem.key_mem[11][16] ),
    .ZN(_18852_));
 NAND4_X2 _24945_ (.A1(_18849_),
    .A2(_18850_),
    .A3(_18851_),
    .A4(_18852_),
    .ZN(_18853_));
 AOI22_X1 _24946_ (.A1(\core.keymem.key_mem[3][16] ),
    .A2(_17683_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][16] ),
    .ZN(_18854_));
 AOI22_X2 _24947_ (.A1(\core.keymem.key_mem[8][16] ),
    .A2(_16453_),
    .B1(_17675_),
    .B2(\core.keymem.key_mem[5][16] ),
    .ZN(_18855_));
 AOI22_X2 _24948_ (.A1(\core.keymem.key_mem[10][16] ),
    .A2(_16433_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][16] ),
    .ZN(_18856_));
 NAND3_X2 _24949_ (.A1(_18854_),
    .A2(_18855_),
    .A3(_18856_),
    .ZN(_18857_));
 NOR3_X4 _24950_ (.A1(_17183_),
    .A2(_18853_),
    .A3(_18857_),
    .ZN(_18858_));
 AOI21_X4 _24951_ (.A(_18858_),
    .B1(_16498_),
    .B2(_00254_),
    .ZN(_18859_));
 XNOR2_X1 _24952_ (.A(\block_reg[3][16] ),
    .B(_18859_),
    .ZN(_18860_));
 AOI22_X1 _24953_ (.A1(\core.keymem.key_mem[4][112] ),
    .A2(_16946_),
    .B1(_16858_),
    .B2(\core.keymem.key_mem[2][112] ),
    .ZN(_18861_));
 AOI21_X1 _24954_ (.A(_16544_),
    .B1(_16461_),
    .B2(\core.keymem.key_mem[9][112] ),
    .ZN(_18862_));
 AOI22_X1 _24955_ (.A1(\core.keymem.key_mem[3][112] ),
    .A2(_16864_),
    .B1(_16431_),
    .B2(\core.keymem.key_mem[10][112] ),
    .ZN(_18863_));
 AOI22_X1 _24956_ (.A1(\core.keymem.key_mem[11][112] ),
    .A2(_16441_),
    .B1(_16471_),
    .B2(\core.keymem.key_mem[13][112] ),
    .ZN(_18864_));
 AND4_X1 _24957_ (.A1(_18861_),
    .A2(_18862_),
    .A3(_18863_),
    .A4(_18864_),
    .ZN(_18865_));
 AOI222_X2 _24958_ (.A1(\core.keymem.key_mem[14][112] ),
    .A2(_16436_),
    .B1(_16519_),
    .B2(\core.keymem.key_mem[6][112] ),
    .C1(_16466_),
    .C2(\core.keymem.key_mem[5][112] ),
    .ZN(_18866_));
 AOI22_X1 _24959_ (.A1(\core.keymem.key_mem[7][112] ),
    .A2(_16406_),
    .B1(_16397_),
    .B2(\core.keymem.key_mem[12][112] ),
    .ZN(_18867_));
 AOI22_X1 _24960_ (.A1(\core.keymem.key_mem[8][112] ),
    .A2(_16451_),
    .B1(_16415_),
    .B2(\core.keymem.key_mem[1][112] ),
    .ZN(_18868_));
 AND3_X1 _24961_ (.A1(_18866_),
    .A2(_18867_),
    .A3(_18868_),
    .ZN(_18869_));
 AOI22_X4 _24962_ (.A1(_00180_),
    .A2(_16871_),
    .B1(_18865_),
    .B2(_18869_),
    .ZN(_18870_));
 XNOR2_X2 _24963_ (.A(\core.dec_block.block_w0_reg[16] ),
    .B(_18870_),
    .ZN(_18871_));
 OAI221_X2 _24964_ (.A(_18329_),
    .B1(_18466_),
    .B2(_18860_),
    .C1(_18871_),
    .C2(_18479_),
    .ZN(_18872_));
 AOI222_X2 _24965_ (.A1(\core.keymem.key_mem[2][6] ),
    .A2(_16993_),
    .B1(_16528_),
    .B2(\core.keymem.key_mem[8][6] ),
    .C1(\core.keymem.key_mem[12][6] ),
    .C2(_16397_),
    .ZN(_18873_));
 AOI22_X2 _24966_ (.A1(\core.keymem.key_mem[4][6] ),
    .A2(_16947_),
    .B1(_17175_),
    .B2(\core.keymem.key_mem[3][6] ),
    .ZN(_18874_));
 AOI22_X2 _24967_ (.A1(\core.keymem.key_mem[11][6] ),
    .A2(_16442_),
    .B1(_16472_),
    .B2(\core.keymem.key_mem[13][6] ),
    .ZN(_18875_));
 NAND3_X2 _24968_ (.A1(_18873_),
    .A2(_18874_),
    .A3(_18875_),
    .ZN(_18876_));
 AOI22_X1 _24969_ (.A1(\core.keymem.key_mem[14][6] ),
    .A2(_16998_),
    .B1(_17736_),
    .B2(\core.keymem.key_mem[7][6] ),
    .ZN(_18877_));
 AOI22_X2 _24970_ (.A1(\core.keymem.key_mem[10][6] ),
    .A2(_16432_),
    .B1(_16524_),
    .B2(\core.keymem.key_mem[1][6] ),
    .ZN(_18878_));
 AOI22_X2 _24971_ (.A1(\core.keymem.key_mem[9][6] ),
    .A2(_17522_),
    .B1(_17004_),
    .B2(\core.keymem.key_mem[5][6] ),
    .ZN(_18879_));
 AOI21_X1 _24972_ (.A(_16494_),
    .B1(_16520_),
    .B2(\core.keymem.key_mem[6][6] ),
    .ZN(_18880_));
 NAND4_X2 _24973_ (.A1(_18877_),
    .A2(_18878_),
    .A3(_18879_),
    .A4(_18880_),
    .ZN(_18881_));
 NOR2_X4 _24974_ (.A1(_18876_),
    .A2(_18881_),
    .ZN(_18882_));
 AOI21_X4 _24975_ (.A(_18882_),
    .B1(_16852_),
    .B2(_00212_),
    .ZN(_18883_));
 XNOR2_X2 _24976_ (.A(\core.dec_block.block_w3_reg[6] ),
    .B(_18883_),
    .ZN(_18884_));
 NAND2_X1 _24977_ (.A1(_00211_),
    .A2(_16496_),
    .ZN(_18885_));
 AOI22_X2 _24978_ (.A1(\core.keymem.key_mem[7][5] ),
    .A2(_17084_),
    .B1(_16855_),
    .B2(\core.keymem.key_mem[1][5] ),
    .ZN(_18886_));
 AOI222_X2 _24979_ (.A1(\core.keymem.key_mem[6][5] ),
    .A2(_16448_),
    .B1(_17175_),
    .B2(\core.keymem.key_mem[3][5] ),
    .C1(_16988_),
    .C2(\core.keymem.key_mem[10][5] ),
    .ZN(_18887_));
 AOI22_X2 _24980_ (.A1(\core.keymem.key_mem[4][5] ),
    .A2(_16457_),
    .B1(_16529_),
    .B2(\core.keymem.key_mem[8][5] ),
    .ZN(_18888_));
 NAND3_X2 _24981_ (.A1(_18886_),
    .A2(_18887_),
    .A3(_18888_),
    .ZN(_18889_));
 AOI22_X1 _24982_ (.A1(\core.keymem.key_mem[12][5] ),
    .A2(_16398_),
    .B1(_16949_),
    .B2(\core.keymem.key_mem[5][5] ),
    .ZN(_18890_));
 AOI21_X1 _24983_ (.A(_16982_),
    .B1(_16860_),
    .B2(\core.keymem.key_mem[2][5] ),
    .ZN(_18891_));
 AOI22_X2 _24984_ (.A1(\core.keymem.key_mem[9][5] ),
    .A2(_16462_),
    .B1(_16472_),
    .B2(\core.keymem.key_mem[13][5] ),
    .ZN(_18892_));
 AOI22_X2 _24985_ (.A1(\core.keymem.key_mem[14][5] ),
    .A2(_16438_),
    .B1(_16442_),
    .B2(\core.keymem.key_mem[11][5] ),
    .ZN(_18893_));
 NAND4_X2 _24986_ (.A1(_18890_),
    .A2(_18891_),
    .A3(_18892_),
    .A4(_18893_),
    .ZN(_18894_));
 OAI21_X4 _24987_ (.A(_18885_),
    .B1(_18889_),
    .B2(_18894_),
    .ZN(_18895_));
 XOR2_X2 _24988_ (.A(\core.dec_block.block_w3_reg[5] ),
    .B(_18895_),
    .Z(_18896_));
 XNOR2_X2 _24989_ (.A(_18884_),
    .B(_18896_),
    .ZN(_18897_));
 AOI22_X2 _24990_ (.A1(\core.keymem.key_mem[2][21] ),
    .A2(_16859_),
    .B1(_16524_),
    .B2(\core.keymem.key_mem[1][21] ),
    .ZN(_18898_));
 AOI22_X2 _24991_ (.A1(\core.keymem.key_mem[9][21] ),
    .A2(_16535_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][21] ),
    .ZN(_18899_));
 AOI22_X2 _24992_ (.A1(\core.keymem.key_mem[8][21] ),
    .A2(_16528_),
    .B1(_16505_),
    .B2(\core.keymem.key_mem[11][21] ),
    .ZN(_18900_));
 AOI22_X2 _24993_ (.A1(\core.keymem.key_mem[7][21] ),
    .A2(_16955_),
    .B1(_17648_),
    .B2(\core.keymem.key_mem[6][21] ),
    .ZN(_18901_));
 NAND4_X2 _24994_ (.A1(_18898_),
    .A2(_18899_),
    .A3(_18900_),
    .A4(_18901_),
    .ZN(_18902_));
 AOI22_X1 _24995_ (.A1(\core.keymem.key_mem[4][21] ),
    .A2(_16499_),
    .B1(_16986_),
    .B2(\core.keymem.key_mem[3][21] ),
    .ZN(_18903_));
 AOI22_X2 _24996_ (.A1(\core.keymem.key_mem[5][21] ),
    .A2(_17004_),
    .B1(_17193_),
    .B2(\core.keymem.key_mem[13][21] ),
    .ZN(_18904_));
 AOI22_X2 _24997_ (.A1(\core.keymem.key_mem[14][21] ),
    .A2(_17191_),
    .B1(_16988_),
    .B2(\core.keymem.key_mem[10][21] ),
    .ZN(_18905_));
 NAND3_X2 _24998_ (.A1(_18903_),
    .A2(_18904_),
    .A3(_18905_),
    .ZN(_18906_));
 NOR3_X4 _24999_ (.A1(_16546_),
    .A2(_18902_),
    .A3(_18906_),
    .ZN(_18907_));
 AOI21_X4 _25000_ (.A(_18907_),
    .B1(_16852_),
    .B2(_00291_),
    .ZN(_18908_));
 XNOR2_X2 _25001_ (.A(\core.dec_block.block_w3_reg[21] ),
    .B(_18908_),
    .ZN(_18909_));
 NAND2_X2 _25002_ (.A1(_00292_),
    .A2(_16871_),
    .ZN(_18910_));
 AOI22_X1 _25003_ (.A1(\core.keymem.key_mem[4][22] ),
    .A2(_16455_),
    .B1(_16954_),
    .B2(\core.keymem.key_mem[7][22] ),
    .ZN(_18911_));
 AOI22_X1 _25004_ (.A1(\core.keymem.key_mem[6][22] ),
    .A2(_16519_),
    .B1(_16460_),
    .B2(\core.keymem.key_mem[9][22] ),
    .ZN(_18912_));
 AOI22_X1 _25005_ (.A1(\core.keymem.key_mem[8][22] ),
    .A2(_16450_),
    .B1(_16431_),
    .B2(\core.keymem.key_mem[10][22] ),
    .ZN(_18913_));
 AOI22_X1 _25006_ (.A1(\core.keymem.key_mem[1][22] ),
    .A2(_16523_),
    .B1(_16470_),
    .B2(\core.keymem.key_mem[13][22] ),
    .ZN(_18914_));
 AND4_X1 _25007_ (.A1(_18911_),
    .A2(_18912_),
    .A3(_18913_),
    .A4(_18914_),
    .ZN(_18915_));
 AOI22_X4 _25008_ (.A1(\core.keymem.key_mem[2][22] ),
    .A2(_16859_),
    .B1(_16505_),
    .B2(\core.keymem.key_mem[11][22] ),
    .ZN(_18916_));
 AOI22_X2 _25009_ (.A1(\core.keymem.key_mem[14][22] ),
    .A2(_17191_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][22] ),
    .ZN(_18917_));
 AOI22_X4 _25010_ (.A1(\core.keymem.key_mem[3][22] ),
    .A2(_16865_),
    .B1(_16467_),
    .B2(\core.keymem.key_mem[5][22] ),
    .ZN(_18918_));
 NAND4_X4 _25011_ (.A1(_18915_),
    .A2(_18916_),
    .A3(_18917_),
    .A4(_18918_),
    .ZN(_18919_));
 OAI21_X4 _25012_ (.A(_18910_),
    .B1(_18919_),
    .B2(_16871_),
    .ZN(_18920_));
 XOR2_X2 _25013_ (.A(\core.dec_block.block_w3_reg[22] ),
    .B(_18920_),
    .Z(_18921_));
 XNOR2_X2 _25014_ (.A(_18909_),
    .B(_18921_),
    .ZN(_18922_));
 XNOR2_X2 _25015_ (.A(_18897_),
    .B(_18922_),
    .ZN(_18923_));
 AOI22_X1 _25016_ (.A1(\core.keymem.key_mem[14][15] ),
    .A2(_17099_),
    .B1(_16902_),
    .B2(\core.keymem.key_mem[2][15] ),
    .ZN(_18924_));
 NOR2_X1 _25017_ (.A1(_16421_),
    .A2(_18924_),
    .ZN(_18925_));
 NAND3_X1 _25018_ (.A1(\core.keymem.key_mem[12][15] ),
    .A2(_16919_),
    .A3(_16931_),
    .ZN(_18926_));
 AOI22_X2 _25019_ (.A1(\core.keymem.key_mem[7][15] ),
    .A2(_16938_),
    .B1(_17025_),
    .B2(\core.keymem.key_mem[6][15] ),
    .ZN(_18927_));
 INV_X1 _25020_ (.A(\core.keymem.key_mem[13][15] ),
    .ZN(_18928_));
 OAI221_X2 _25021_ (.A(_18926_),
    .B1(_18927_),
    .B2(_17042_),
    .C1(_18928_),
    .C2(_17638_),
    .ZN(_18929_));
 OAI211_X2 _25022_ (.A(\core.keymem.key_mem[8][15] ),
    .B(_16921_),
    .C1(_16922_),
    .C2(_16923_),
    .ZN(_18930_));
 OAI211_X2 _25023_ (.A(\core.keymem.key_mem[4][15] ),
    .B(_16921_),
    .C1(_16933_),
    .C2(_16934_),
    .ZN(_18931_));
 OAI211_X2 _25024_ (.A(\core.keymem.key_mem[11][15] ),
    .B(_16938_),
    .C1(_16885_),
    .C2(_16889_),
    .ZN(_18932_));
 NAND3_X1 _25025_ (.A1(\core.keymem.key_mem[3][15] ),
    .A2(_16938_),
    .A3(_16969_),
    .ZN(_18933_));
 NAND4_X2 _25026_ (.A1(_18930_),
    .A2(_18931_),
    .A3(_18932_),
    .A4(_18933_),
    .ZN(_18934_));
 OAI221_X2 _25027_ (.A(\core.keymem.key_mem[9][15] ),
    .B1(_16926_),
    .B2(_16928_),
    .C1(_17018_),
    .C2(_17020_),
    .ZN(_18935_));
 OAI211_X2 _25028_ (.A(\core.keymem.key_mem[10][15] ),
    .B(_17015_),
    .C1(_16885_),
    .C2(_16889_),
    .ZN(_18936_));
 OAI211_X2 _25029_ (.A(\core.keymem.key_mem[1][15] ),
    .B(_16969_),
    .C1(_17018_),
    .C2(_17020_),
    .ZN(_18937_));
 OAI221_X2 _25030_ (.A(\core.keymem.key_mem[5][15] ),
    .B1(_16895_),
    .B2(_16898_),
    .C1(_17018_),
    .C2(_17020_),
    .ZN(_18938_));
 NAND4_X2 _25031_ (.A1(_18935_),
    .A2(_18936_),
    .A3(_18937_),
    .A4(_18938_),
    .ZN(_18939_));
 NOR4_X4 _25032_ (.A1(_18925_),
    .A2(_18929_),
    .A3(_18934_),
    .A4(_18939_),
    .ZN(_18940_));
 MUX2_X2 _25033_ (.A(_00253_),
    .B(_18940_),
    .S(_16487_),
    .Z(_18941_));
 XOR2_X2 _25034_ (.A(\core.dec_block.block_w3_reg[15] ),
    .B(_18941_),
    .Z(_18942_));
 AOI22_X1 _25035_ (.A1(\core.keymem.key_mem[9][23] ),
    .A2(_17914_),
    .B1(_17768_),
    .B2(\core.keymem.key_mem[11][23] ),
    .ZN(_18943_));
 AOI22_X1 _25036_ (.A1(\core.keymem.key_mem[4][23] ),
    .A2(_16500_),
    .B1(_17084_),
    .B2(\core.keymem.key_mem[7][23] ),
    .ZN(_18944_));
 AOI22_X1 _25037_ (.A1(\core.keymem.key_mem[3][23] ),
    .A2(_16987_),
    .B1(_17720_),
    .B2(\core.keymem.key_mem[12][23] ),
    .ZN(_18945_));
 AOI21_X1 _25038_ (.A(_17013_),
    .B1(_17675_),
    .B2(\core.keymem.key_mem[5][23] ),
    .ZN(_18946_));
 NAND4_X1 _25039_ (.A1(_18943_),
    .A2(_18944_),
    .A3(_18945_),
    .A4(_18946_),
    .ZN(_18947_));
 MUX2_X1 _25040_ (.A(\core.keymem.key_mem[6][23] ),
    .B(\core.keymem.key_mem[14][23] ),
    .S(_17054_),
    .Z(_18948_));
 AOI22_X1 _25041_ (.A1(\core.keymem.key_mem[10][23] ),
    .A2(_17067_),
    .B1(_17051_),
    .B2(_18948_),
    .ZN(_18949_));
 NOR2_X1 _25042_ (.A1(_16968_),
    .A2(_18949_),
    .ZN(_18950_));
 AOI22_X1 _25043_ (.A1(\core.keymem.key_mem[2][23] ),
    .A2(_16994_),
    .B1(_17781_),
    .B2(\core.keymem.key_mem[8][23] ),
    .ZN(_18951_));
 AOI22_X1 _25044_ (.A1(\core.keymem.key_mem[1][23] ),
    .A2(_17003_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][23] ),
    .ZN(_18952_));
 NAND2_X1 _25045_ (.A1(_18951_),
    .A2(_18952_),
    .ZN(_18953_));
 NOR3_X2 _25046_ (.A1(_18947_),
    .A2(_18950_),
    .A3(_18953_),
    .ZN(_18954_));
 AOI21_X4 _25047_ (.A(_18954_),
    .B1(_16548_),
    .B2(_00293_),
    .ZN(_18955_));
 XNOR2_X2 _25048_ (.A(_18576_),
    .B(_18955_),
    .ZN(_18956_));
 XNOR2_X2 _25049_ (.A(_18942_),
    .B(_18956_),
    .ZN(_18957_));
 XNOR2_X1 _25050_ (.A(_18923_),
    .B(_18957_),
    .ZN(_18958_));
 NAND2_X1 _25051_ (.A1(_00251_),
    .A2(_16984_),
    .ZN(_18959_));
 AOI22_X2 _25052_ (.A1(\core.keymem.key_mem[2][13] ),
    .A2(_16424_),
    .B1(_17175_),
    .B2(\core.keymem.key_mem[3][13] ),
    .ZN(_18960_));
 AOI22_X1 _25053_ (.A1(\core.keymem.key_mem[4][13] ),
    .A2(_16947_),
    .B1(_16520_),
    .B2(\core.keymem.key_mem[6][13] ),
    .ZN(_18961_));
 AOI22_X1 _25054_ (.A1(\core.keymem.key_mem[7][13] ),
    .A2(_16407_),
    .B1(_17506_),
    .B2(\core.keymem.key_mem[8][13] ),
    .ZN(_18962_));
 AOI22_X1 _25055_ (.A1(\core.keymem.key_mem[5][13] ),
    .A2(_16949_),
    .B1(_16472_),
    .B2(\core.keymem.key_mem[13][13] ),
    .ZN(_18963_));
 AND4_X1 _25056_ (.A1(_18960_),
    .A2(_18961_),
    .A3(_18962_),
    .A4(_18963_),
    .ZN(_18964_));
 AOI22_X2 _25057_ (.A1(\core.keymem.key_mem[14][13] ),
    .A2(_16439_),
    .B1(_16417_),
    .B2(\core.keymem.key_mem[1][13] ),
    .ZN(_18965_));
 AOI22_X2 _25058_ (.A1(\core.keymem.key_mem[9][13] ),
    .A2(_16463_),
    .B1(_16443_),
    .B2(\core.keymem.key_mem[11][13] ),
    .ZN(_18966_));
 AOI22_X4 _25059_ (.A1(\core.keymem.key_mem[10][13] ),
    .A2(_16433_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][13] ),
    .ZN(_18967_));
 NAND4_X4 _25060_ (.A1(_18964_),
    .A2(_18965_),
    .A3(_18966_),
    .A4(_18967_),
    .ZN(_18968_));
 OAI21_X4 _25061_ (.A(_18959_),
    .B1(_18968_),
    .B2(_16497_),
    .ZN(_18969_));
 XOR2_X2 _25062_ (.A(\core.dec_block.block_w3_reg[13] ),
    .B(_18969_),
    .Z(_18970_));
 NAND2_X1 _25063_ (.A1(_00294_),
    .A2(_16873_),
    .ZN(_18971_));
 AOI222_X2 _25064_ (.A1(\core.keymem.key_mem[6][24] ),
    .A2(_16449_),
    .B1(_16537_),
    .B2(\core.keymem.key_mem[9][24] ),
    .C1(\core.keymem.key_mem[11][24] ),
    .C2(_17768_),
    .ZN(_18972_));
 AOI22_X2 _25065_ (.A1(\core.keymem.key_mem[3][24] ),
    .A2(_17091_),
    .B1(_16516_),
    .B2(\core.keymem.key_mem[10][24] ),
    .ZN(_18973_));
 AOI22_X2 _25066_ (.A1(\core.keymem.key_mem[7][24] ),
    .A2(_17085_),
    .B1(_16540_),
    .B2(\core.keymem.key_mem[12][24] ),
    .ZN(_18974_));
 NAND3_X2 _25067_ (.A1(_18972_),
    .A2(_18973_),
    .A3(_18974_),
    .ZN(_18975_));
 AOI21_X2 _25068_ (.A(_16496_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][24] ),
    .ZN(_18976_));
 AOI22_X2 _25069_ (.A1(\core.keymem.key_mem[5][24] ),
    .A2(_16510_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][24] ),
    .ZN(_18977_));
 AOI22_X2 _25070_ (.A1(\core.keymem.key_mem[14][24] ),
    .A2(_16502_),
    .B1(_16453_),
    .B2(\core.keymem.key_mem[8][24] ),
    .ZN(_18978_));
 AOI22_X2 _25071_ (.A1(\core.keymem.key_mem[4][24] ),
    .A2(_16458_),
    .B1(_16425_),
    .B2(\core.keymem.key_mem[2][24] ),
    .ZN(_18979_));
 NAND4_X2 _25072_ (.A1(_18976_),
    .A2(_18977_),
    .A3(_18978_),
    .A4(_18979_),
    .ZN(_18980_));
 OAI21_X4 _25073_ (.A(_18971_),
    .B1(_18975_),
    .B2(_18980_),
    .ZN(_18981_));
 XOR2_X2 _25074_ (.A(\core.dec_block.block_w3_reg[24] ),
    .B(_18981_),
    .Z(_18982_));
 MUX2_X1 _25075_ (.A(\core.keymem.key_mem[9][29] ),
    .B(\core.keymem.key_mem[13][29] ),
    .S(_16960_),
    .Z(_18983_));
 NAND3_X1 _25076_ (.A1(_16964_),
    .A2(_17054_),
    .A3(_18983_),
    .ZN(_18984_));
 NOR2_X2 _25077_ (.A1(_16421_),
    .A2(_17054_),
    .ZN(_18985_));
 MUX2_X1 _25078_ (.A(\core.keymem.key_mem[2][29] ),
    .B(\core.keymem.key_mem[6][29] ),
    .S(_16961_),
    .Z(_18986_));
 NAND2_X1 _25079_ (.A1(_18985_),
    .A2(_18986_),
    .ZN(_18987_));
 AOI22_X2 _25080_ (.A1(\core.keymem.key_mem[14][29] ),
    .A2(_16437_),
    .B1(_16948_),
    .B2(\core.keymem.key_mem[5][29] ),
    .ZN(_18988_));
 NAND3_X2 _25081_ (.A1(_18984_),
    .A2(_18987_),
    .A3(_18988_),
    .ZN(_18989_));
 AOI22_X1 _25082_ (.A1(\core.keymem.key_mem[4][29] ),
    .A2(_17513_),
    .B1(_17067_),
    .B2(\core.keymem.key_mem[8][29] ),
    .ZN(_18990_));
 NOR2_X1 _25083_ (.A1(_16394_),
    .A2(_18990_),
    .ZN(_18991_));
 AOI221_X2 _25084_ (.A(_16383_),
    .B1(_16963_),
    .B2(\core.keymem.key_mem[1][29] ),
    .C1(_16480_),
    .C2(\core.keymem.key_mem[3][29] ),
    .ZN(_18992_));
 NAND3_X1 _25085_ (.A1(\core.keymem.key_mem[10][29] ),
    .A2(_16907_),
    .A3(_17043_),
    .ZN(_18993_));
 AOI21_X1 _25086_ (.A(_16958_),
    .B1(_16481_),
    .B2(\core.keymem.key_mem[7][29] ),
    .ZN(_18994_));
 OR2_X1 _25087_ (.A1(_16972_),
    .A2(_18994_),
    .ZN(_18995_));
 AOI21_X2 _25088_ (.A(_18992_),
    .B1(_18993_),
    .B2(_18995_),
    .ZN(_18996_));
 NAND3_X1 _25089_ (.A1(\core.keymem.key_mem[11][29] ),
    .A2(_16901_),
    .A3(_16958_),
    .ZN(_18997_));
 NAND3_X1 _25090_ (.A1(\core.keymem.key_mem[12][29] ),
    .A2(_16931_),
    .A3(_16961_),
    .ZN(_18998_));
 AOI21_X2 _25091_ (.A(_16967_),
    .B1(_18997_),
    .B2(_18998_),
    .ZN(_18999_));
 NOR4_X4 _25092_ (.A1(_18989_),
    .A2(_18991_),
    .A3(_18996_),
    .A4(_18999_),
    .ZN(_19000_));
 MUX2_X2 _25093_ (.A(_00295_),
    .B(_19000_),
    .S(_16487_),
    .Z(_19001_));
 XOR2_X2 _25094_ (.A(\core.dec_block.block_w3_reg[29] ),
    .B(_19001_),
    .Z(_19002_));
 XNOR2_X2 _25095_ (.A(_18982_),
    .B(_19002_),
    .ZN(_19003_));
 XNOR2_X2 _25096_ (.A(_18970_),
    .B(_19003_),
    .ZN(_19004_));
 AOI222_X2 _25097_ (.A1(\core.keymem.key_mem[12][8] ),
    .A2(_16540_),
    .B1(_16469_),
    .B2(\core.keymem.key_mem[5][8] ),
    .C1(\core.keymem.key_mem[4][8] ),
    .C2(_18232_),
    .ZN(_19005_));
 AOI22_X1 _25098_ (.A1(\core.keymem.key_mem[9][8] ),
    .A2(_17585_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][8] ),
    .ZN(_19006_));
 AOI22_X1 _25099_ (.A1(\core.keymem.key_mem[2][8] ),
    .A2(_16425_),
    .B1(_16507_),
    .B2(\core.keymem.key_mem[11][8] ),
    .ZN(_19007_));
 NAND3_X1 _25100_ (.A1(_19005_),
    .A2(_19006_),
    .A3(_19007_),
    .ZN(_19008_));
 AOI22_X1 _25101_ (.A1(\core.keymem.key_mem[6][8] ),
    .A2(_16522_),
    .B1(_16387_),
    .B2(\core.keymem.key_mem[3][8] ),
    .ZN(_19009_));
 AOI22_X1 _25102_ (.A1(\core.keymem.key_mem[7][8] ),
    .A2(_17085_),
    .B1(_16530_),
    .B2(\core.keymem.key_mem[8][8] ),
    .ZN(_19010_));
 AOI22_X1 _25103_ (.A1(\core.keymem.key_mem[14][8] ),
    .A2(_16502_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][8] ),
    .ZN(_19011_));
 AOI21_X1 _25104_ (.A(_17014_),
    .B1(_16516_),
    .B2(\core.keymem.key_mem[10][8] ),
    .ZN(_19012_));
 NAND4_X1 _25105_ (.A1(_19009_),
    .A2(_19010_),
    .A3(_19011_),
    .A4(_19012_),
    .ZN(_19013_));
 NOR2_X2 _25106_ (.A1(_19008_),
    .A2(_19013_),
    .ZN(_19014_));
 AOI21_X4 _25107_ (.A(_19014_),
    .B1(_16549_),
    .B2(_00214_),
    .ZN(_19015_));
 XNOR2_X2 _25108_ (.A(\core.dec_block.block_w3_reg[8] ),
    .B(_19015_),
    .ZN(_19016_));
 AOI22_X1 _25109_ (.A1(\core.keymem.key_mem[6][0] ),
    .A2(_16447_),
    .B1(_16397_),
    .B2(\core.keymem.key_mem[12][0] ),
    .ZN(_19017_));
 AOI21_X1 _25110_ (.A(_16544_),
    .B1(_16451_),
    .B2(\core.keymem.key_mem[8][0] ),
    .ZN(_19018_));
 AOI22_X1 _25111_ (.A1(\core.keymem.key_mem[14][0] ),
    .A2(_16437_),
    .B1(_16441_),
    .B2(\core.keymem.key_mem[11][0] ),
    .ZN(_19019_));
 AOI22_X1 _25112_ (.A1(\core.keymem.key_mem[7][0] ),
    .A2(_16406_),
    .B1(_16471_),
    .B2(\core.keymem.key_mem[13][0] ),
    .ZN(_19020_));
 AND4_X1 _25113_ (.A1(_19017_),
    .A2(_19018_),
    .A3(_19019_),
    .A4(_19020_),
    .ZN(_19021_));
 AOI222_X2 _25114_ (.A1(\core.keymem.key_mem[4][0] ),
    .A2(_16946_),
    .B1(_16858_),
    .B2(\core.keymem.key_mem[2][0] ),
    .C1(_16466_),
    .C2(\core.keymem.key_mem[5][0] ),
    .ZN(_19022_));
 AOI22_X1 _25115_ (.A1(\core.keymem.key_mem[10][0] ),
    .A2(_16514_),
    .B1(_16415_),
    .B2(\core.keymem.key_mem[1][0] ),
    .ZN(_19023_));
 AOI22_X1 _25116_ (.A1(\core.keymem.key_mem[3][0] ),
    .A2(_16385_),
    .B1(_16461_),
    .B2(\core.keymem.key_mem[9][0] ),
    .ZN(_19024_));
 AND3_X1 _25117_ (.A1(_19022_),
    .A2(_19023_),
    .A3(_19024_),
    .ZN(_19025_));
 AOI22_X4 _25118_ (.A1(_00173_),
    .A2(_16546_),
    .B1(_19021_),
    .B2(_19025_),
    .ZN(_19026_));
 XNOR2_X2 _25119_ (.A(\core.dec_block.block_w3_reg[0] ),
    .B(_19026_),
    .ZN(_19027_));
 XOR2_X1 _25120_ (.A(_19016_),
    .B(_19027_),
    .Z(_19028_));
 XNOR2_X1 _25121_ (.A(_19004_),
    .B(_19028_),
    .ZN(_19029_));
 XNOR2_X1 _25122_ (.A(_18958_),
    .B(_19029_),
    .ZN(_19030_));
 BUF_X4 _25123_ (.A(_17748_),
    .Z(_19031_));
 AOI21_X1 _25124_ (.A(_18872_),
    .B1(_19030_),
    .B2(_19031_),
    .ZN(_19032_));
 AOI21_X1 _25125_ (.A(_18565_),
    .B1(_18848_),
    .B2(_19032_),
    .ZN(_00574_));
 INV_X1 _25126_ (.A(\core.dec_block.block_w0_reg[17] ),
    .ZN(_19033_));
 BUF_X4 _25127_ (.A(_18573_),
    .Z(_19034_));
 NOR2_X1 _25128_ (.A1(_19034_),
    .A2(_18743_),
    .ZN(_19035_));
 NOR3_X1 _25129_ (.A1(_18763_),
    .A2(_18609_),
    .A3(_18721_),
    .ZN(_19036_));
 OAI21_X1 _25130_ (.A(_18788_),
    .B1(_19035_),
    .B2(_19036_),
    .ZN(_19037_));
 NAND3_X1 _25131_ (.A1(_18715_),
    .A2(_18662_),
    .A3(_18719_),
    .ZN(_19038_));
 AOI21_X1 _25132_ (.A(_18842_),
    .B1(_18783_),
    .B2(_18816_),
    .ZN(_19039_));
 BUF_X4 _25133_ (.A(_18670_),
    .Z(_19040_));
 OAI221_X2 _25134_ (.A(_19037_),
    .B1(_19038_),
    .B2(_18788_),
    .C1(_19039_),
    .C2(_19040_),
    .ZN(_19041_));
 AOI21_X1 _25135_ (.A(_18670_),
    .B1(_18721_),
    .B2(_18665_),
    .ZN(_19042_));
 AOI221_X2 _25136_ (.A(_19042_),
    .B1(_18726_),
    .B2(_18774_),
    .C1(_18702_),
    .C2(_18802_),
    .ZN(_19043_));
 OAI21_X1 _25137_ (.A(_18619_),
    .B1(_18596_),
    .B2(_18755_),
    .ZN(_19044_));
 NAND2_X2 _25138_ (.A1(_18596_),
    .A2(_18633_),
    .ZN(_19045_));
 NAND3_X1 _25139_ (.A1(_18645_),
    .A2(_19044_),
    .A3(_19045_),
    .ZN(_19046_));
 MUX2_X1 _25140_ (.A(_18585_),
    .B(_18752_),
    .S(_18619_),
    .Z(_19047_));
 AOI21_X1 _25141_ (.A(_19046_),
    .B1(_19047_),
    .B2(_18626_),
    .ZN(_19048_));
 OAI22_X2 _25142_ (.A1(_18633_),
    .A2(_18684_),
    .B1(_19045_),
    .B2(_18629_),
    .ZN(_19049_));
 NOR3_X1 _25143_ (.A1(_18645_),
    .A2(_18745_),
    .A3(_18725_),
    .ZN(_19050_));
 AOI221_X2 _25144_ (.A(_19048_),
    .B1(_19049_),
    .B2(_19050_),
    .C1(_18636_),
    .C2(_18620_),
    .ZN(_19051_));
 BUF_X4 _25145_ (.A(_18773_),
    .Z(_19052_));
 NOR2_X2 _25146_ (.A1(_19052_),
    .A2(_18681_),
    .ZN(_19053_));
 AOI22_X2 _25147_ (.A1(_18708_),
    .A2(_18740_),
    .B1(_19053_),
    .B2(_18779_),
    .ZN(_19054_));
 NAND3_X1 _25148_ (.A1(_18642_),
    .A2(_18633_),
    .A3(_18688_),
    .ZN(_19055_));
 AOI21_X1 _25149_ (.A(_19055_),
    .B1(_18581_),
    .B2(_18750_),
    .ZN(_19056_));
 OAI21_X1 _25150_ (.A(_18814_),
    .B1(_18695_),
    .B2(_18755_),
    .ZN(_19057_));
 AOI22_X1 _25151_ (.A1(_18624_),
    .A2(_18629_),
    .B1(_18645_),
    .B2(_18573_),
    .ZN(_19058_));
 OAI21_X1 _25152_ (.A(_19057_),
    .B1(_19058_),
    .B2(_18633_),
    .ZN(_19059_));
 AOI221_X1 _25153_ (.A(_19056_),
    .B1(_19059_),
    .B2(_18750_),
    .C1(_18662_),
    .C2(_18761_),
    .ZN(_19060_));
 NAND4_X1 _25154_ (.A1(_19043_),
    .A2(_19051_),
    .A3(_19054_),
    .A4(_19060_),
    .ZN(_19061_));
 NOR3_X1 _25155_ (.A1(_18629_),
    .A2(_18581_),
    .A3(_19045_),
    .ZN(_19062_));
 AOI21_X1 _25156_ (.A(_19062_),
    .B1(_18650_),
    .B2(_18631_),
    .ZN(_19063_));
 NOR2_X1 _25157_ (.A1(_18658_),
    .A2(_19063_),
    .ZN(_19064_));
 AOI21_X1 _25158_ (.A(_18634_),
    .B1(_18695_),
    .B2(_18750_),
    .ZN(_19065_));
 NOR3_X1 _25159_ (.A1(_18621_),
    .A2(_18629_),
    .A3(_19065_),
    .ZN(_19066_));
 OAI21_X1 _25160_ (.A(_18805_),
    .B1(_19064_),
    .B2(_19066_),
    .ZN(_19067_));
 OAI21_X1 _25161_ (.A(_18746_),
    .B1(_18707_),
    .B2(_18779_),
    .ZN(_19068_));
 AOI22_X2 _25162_ (.A1(_18670_),
    .A2(_18705_),
    .B1(_18801_),
    .B2(_19068_),
    .ZN(_19069_));
 NOR2_X2 _25163_ (.A1(_18674_),
    .A2(_18675_),
    .ZN(_19070_));
 NOR2_X4 _25164_ (.A1(_18679_),
    .A2(_18706_),
    .ZN(_19071_));
 NOR2_X1 _25165_ (.A1(_18639_),
    .A2(_18728_),
    .ZN(_19072_));
 AOI221_X2 _25166_ (.A(_19069_),
    .B1(_19070_),
    .B2(_18765_),
    .C1(_19071_),
    .C2(_19072_),
    .ZN(_19073_));
 AOI21_X1 _25167_ (.A(_18639_),
    .B1(_18727_),
    .B2(_18666_),
    .ZN(_19074_));
 NOR2_X1 _25168_ (.A1(_18621_),
    .A2(_18717_),
    .ZN(_19075_));
 NAND2_X1 _25169_ (.A1(_19034_),
    .A2(_18779_),
    .ZN(_19076_));
 OAI21_X1 _25170_ (.A(_19076_),
    .B1(_18766_),
    .B2(_18736_),
    .ZN(_19077_));
 AOI21_X2 _25171_ (.A(_19074_),
    .B1(_19075_),
    .B2(_19077_),
    .ZN(_19078_));
 NAND3_X1 _25172_ (.A1(_19067_),
    .A2(_19073_),
    .A3(_19078_),
    .ZN(_19079_));
 NOR3_X1 _25173_ (.A1(_19041_),
    .A2(_19061_),
    .A3(_19079_),
    .ZN(_19080_));
 NOR2_X2 _25174_ (.A1(_18675_),
    .A2(_19052_),
    .ZN(_19081_));
 NOR2_X2 _25175_ (.A1(_18676_),
    .A2(_18639_),
    .ZN(_19082_));
 OAI21_X1 _25176_ (.A(_18778_),
    .B1(_19081_),
    .B2(_19082_),
    .ZN(_19083_));
 NOR2_X1 _25177_ (.A1(_18623_),
    .A2(_18651_),
    .ZN(_19084_));
 NOR2_X1 _25178_ (.A1(_18842_),
    .A2(_19084_),
    .ZN(_19085_));
 OAI221_X2 _25179_ (.A(_19083_),
    .B1(_18733_),
    .B2(_18729_),
    .C1(_19052_),
    .C2(_19085_),
    .ZN(_19086_));
 OAI22_X1 _25180_ (.A1(_18796_),
    .A2(_18651_),
    .B1(_18736_),
    .B2(_18819_),
    .ZN(_19087_));
 NAND2_X1 _25181_ (.A1(_18796_),
    .A2(_18765_),
    .ZN(_19088_));
 NAND2_X1 _25182_ (.A1(_18810_),
    .A2(_19088_),
    .ZN(_19089_));
 AOI221_X2 _25183_ (.A(_19086_),
    .B1(_19087_),
    .B2(_18703_),
    .C1(_18815_),
    .C2(_19089_),
    .ZN(_19090_));
 OAI21_X1 _25184_ (.A(_19034_),
    .B1(_18765_),
    .B2(_19084_),
    .ZN(_19091_));
 AOI21_X1 _25185_ (.A(_18658_),
    .B1(_18696_),
    .B2(_19091_),
    .ZN(_19092_));
 NAND2_X1 _25186_ (.A1(_18695_),
    .A2(_18597_),
    .ZN(_19093_));
 BUF_X4 _25187_ (.A(_19093_),
    .Z(_19094_));
 NOR3_X1 _25188_ (.A1(_18620_),
    .A2(_18697_),
    .A3(_19094_),
    .ZN(_19095_));
 AOI21_X1 _25189_ (.A(_19095_),
    .B1(_18712_),
    .B2(_18620_),
    .ZN(_19096_));
 OAI22_X2 _25190_ (.A1(_19052_),
    .A2(_18801_),
    .B1(_19096_),
    .B2(_19034_),
    .ZN(_19097_));
 NOR2_X2 _25191_ (.A1(_18675_),
    .A2(_18801_),
    .ZN(_19098_));
 AOI21_X1 _25192_ (.A(_19098_),
    .B1(_18726_),
    .B2(_18738_),
    .ZN(_19099_));
 OAI22_X2 _25193_ (.A1(_19040_),
    .A2(_19088_),
    .B1(_19099_),
    .B2(_18763_),
    .ZN(_19100_));
 AOI221_X2 _25194_ (.A(_19092_),
    .B1(_19097_),
    .B2(_18654_),
    .C1(_18699_),
    .C2(_19100_),
    .ZN(_19101_));
 NAND4_X2 _25195_ (.A1(_18838_),
    .A2(_19080_),
    .A3(_19090_),
    .A4(_19101_),
    .ZN(_19102_));
 OAI21_X1 _25196_ (.A(_18647_),
    .B1(_18677_),
    .B2(_18740_),
    .ZN(_19103_));
 NOR2_X4 _25197_ (.A1(_18642_),
    .A2(_18635_),
    .ZN(_19104_));
 NAND2_X1 _25198_ (.A1(_19104_),
    .A2(_19053_),
    .ZN(_19105_));
 AOI222_X2 _25199_ (.A1(_18662_),
    .A2(_18682_),
    .B1(_18774_),
    .B2(_18783_),
    .C1(_18677_),
    .C2(_18780_),
    .ZN(_19106_));
 NAND4_X4 _25200_ (.A1(_19102_),
    .A2(_19103_),
    .A3(_19105_),
    .A4(_19106_),
    .ZN(_19107_));
 NAND2_X1 _25201_ (.A1(_18717_),
    .A2(_19104_),
    .ZN(_19108_));
 OAI21_X1 _25202_ (.A(_18807_),
    .B1(_18780_),
    .B2(_19098_),
    .ZN(_19109_));
 AOI21_X1 _25203_ (.A(_18640_),
    .B1(_19108_),
    .B2(_19109_),
    .ZN(_19110_));
 NOR2_X1 _25204_ (.A1(_18639_),
    .A2(_18721_),
    .ZN(_19111_));
 AOI21_X1 _25205_ (.A(_18768_),
    .B1(_19111_),
    .B2(_18823_),
    .ZN(_19112_));
 NAND2_X1 _25206_ (.A1(_18815_),
    .A2(_18653_),
    .ZN(_19113_));
 AOI21_X1 _25207_ (.A(_19112_),
    .B1(_19113_),
    .B2(_18640_),
    .ZN(_19114_));
 NAND2_X1 _25208_ (.A1(_18750_),
    .A2(_18634_),
    .ZN(_19115_));
 NOR3_X1 _25209_ (.A1(_18741_),
    .A2(_18676_),
    .A3(_19115_),
    .ZN(_19116_));
 XNOR2_X1 _25210_ (.A(_18645_),
    .B(_18648_),
    .ZN(_19117_));
 NAND4_X1 _25211_ (.A1(_18631_),
    .A2(_18633_),
    .A3(_18654_),
    .A4(_19117_),
    .ZN(_19118_));
 OAI21_X1 _25212_ (.A(_19118_),
    .B1(_19115_),
    .B2(_18807_),
    .ZN(_19119_));
 AOI21_X1 _25213_ (.A(_19116_),
    .B1(_19119_),
    .B2(_18741_),
    .ZN(_19120_));
 OAI21_X1 _25214_ (.A(_19073_),
    .B1(_19120_),
    .B2(_19052_),
    .ZN(_19121_));
 NAND2_X1 _25215_ (.A1(_18698_),
    .A2(_18711_),
    .ZN(_19122_));
 NOR3_X1 _25216_ (.A1(_18788_),
    .A2(_18654_),
    .A3(_19122_),
    .ZN(_19123_));
 NAND2_X1 _25217_ (.A1(_18711_),
    .A2(_18609_),
    .ZN(_19124_));
 AOI21_X1 _25218_ (.A(_18658_),
    .B1(_18693_),
    .B2(_19124_),
    .ZN(_19125_));
 OAI21_X1 _25219_ (.A(_18716_),
    .B1(_19123_),
    .B2(_19125_),
    .ZN(_19126_));
 AOI21_X1 _25220_ (.A(_18774_),
    .B1(_18753_),
    .B2(_18707_),
    .ZN(_19127_));
 AOI21_X1 _25221_ (.A(_19127_),
    .B1(_18733_),
    .B2(_18651_),
    .ZN(_19128_));
 NAND2_X1 _25222_ (.A1(_18694_),
    .A2(_18676_),
    .ZN(_19129_));
 OAI22_X2 _25223_ (.A1(_18718_),
    .A2(_18733_),
    .B1(_19094_),
    .B2(_19129_),
    .ZN(_19130_));
 NAND2_X1 _25224_ (.A1(_18624_),
    .A2(_18623_),
    .ZN(_19131_));
 NOR2_X1 _25225_ (.A1(_19034_),
    .A2(_19131_),
    .ZN(_19132_));
 AOI221_X2 _25226_ (.A(_19128_),
    .B1(_19130_),
    .B2(_18746_),
    .C1(_19132_),
    .C2(_18818_),
    .ZN(_19133_));
 NAND2_X4 _25227_ (.A1(_18629_),
    .A2(_18691_),
    .ZN(_19134_));
 NAND2_X4 _25228_ (.A1(_18613_),
    .A2(_18702_),
    .ZN(_19135_));
 NAND2_X2 _25229_ (.A1(_18648_),
    .A2(_18628_),
    .ZN(_19136_));
 OAI22_X1 _25230_ (.A1(_19134_),
    .A2(_19135_),
    .B1(_19136_),
    .B2(_18722_),
    .ZN(_19137_));
 AOI21_X1 _25231_ (.A(_19137_),
    .B1(_18740_),
    .B2(_18686_),
    .ZN(_19138_));
 NAND2_X2 _25232_ (.A1(_18815_),
    .A2(_18717_),
    .ZN(_19139_));
 NOR2_X1 _25233_ (.A1(_18647_),
    .A2(_18685_),
    .ZN(_19140_));
 AOI21_X1 _25234_ (.A(_19139_),
    .B1(_19140_),
    .B2(_18696_),
    .ZN(_19141_));
 NOR2_X2 _25235_ (.A1(_18674_),
    .A2(_18697_),
    .ZN(_19142_));
 AOI22_X1 _25236_ (.A1(_18779_),
    .A2(_19081_),
    .B1(_19142_),
    .B2(_18662_),
    .ZN(_19143_));
 NAND2_X2 _25237_ (.A1(_18688_),
    .A2(_18717_),
    .ZN(_19144_));
 OAI21_X1 _25238_ (.A(_19143_),
    .B1(_19144_),
    .B2(_19094_),
    .ZN(_19145_));
 NOR2_X1 _25239_ (.A1(_19141_),
    .A2(_19145_),
    .ZN(_19146_));
 NAND4_X1 _25240_ (.A1(_19126_),
    .A2(_19133_),
    .A3(_19138_),
    .A4(_19146_),
    .ZN(_19147_));
 NOR4_X2 _25241_ (.A1(_19110_),
    .A2(_19114_),
    .A3(_19121_),
    .A4(_19147_),
    .ZN(_19148_));
 OAI33_X1 _25242_ (.A1(_18782_),
    .A2(_18717_),
    .A3(_18722_),
    .B1(_18725_),
    .B2(_18801_),
    .B3(_18816_),
    .ZN(_19149_));
 NAND2_X2 _25243_ (.A1(_18746_),
    .A2(_18717_),
    .ZN(_19150_));
 AOI21_X1 _25244_ (.A(_19134_),
    .B1(_19113_),
    .B2(_19150_),
    .ZN(_19151_));
 AOI221_X2 _25245_ (.A(_19151_),
    .B1(_18680_),
    .B2(_18628_),
    .C1(_18815_),
    .C2(_18783_),
    .ZN(_19152_));
 AOI22_X2 _25246_ (.A1(_18686_),
    .A2(_18668_),
    .B1(_18842_),
    .B2(_18736_),
    .ZN(_19153_));
 NOR3_X1 _25247_ (.A1(_18805_),
    .A2(_18609_),
    .A3(_18696_),
    .ZN(_19154_));
 NOR2_X1 _25248_ (.A1(_18808_),
    .A2(_18693_),
    .ZN(_19155_));
 AOI21_X1 _25249_ (.A(_19154_),
    .B1(_19155_),
    .B2(_18806_),
    .ZN(_19156_));
 OAI221_X2 _25250_ (.A(_19152_),
    .B1(_19153_),
    .B2(_19040_),
    .C1(_19156_),
    .C2(_18659_),
    .ZN(_19157_));
 NOR2_X2 _25251_ (.A1(_19149_),
    .A2(_19157_),
    .ZN(_19158_));
 OAI22_X1 _25252_ (.A1(_18816_),
    .A2(_18744_),
    .B1(_18668_),
    .B2(_18810_),
    .ZN(_19159_));
 AOI22_X2 _25253_ (.A1(_18708_),
    .A2(_18677_),
    .B1(_19159_),
    .B2(_18703_),
    .ZN(_19160_));
 NOR3_X1 _25254_ (.A1(_18819_),
    .A2(_18670_),
    .A3(_18719_),
    .ZN(_19161_));
 AOI221_X2 _25255_ (.A(_19161_),
    .B1(_18740_),
    .B2(_18778_),
    .C1(_18708_),
    .C2(_19082_),
    .ZN(_19162_));
 NAND2_X1 _25256_ (.A1(_18780_),
    .A2(_19070_),
    .ZN(_19163_));
 NAND2_X2 _25257_ (.A1(_18815_),
    .A2(_18668_),
    .ZN(_19164_));
 AOI21_X1 _25258_ (.A(_18810_),
    .B1(_19164_),
    .B2(_18689_),
    .ZN(_19165_));
 AOI221_X2 _25259_ (.A(_19165_),
    .B1(_19071_),
    .B2(_18677_),
    .C1(_18647_),
    .C2(_18628_),
    .ZN(_19166_));
 NAND4_X2 _25260_ (.A1(_19160_),
    .A2(_19162_),
    .A3(_19163_),
    .A4(_19166_),
    .ZN(_19167_));
 NAND2_X2 _25261_ (.A1(_18664_),
    .A2(_18650_),
    .ZN(_19168_));
 OAI21_X1 _25262_ (.A(_18670_),
    .B1(_18639_),
    .B2(_18648_),
    .ZN(_19169_));
 AOI221_X1 _25263_ (.A(_18761_),
    .B1(_19169_),
    .B2(_18796_),
    .C1(_18698_),
    .C2(_18746_),
    .ZN(_19170_));
 NOR2_X1 _25264_ (.A1(_19168_),
    .A2(_19170_),
    .ZN(_19171_));
 NAND2_X1 _25265_ (.A1(_18702_),
    .A2(_18778_),
    .ZN(_19172_));
 NAND3_X1 _25266_ (.A1(_18815_),
    .A2(_18808_),
    .A3(_18768_),
    .ZN(_19173_));
 AOI21_X1 _25267_ (.A(_18807_),
    .B1(_19172_),
    .B2(_19173_),
    .ZN(_19174_));
 NAND2_X1 _25268_ (.A1(_18686_),
    .A2(_18753_),
    .ZN(_19175_));
 OAI221_X2 _25269_ (.A(_19175_),
    .B1(_19134_),
    .B2(_18775_),
    .C1(_18693_),
    .C2(_19144_),
    .ZN(_19176_));
 NOR4_X2 _25270_ (.A1(_19167_),
    .A2(_19171_),
    .A3(_19174_),
    .A4(_19176_),
    .ZN(_19177_));
 NAND4_X2 _25271_ (.A1(_18669_),
    .A2(_19148_),
    .A3(_19158_),
    .A4(_19177_),
    .ZN(_19178_));
 OAI21_X2 _25272_ (.A(_18416_),
    .B1(_19107_),
    .B2(_19178_),
    .ZN(_19179_));
 BUF_X4 _25273_ (.A(_16554_),
    .Z(_19180_));
 NAND2_X1 _25274_ (.A1(_00191_),
    .A2(_17578_),
    .ZN(_19181_));
 AOI22_X1 _25275_ (.A1(\core.keymem.key_mem[10][113] ),
    .A2(_16516_),
    .B1(_17178_),
    .B2(\core.keymem.key_mem[1][113] ),
    .ZN(_19182_));
 AOI22_X1 _25276_ (.A1(\core.keymem.key_mem[3][113] ),
    .A2(_16387_),
    .B1(_16463_),
    .B2(\core.keymem.key_mem[9][113] ),
    .ZN(_19183_));
 AOI22_X1 _25277_ (.A1(\core.keymem.key_mem[7][113] ),
    .A2(_16513_),
    .B1(_17675_),
    .B2(\core.keymem.key_mem[5][113] ),
    .ZN(_19184_));
 AOI22_X1 _25278_ (.A1(\core.keymem.key_mem[4][113] ),
    .A2(_16458_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][113] ),
    .ZN(_19185_));
 AND4_X1 _25279_ (.A1(_19182_),
    .A2(_19183_),
    .A3(_19184_),
    .A4(_19185_),
    .ZN(_19186_));
 AOI22_X2 _25280_ (.A1(\core.keymem.key_mem[6][113] ),
    .A2(_16522_),
    .B1(_17769_),
    .B2(\core.keymem.key_mem[11][113] ),
    .ZN(_19187_));
 AOI22_X2 _25281_ (.A1(\core.keymem.key_mem[2][113] ),
    .A2(_17086_),
    .B1(_17765_),
    .B2(\core.keymem.key_mem[8][113] ),
    .ZN(_19188_));
 AOI22_X2 _25282_ (.A1(\core.keymem.key_mem[14][113] ),
    .A2(_17581_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][113] ),
    .ZN(_19189_));
 NAND4_X2 _25283_ (.A1(_19186_),
    .A2(_19187_),
    .A3(_19188_),
    .A4(_19189_),
    .ZN(_19190_));
 OAI21_X4 _25284_ (.A(_19181_),
    .B1(_19190_),
    .B2(_16549_),
    .ZN(_19191_));
 XNOR2_X2 _25285_ (.A(_19033_),
    .B(_19191_),
    .ZN(_19192_));
 AND2_X1 _25286_ (.A1(_00267_),
    .A2(_16496_),
    .ZN(_19193_));
 INV_X1 _25287_ (.A(\core.keymem.key_mem[12][17] ),
    .ZN(_19194_));
 INV_X1 _25288_ (.A(\core.keymem.key_mem[2][17] ),
    .ZN(_19195_));
 OAI33_X1 _25289_ (.A1(_19194_),
    .A2(_16390_),
    .A3(_16394_),
    .B1(_16383_),
    .B2(_16421_),
    .B3(_19195_),
    .ZN(_19196_));
 AOI221_X1 _25290_ (.A(_19196_),
    .B1(_16415_),
    .B2(\core.keymem.key_mem[1][17] ),
    .C1(\core.keymem.key_mem[3][17] ),
    .C2(_16865_),
    .ZN(_19197_));
 OAI211_X2 _25291_ (.A(\core.keymem.key_mem[13][17] ),
    .B(_16882_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_19198_));
 OAI211_X2 _25292_ (.A(\core.keymem.key_mem[7][17] ),
    .B(_17048_),
    .C1(_17114_),
    .C2(_17115_),
    .ZN(_19199_));
 NAND3_X1 _25293_ (.A1(\core.keymem.key_mem[14][17] ),
    .A2(_16882_),
    .A3(_17016_),
    .ZN(_19200_));
 OAI211_X2 _25294_ (.A(\core.keymem.key_mem[10][17] ),
    .B(_17156_),
    .C1(_16886_),
    .C2(_16890_),
    .ZN(_19201_));
 AND4_X1 _25295_ (.A1(_19198_),
    .A2(_19199_),
    .A3(_19200_),
    .A4(_19201_),
    .ZN(_19202_));
 OAI211_X2 _25296_ (.A(\core.keymem.key_mem[6][17] ),
    .B(_17156_),
    .C1(_17115_),
    .C2(_17146_),
    .ZN(_19203_));
 OAI211_X2 _25297_ (.A(\core.keymem.key_mem[11][17] ),
    .B(_17111_),
    .C1(_17128_),
    .C2(_17129_),
    .ZN(_19204_));
 OAI211_X2 _25298_ (.A(\core.keymem.key_mem[8][17] ),
    .B(_17527_),
    .C1(_16886_),
    .C2(_16890_),
    .ZN(_19205_));
 OAI221_X1 _25299_ (.A(\core.keymem.key_mem[9][17] ),
    .B1(_17035_),
    .B2(_17036_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_19206_));
 AND4_X1 _25300_ (.A1(_19203_),
    .A2(_19204_),
    .A3(_19205_),
    .A4(_19206_),
    .ZN(_19207_));
 AOI22_X1 _25301_ (.A1(\core.keymem.key_mem[4][17] ),
    .A2(_17713_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][17] ),
    .ZN(_19208_));
 AND4_X2 _25302_ (.A1(_19197_),
    .A2(_19202_),
    .A3(_19207_),
    .A4(_19208_),
    .ZN(_19209_));
 AOI21_X4 _25303_ (.A(_19193_),
    .B1(_19209_),
    .B2(_16489_),
    .ZN(_19210_));
 XNOR2_X2 _25304_ (.A(\block_reg[3][17] ),
    .B(_19210_),
    .ZN(_19211_));
 OAI221_X2 _25305_ (.A(_16364_),
    .B1(_19180_),
    .B2(_19192_),
    .C1(_19211_),
    .C2(_17710_),
    .ZN(_19212_));
 NAND2_X1 _25306_ (.A1(_00252_),
    .A2(_16497_),
    .ZN(_19213_));
 AOI22_X4 _25307_ (.A1(\core.keymem.key_mem[2][14] ),
    .A2(_16424_),
    .B1(_16386_),
    .B2(\core.keymem.key_mem[3][14] ),
    .ZN(_19214_));
 AOI22_X1 _25308_ (.A1(\core.keymem.key_mem[8][14] ),
    .A2(_16452_),
    .B1(_16432_),
    .B2(\core.keymem.key_mem[10][14] ),
    .ZN(_19215_));
 AOI22_X1 _25309_ (.A1(\core.keymem.key_mem[6][14] ),
    .A2(_16520_),
    .B1(_16472_),
    .B2(\core.keymem.key_mem[13][14] ),
    .ZN(_19216_));
 AOI22_X1 _25310_ (.A1(\core.keymem.key_mem[4][14] ),
    .A2(_16947_),
    .B1(_17736_),
    .B2(\core.keymem.key_mem[7][14] ),
    .ZN(_19217_));
 AND4_X1 _25311_ (.A1(_19214_),
    .A2(_19215_),
    .A3(_19216_),
    .A4(_19217_),
    .ZN(_19218_));
 AOI22_X4 _25312_ (.A1(\core.keymem.key_mem[12][14] ),
    .A2(_16540_),
    .B1(_16417_),
    .B2(\core.keymem.key_mem[1][14] ),
    .ZN(_19219_));
 AOI22_X2 _25313_ (.A1(\core.keymem.key_mem[9][14] ),
    .A2(_16463_),
    .B1(_17675_),
    .B2(\core.keymem.key_mem[5][14] ),
    .ZN(_19220_));
 AOI22_X2 _25314_ (.A1(\core.keymem.key_mem[14][14] ),
    .A2(_16439_),
    .B1(_16443_),
    .B2(\core.keymem.key_mem[11][14] ),
    .ZN(_19221_));
 NAND4_X4 _25315_ (.A1(_19218_),
    .A2(_19219_),
    .A3(_19220_),
    .A4(_19221_),
    .ZN(_19222_));
 OAI21_X4 _25316_ (.A(_19213_),
    .B1(_19222_),
    .B2(_16497_),
    .ZN(_19223_));
 XOR2_X2 _25317_ (.A(_17248_),
    .B(_19223_),
    .Z(_19224_));
 XNOR2_X2 _25318_ (.A(_18970_),
    .B(_19224_),
    .ZN(_19225_));
 XNOR2_X2 _25319_ (.A(\core.dec_block.block_w3_reg[16] ),
    .B(_18859_),
    .ZN(_19226_));
 XOR2_X1 _25320_ (.A(_18909_),
    .B(_19226_),
    .Z(_19227_));
 XNOR2_X1 _25321_ (.A(_19225_),
    .B(_19227_),
    .ZN(_19228_));
 XNOR2_X2 _25322_ (.A(_19016_),
    .B(_19228_),
    .ZN(_19229_));
 AOI22_X1 _25323_ (.A1(\core.keymem.key_mem[7][30] ),
    .A2(_16954_),
    .B1(_16450_),
    .B2(\core.keymem.key_mem[8][30] ),
    .ZN(_19230_));
 AOI22_X1 _25324_ (.A1(\core.keymem.key_mem[11][30] ),
    .A2(_16504_),
    .B1(_16470_),
    .B2(\core.keymem.key_mem[13][30] ),
    .ZN(_19231_));
 NAND2_X1 _25325_ (.A1(_19230_),
    .A2(_19231_),
    .ZN(_19232_));
 AOI221_X2 _25326_ (.A(_16967_),
    .B1(_16483_),
    .B2(\core.keymem.key_mem[12][30] ),
    .C1(\core.keymem.key_mem[14][30] ),
    .C2(_16906_),
    .ZN(_19233_));
 AOI21_X1 _25327_ (.A(_16972_),
    .B1(_16484_),
    .B2(\core.keymem.key_mem[4][30] ),
    .ZN(_19234_));
 OAI21_X1 _25328_ (.A(_16961_),
    .B1(_19233_),
    .B2(_19234_),
    .ZN(_19235_));
 NAND3_X1 _25329_ (.A1(\core.keymem.key_mem[1][30] ),
    .A2(_16964_),
    .A3(_16967_),
    .ZN(_19236_));
 NAND3_X1 _25330_ (.A1(\core.keymem.key_mem[10][30] ),
    .A2(_17025_),
    .A3(_16972_),
    .ZN(_19237_));
 NAND3_X1 _25331_ (.A1(_16958_),
    .A2(_19236_),
    .A3(_19237_),
    .ZN(_19238_));
 INV_X1 _25332_ (.A(\core.keymem.key_mem[5][30] ),
    .ZN(_19239_));
 INV_X1 _25333_ (.A(\core.keymem.key_mem[9][30] ),
    .ZN(_19240_));
 OAI22_X2 _25334_ (.A1(_19239_),
    .A2(_17042_),
    .B1(_17529_),
    .B2(_19240_),
    .ZN(_19241_));
 AOI221_X2 _25335_ (.A(_19232_),
    .B1(_19235_),
    .B2(_19238_),
    .C1(_16964_),
    .C2(_19241_),
    .ZN(_19242_));
 MUX2_X1 _25336_ (.A(\core.keymem.key_mem[2][30] ),
    .B(\core.keymem.key_mem[6][30] ),
    .S(_16960_),
    .Z(_19243_));
 AOI221_X2 _25337_ (.A(_16544_),
    .B1(_18985_),
    .B2(_19243_),
    .C1(_16986_),
    .C2(\core.keymem.key_mem[3][30] ),
    .ZN(_19244_));
 AOI22_X4 _25338_ (.A1(_00296_),
    .A2(_16496_),
    .B1(_19242_),
    .B2(_19244_),
    .ZN(_19245_));
 XNOR2_X2 _25339_ (.A(\core.dec_block.block_w3_reg[30] ),
    .B(_19245_),
    .ZN(_19246_));
 XNOR2_X2 _25340_ (.A(_19002_),
    .B(_19246_),
    .ZN(_19247_));
 XNOR2_X2 _25341_ (.A(_19229_),
    .B(_19247_),
    .ZN(_19248_));
 NAND2_X1 _25342_ (.A1(_00213_),
    .A2(_17014_),
    .ZN(_19249_));
 AOI22_X1 _25343_ (.A1(\core.keymem.key_mem[10][7] ),
    .A2(_16514_),
    .B1(_16854_),
    .B2(\core.keymem.key_mem[1][7] ),
    .ZN(_19250_));
 AOI22_X1 _25344_ (.A1(\core.keymem.key_mem[3][7] ),
    .A2(_16865_),
    .B1(_16535_),
    .B2(\core.keymem.key_mem[9][7] ),
    .ZN(_19251_));
 AOI22_X1 _25345_ (.A1(\core.keymem.key_mem[7][7] ),
    .A2(_16955_),
    .B1(_16467_),
    .B2(\core.keymem.key_mem[5][7] ),
    .ZN(_19252_));
 AOI22_X1 _25346_ (.A1(\core.keymem.key_mem[4][7] ),
    .A2(_16946_),
    .B1(_16397_),
    .B2(\core.keymem.key_mem[12][7] ),
    .ZN(_19253_));
 AND4_X1 _25347_ (.A1(_19250_),
    .A2(_19251_),
    .A3(_19252_),
    .A4(_19253_),
    .ZN(_19254_));
 AOI22_X2 _25348_ (.A1(\core.keymem.key_mem[6][7] ),
    .A2(_17695_),
    .B1(_16442_),
    .B2(\core.keymem.key_mem[11][7] ),
    .ZN(_19255_));
 AOI22_X4 _25349_ (.A1(\core.keymem.key_mem[2][7] ),
    .A2(_16860_),
    .B1(_16529_),
    .B2(\core.keymem.key_mem[8][7] ),
    .ZN(_19256_));
 AOI22_X2 _25350_ (.A1(\core.keymem.key_mem[14][7] ),
    .A2(_17719_),
    .B1(_16532_),
    .B2(\core.keymem.key_mem[13][7] ),
    .ZN(_19257_));
 NAND4_X4 _25351_ (.A1(_19254_),
    .A2(_19255_),
    .A3(_19256_),
    .A4(_19257_),
    .ZN(_19258_));
 OAI21_X4 _25352_ (.A(_19249_),
    .B1(_19258_),
    .B2(_16872_),
    .ZN(_19259_));
 XOR2_X2 _25353_ (.A(\core.dec_block.block_w3_reg[7] ),
    .B(_19259_),
    .Z(_19260_));
 XNOR2_X2 _25354_ (.A(_18896_),
    .B(_18942_),
    .ZN(_19261_));
 XNOR2_X2 _25355_ (.A(_19260_),
    .B(_19261_),
    .ZN(_19262_));
 NAND2_X2 _25356_ (.A1(_00227_),
    .A2(_17183_),
    .ZN(_19263_));
 AOI222_X2 _25357_ (.A1(\core.keymem.key_mem[6][9] ),
    .A2(_16449_),
    .B1(_16994_),
    .B2(\core.keymem.key_mem[2][9] ),
    .C1(_17005_),
    .C2(\core.keymem.key_mem[5][9] ),
    .ZN(_19264_));
 AOI22_X2 _25358_ (.A1(\core.keymem.key_mem[11][9] ),
    .A2(_16507_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][9] ),
    .ZN(_19265_));
 AOI22_X2 _25359_ (.A1(\core.keymem.key_mem[7][9] ),
    .A2(_16513_),
    .B1(_16537_),
    .B2(\core.keymem.key_mem[9][9] ),
    .ZN(_19266_));
 NAND3_X2 _25360_ (.A1(_19264_),
    .A2(_19265_),
    .A3(_19266_),
    .ZN(_19267_));
 AOI21_X1 _25361_ (.A(_16983_),
    .B1(_17178_),
    .B2(\core.keymem.key_mem[1][9] ),
    .ZN(_19268_));
 AOI22_X2 _25362_ (.A1(\core.keymem.key_mem[3][9] ),
    .A2(_16387_),
    .B1(_16433_),
    .B2(\core.keymem.key_mem[10][9] ),
    .ZN(_19269_));
 AOI22_X2 _25363_ (.A1(\core.keymem.key_mem[8][9] ),
    .A2(_16453_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][9] ),
    .ZN(_19270_));
 AOI22_X2 _25364_ (.A1(\core.keymem.key_mem[4][9] ),
    .A2(_16458_),
    .B1(_16439_),
    .B2(\core.keymem.key_mem[14][9] ),
    .ZN(_19271_));
 NAND4_X2 _25365_ (.A1(_19268_),
    .A2(_19269_),
    .A3(_19270_),
    .A4(_19271_),
    .ZN(_19272_));
 OAI21_X4 _25366_ (.A(_19263_),
    .B1(_19267_),
    .B2(_19272_),
    .ZN(_19273_));
 XOR2_X2 _25367_ (.A(\core.dec_block.block_w3_reg[9] ),
    .B(_19273_),
    .Z(_19274_));
 AOI222_X2 _25368_ (.A1(\core.keymem.key_mem[14][1] ),
    .A2(_17719_),
    .B1(_16424_),
    .B2(\core.keymem.key_mem[2][1] ),
    .C1(_17175_),
    .C2(\core.keymem.key_mem[3][1] ),
    .ZN(_19275_));
 AOI22_X1 _25369_ (.A1(\core.keymem.key_mem[10][1] ),
    .A2(_16989_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][1] ),
    .ZN(_19276_));
 AOI22_X1 _25370_ (.A1(\core.keymem.key_mem[4][1] ),
    .A2(_17713_),
    .B1(_17720_),
    .B2(\core.keymem.key_mem[12][1] ),
    .ZN(_19277_));
 AND3_X1 _25371_ (.A1(_19275_),
    .A2(_19276_),
    .A3(_19277_),
    .ZN(_19278_));
 AOI22_X1 _25372_ (.A1(\core.keymem.key_mem[11][1] ),
    .A2(_17008_),
    .B1(_16855_),
    .B2(\core.keymem.key_mem[1][1] ),
    .ZN(_19279_));
 AOI22_X1 _25373_ (.A1(\core.keymem.key_mem[6][1] ),
    .A2(_17695_),
    .B1(_16529_),
    .B2(\core.keymem.key_mem[8][1] ),
    .ZN(_19280_));
 AOI22_X1 _25374_ (.A1(\core.keymem.key_mem[7][1] ),
    .A2(_16512_),
    .B1(_16462_),
    .B2(\core.keymem.key_mem[9][1] ),
    .ZN(_19281_));
 AOI21_X1 _25375_ (.A(_16982_),
    .B1(_16509_),
    .B2(\core.keymem.key_mem[5][1] ),
    .ZN(_19282_));
 AND4_X1 _25376_ (.A1(_19279_),
    .A2(_19280_),
    .A3(_19281_),
    .A4(_19282_),
    .ZN(_19283_));
 AOI22_X4 _25377_ (.A1(_00187_),
    .A2(_16497_),
    .B1(_19278_),
    .B2(_19283_),
    .ZN(_19284_));
 XNOR2_X2 _25378_ (.A(\core.dec_block.block_w3_reg[1] ),
    .B(_19284_),
    .ZN(_19285_));
 AOI22_X1 _25379_ (.A1(\core.keymem.key_mem[11][25] ),
    .A2(_17008_),
    .B1(_16855_),
    .B2(\core.keymem.key_mem[1][25] ),
    .ZN(_19286_));
 AOI22_X1 _25380_ (.A1(\core.keymem.key_mem[8][25] ),
    .A2(_17666_),
    .B1(_16536_),
    .B2(\core.keymem.key_mem[9][25] ),
    .ZN(_19287_));
 AOI22_X1 _25381_ (.A1(\core.keymem.key_mem[4][25] ),
    .A2(_17713_),
    .B1(_16512_),
    .B2(\core.keymem.key_mem[7][25] ),
    .ZN(_19288_));
 AOI21_X1 _25382_ (.A(_16495_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][25] ),
    .ZN(_19289_));
 NAND4_X1 _25383_ (.A1(_19286_),
    .A2(_19287_),
    .A3(_19288_),
    .A4(_19289_),
    .ZN(_19290_));
 MUX2_X1 _25384_ (.A(\core.keymem.key_mem[6][25] ),
    .B(\core.keymem.key_mem[14][25] ),
    .S(_17054_),
    .Z(_19291_));
 AOI22_X1 _25385_ (.A1(\core.keymem.key_mem[2][25] ),
    .A2(_17121_),
    .B1(_17051_),
    .B2(_19291_),
    .ZN(_19292_));
 NOR2_X1 _25386_ (.A1(_16968_),
    .A2(_19292_),
    .ZN(_19293_));
 AOI22_X1 _25387_ (.A1(\core.keymem.key_mem[10][25] ),
    .A2(_17715_),
    .B1(_16509_),
    .B2(\core.keymem.key_mem[5][25] ),
    .ZN(_19294_));
 AOI22_X1 _25388_ (.A1(\core.keymem.key_mem[3][25] ),
    .A2(_16866_),
    .B1(_16539_),
    .B2(\core.keymem.key_mem[12][25] ),
    .ZN(_19295_));
 NAND2_X1 _25389_ (.A1(_19294_),
    .A2(_19295_),
    .ZN(_19296_));
 NOR3_X2 _25390_ (.A1(_19290_),
    .A2(_19293_),
    .A3(_19296_),
    .ZN(_19297_));
 AOI21_X4 _25391_ (.A(_19297_),
    .B1(_16873_),
    .B2(_00298_),
    .ZN(_19298_));
 XNOR2_X2 _25392_ (.A(\core.dec_block.block_w3_reg[25] ),
    .B(_19298_),
    .ZN(_19299_));
 XNOR2_X2 _25393_ (.A(_19285_),
    .B(_19299_),
    .ZN(_19300_));
 XNOR2_X1 _25394_ (.A(_19274_),
    .B(_19300_),
    .ZN(_19301_));
 XNOR2_X1 _25395_ (.A(_19262_),
    .B(_19301_),
    .ZN(_19302_));
 XNOR2_X1 _25396_ (.A(_19248_),
    .B(_19302_),
    .ZN(_19303_));
 AOI21_X1 _25397_ (.A(_19212_),
    .B1(_19303_),
    .B2(_18332_),
    .ZN(_19304_));
 AOI22_X1 _25398_ (.A1(_19033_),
    .A2(_17744_),
    .B1(_19179_),
    .B2(_19304_),
    .ZN(_00575_));
 NOR2_X1 _25399_ (.A1(\core.dec_block.block_w0_reg[18] ),
    .A2(_18330_),
    .ZN(_19305_));
 OAI21_X1 _25400_ (.A(_18629_),
    .B1(_18740_),
    .B2(_18806_),
    .ZN(_19306_));
 NOR2_X1 _25401_ (.A1(_18629_),
    .A2(_18770_),
    .ZN(_19307_));
 NAND3_X1 _25402_ (.A1(_18716_),
    .A2(_18699_),
    .A3(_19307_),
    .ZN(_19308_));
 AOI21_X1 _25403_ (.A(_18635_),
    .B1(_19306_),
    .B2(_19308_),
    .ZN(_19309_));
 OAI22_X1 _25404_ (.A1(_18820_),
    .A2(_18747_),
    .B1(_19150_),
    .B2(_18666_),
    .ZN(_19310_));
 AOI21_X1 _25405_ (.A(_19310_),
    .B1(_19142_),
    .B2(_18680_),
    .ZN(_19311_));
 OAI221_X2 _25406_ (.A(_19311_),
    .B1(_19136_),
    .B2(_18744_),
    .C1(_18693_),
    .C2(_19164_),
    .ZN(_19312_));
 MUX2_X1 _25407_ (.A(_18820_),
    .B(_19134_),
    .S(_18658_),
    .Z(_19313_));
 NAND2_X2 _25408_ (.A1(_19034_),
    .A2(_18796_),
    .ZN(_19314_));
 OAI21_X1 _25409_ (.A(_19138_),
    .B1(_19313_),
    .B2(_19314_),
    .ZN(_19315_));
 OR3_X1 _25410_ (.A1(_19309_),
    .A2(_19312_),
    .A3(_19315_),
    .ZN(_19316_));
 NAND2_X4 _25411_ (.A1(_18623_),
    .A2(_18746_),
    .ZN(_19317_));
 OAI22_X1 _25412_ (.A1(_18705_),
    .A2(_18801_),
    .B1(_19317_),
    .B2(_18693_),
    .ZN(_19318_));
 NAND2_X1 _25413_ (.A1(_18700_),
    .A2(_19318_),
    .ZN(_19319_));
 NOR3_X1 _25414_ (.A1(_18699_),
    .A2(_19052_),
    .A3(_18722_),
    .ZN(_19320_));
 OAI21_X1 _25415_ (.A(_18722_),
    .B1(_18672_),
    .B2(_18659_),
    .ZN(_19321_));
 NOR2_X4 _25416_ (.A1(_18573_),
    .A2(_18612_),
    .ZN(_19322_));
 AOI21_X1 _25417_ (.A(_19320_),
    .B1(_19321_),
    .B2(_19322_),
    .ZN(_19323_));
 OAI21_X1 _25418_ (.A(_19319_),
    .B1(_19323_),
    .B2(_18817_),
    .ZN(_19324_));
 NAND2_X1 _25419_ (.A1(_18723_),
    .A2(_18780_),
    .ZN(_19325_));
 OAI21_X1 _25420_ (.A(_18823_),
    .B1(_18780_),
    .B2(_18765_),
    .ZN(_19326_));
 AOI21_X1 _25421_ (.A(_19052_),
    .B1(_19325_),
    .B2(_19326_),
    .ZN(_19327_));
 NAND3_X1 _25422_ (.A1(_18647_),
    .A2(_18654_),
    .A3(_18774_),
    .ZN(_19328_));
 AOI22_X1 _25423_ (.A1(_18688_),
    .A2(_18680_),
    .B1(_18726_),
    .B2(_18702_),
    .ZN(_19329_));
 OAI21_X1 _25424_ (.A(_19328_),
    .B1(_19329_),
    .B2(_18654_),
    .ZN(_19330_));
 NOR4_X1 _25425_ (.A1(_19316_),
    .A2(_19324_),
    .A3(_19327_),
    .A4(_19330_),
    .ZN(_19331_));
 MUX2_X1 _25426_ (.A(_18712_),
    .B(_18765_),
    .S(_18823_),
    .Z(_19332_));
 NAND3_X1 _25427_ (.A1(_18789_),
    .A2(_18700_),
    .A3(_19332_),
    .ZN(_19333_));
 NOR2_X2 _25428_ (.A1(_18653_),
    .A2(_18692_),
    .ZN(_19334_));
 AOI21_X1 _25429_ (.A(_18731_),
    .B1(_18597_),
    .B2(_18719_),
    .ZN(_19335_));
 NAND2_X1 _25430_ (.A1(_18581_),
    .A2(_18796_),
    .ZN(_19336_));
 OAI33_X1 _25431_ (.A1(_18581_),
    .A2(_18717_),
    .A3(_19335_),
    .B1(_19336_),
    .B2(_18741_),
    .B3(_18750_),
    .ZN(_19337_));
 AOI221_X2 _25432_ (.A(_19334_),
    .B1(_19337_),
    .B2(_18633_),
    .C1(_18823_),
    .C2(_18708_),
    .ZN(_19338_));
 OAI21_X1 _25433_ (.A(_19333_),
    .B1(_19338_),
    .B2(_18789_),
    .ZN(_19339_));
 NAND2_X1 _25434_ (.A1(_18806_),
    .A2(_19339_),
    .ZN(_19340_));
 NOR3_X1 _25435_ (.A1(_18816_),
    .A2(_18699_),
    .A3(_19172_),
    .ZN(_19341_));
 AOI21_X1 _25436_ (.A(_19111_),
    .B1(_18688_),
    .B2(_18708_),
    .ZN(_19342_));
 OAI22_X1 _25437_ (.A1(_18598_),
    .A2(_19052_),
    .B1(_19342_),
    .B2(_18723_),
    .ZN(_19343_));
 AOI21_X2 _25438_ (.A(_19341_),
    .B1(_19343_),
    .B2(_18817_),
    .ZN(_19344_));
 OAI22_X1 _25439_ (.A1(_18640_),
    .A2(_18672_),
    .B1(_19168_),
    .B2(_19040_),
    .ZN(_19345_));
 AOI222_X2 _25440_ (.A1(_18842_),
    .A2(_19053_),
    .B1(_19345_),
    .B2(_18736_),
    .C1(_19070_),
    .C2(_18686_),
    .ZN(_19346_));
 AOI21_X1 _25441_ (.A(_18599_),
    .B1(_18636_),
    .B2(_19034_),
    .ZN(_19347_));
 OR3_X1 _25442_ (.A1(_18832_),
    .A2(_18808_),
    .A3(_19347_),
    .ZN(_19348_));
 NAND3_X2 _25443_ (.A1(_19344_),
    .A2(_19346_),
    .A3(_19348_),
    .ZN(_19349_));
 NOR2_X1 _25444_ (.A1(_18655_),
    .A2(_18708_),
    .ZN(_19350_));
 AOI221_X2 _25445_ (.A(_18782_),
    .B1(_18655_),
    .B2(_18820_),
    .C1(_19122_),
    .C2(_19350_),
    .ZN(_19351_));
 NOR4_X1 _25446_ (.A1(_18823_),
    .A2(_18807_),
    .A3(_19040_),
    .A4(_18810_),
    .ZN(_19352_));
 NAND3_X1 _25447_ (.A1(_18666_),
    .A2(_18651_),
    .A3(_18810_),
    .ZN(_19353_));
 AOI21_X1 _25448_ (.A(_19352_),
    .B1(_19353_),
    .B2(_18761_),
    .ZN(_19354_));
 NOR2_X2 _25449_ (.A1(_18694_),
    .A2(_18638_),
    .ZN(_19355_));
 OAI21_X1 _25450_ (.A(_18783_),
    .B1(_18753_),
    .B2(_19355_),
    .ZN(_19356_));
 NOR2_X1 _25451_ (.A1(_18620_),
    .A2(_18723_),
    .ZN(_19357_));
 NOR2_X2 _25452_ (.A1(_18745_),
    .A2(_18732_),
    .ZN(_19358_));
 OAI221_X1 _25453_ (.A(_19357_),
    .B1(_19358_),
    .B2(_18768_),
    .C1(_18806_),
    .C2(_18817_),
    .ZN(_19359_));
 NAND3_X1 _25454_ (.A1(_19354_),
    .A2(_19356_),
    .A3(_19359_),
    .ZN(_19360_));
 NOR4_X2 _25455_ (.A1(_18772_),
    .A2(_19349_),
    .A3(_19351_),
    .A4(_19360_),
    .ZN(_19361_));
 OAI21_X1 _25456_ (.A(_18779_),
    .B1(_19082_),
    .B2(_19355_),
    .ZN(_19362_));
 NAND2_X2 _25457_ (.A1(_18697_),
    .A2(_19081_),
    .ZN(_19363_));
 NAND2_X1 _25458_ (.A1(_18815_),
    .A2(_18609_),
    .ZN(_19364_));
 OAI221_X2 _25459_ (.A(_19362_),
    .B1(_19363_),
    .B2(_18810_),
    .C1(_18693_),
    .C2(_19364_),
    .ZN(_19365_));
 OAI21_X1 _25460_ (.A(_18681_),
    .B1(_18719_),
    .B2(_19034_),
    .ZN(_19366_));
 MUX2_X1 _25461_ (.A(_18793_),
    .B(_19366_),
    .S(_18621_),
    .Z(_19367_));
 OAI21_X1 _25462_ (.A(_18709_),
    .B1(_19168_),
    .B2(_18807_),
    .ZN(_19368_));
 AOI221_X2 _25463_ (.A(_19365_),
    .B1(_19367_),
    .B2(_19071_),
    .C1(_18628_),
    .C2(_19368_),
    .ZN(_19369_));
 AND2_X1 _25464_ (.A1(_19101_),
    .A2(_19369_),
    .ZN(_19370_));
 AND4_X2 _25465_ (.A1(_19331_),
    .A2(_19340_),
    .A3(_19361_),
    .A4(_19370_),
    .ZN(_19371_));
 AOI22_X1 _25466_ (.A1(\core.keymem.key_mem[11][114] ),
    .A2(_16443_),
    .B1(_17675_),
    .B2(\core.keymem.key_mem[5][114] ),
    .ZN(_19372_));
 AOI22_X1 _25467_ (.A1(\core.keymem.key_mem[4][114] ),
    .A2(_18232_),
    .B1(_17781_),
    .B2(\core.keymem.key_mem[8][114] ),
    .ZN(_19373_));
 AOI22_X1 _25468_ (.A1(\core.keymem.key_mem[7][114] ),
    .A2(_16408_),
    .B1(_16433_),
    .B2(\core.keymem.key_mem[10][114] ),
    .ZN(_19374_));
 AOI21_X1 _25469_ (.A(_16871_),
    .B1(_16417_),
    .B2(\core.keymem.key_mem[1][114] ),
    .ZN(_19375_));
 NAND4_X1 _25470_ (.A1(_19372_),
    .A2(_19373_),
    .A3(_19374_),
    .A4(_19375_),
    .ZN(_19376_));
 MUX2_X1 _25471_ (.A(\core.keymem.key_mem[6][114] ),
    .B(\core.keymem.key_mem[14][114] ),
    .S(_17054_),
    .Z(_19377_));
 AOI22_X1 _25472_ (.A1(\core.keymem.key_mem[2][114] ),
    .A2(_17121_),
    .B1(_17051_),
    .B2(_19377_),
    .ZN(_19378_));
 NOR2_X1 _25473_ (.A1(_16968_),
    .A2(_19378_),
    .ZN(_19379_));
 AOI22_X1 _25474_ (.A1(\core.keymem.key_mem[3][114] ),
    .A2(_17683_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][114] ),
    .ZN(_19380_));
 AOI22_X1 _25475_ (.A1(\core.keymem.key_mem[9][114] ),
    .A2(_16463_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][114] ),
    .ZN(_19381_));
 NAND2_X1 _25476_ (.A1(_19380_),
    .A2(_19381_),
    .ZN(_19382_));
 NOR3_X2 _25477_ (.A1(_19376_),
    .A2(_19379_),
    .A3(_19382_),
    .ZN(_19383_));
 AOI21_X4 _25478_ (.A(_19383_),
    .B1(_16548_),
    .B2(_00197_),
    .ZN(_19384_));
 XNOR2_X2 _25479_ (.A(\core.dec_block.block_w0_reg[18] ),
    .B(_19384_),
    .ZN(_19385_));
 AOI222_X2 _25480_ (.A1(\core.keymem.key_mem[14][18] ),
    .A2(_16439_),
    .B1(_17781_),
    .B2(\core.keymem.key_mem[8][18] ),
    .C1(\core.keymem.key_mem[4][18] ),
    .C2(_17713_),
    .ZN(_19386_));
 AOI22_X1 _25481_ (.A1(\core.keymem.key_mem[1][18] ),
    .A2(_17178_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][18] ),
    .ZN(_19387_));
 AOI22_X1 _25482_ (.A1(\core.keymem.key_mem[7][18] ),
    .A2(_16513_),
    .B1(_16516_),
    .B2(\core.keymem.key_mem[10][18] ),
    .ZN(_19388_));
 NAND3_X1 _25483_ (.A1(_19386_),
    .A2(_19387_),
    .A3(_19388_),
    .ZN(_19389_));
 AOI22_X1 _25484_ (.A1(\core.keymem.key_mem[6][18] ),
    .A2(_16449_),
    .B1(_16443_),
    .B2(\core.keymem.key_mem[11][18] ),
    .ZN(_19390_));
 AOI22_X1 _25485_ (.A1(\core.keymem.key_mem[2][18] ),
    .A2(_16425_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][18] ),
    .ZN(_19391_));
 AOI22_X1 _25486_ (.A1(\core.keymem.key_mem[3][18] ),
    .A2(_17683_),
    .B1(_17675_),
    .B2(\core.keymem.key_mem[5][18] ),
    .ZN(_19392_));
 AOI21_X1 _25487_ (.A(_16546_),
    .B1(_16537_),
    .B2(\core.keymem.key_mem[9][18] ),
    .ZN(_19393_));
 NAND4_X1 _25488_ (.A1(_19390_),
    .A2(_19391_),
    .A3(_19392_),
    .A4(_19393_),
    .ZN(_19394_));
 NOR2_X2 _25489_ (.A1(_19389_),
    .A2(_19394_),
    .ZN(_19395_));
 AOI21_X4 _25490_ (.A(_19395_),
    .B1(_16498_),
    .B2(_00275_),
    .ZN(_19396_));
 XNOR2_X2 _25491_ (.A(\block_reg[3][18] ),
    .B(_19396_),
    .ZN(_19397_));
 OAI221_X2 _25492_ (.A(_18329_),
    .B1(_17741_),
    .B2(_19385_),
    .C1(_19397_),
    .C2(_18553_),
    .ZN(_19398_));
 AOI22_X1 _25493_ (.A1(\core.keymem.key_mem[4][10] ),
    .A2(_17513_),
    .B1(_17067_),
    .B2(\core.keymem.key_mem[8][10] ),
    .ZN(_19399_));
 NOR2_X1 _25494_ (.A1(_16394_),
    .A2(_19399_),
    .ZN(_19400_));
 AOI22_X1 _25495_ (.A1(\core.keymem.key_mem[6][10] ),
    .A2(_16447_),
    .B1(_16385_),
    .B2(\core.keymem.key_mem[3][10] ),
    .ZN(_19401_));
 AOI22_X1 _25496_ (.A1(\core.keymem.key_mem[10][10] ),
    .A2(_16431_),
    .B1(_16471_),
    .B2(\core.keymem.key_mem[13][10] ),
    .ZN(_19402_));
 NAND2_X1 _25497_ (.A1(_19401_),
    .A2(_19402_),
    .ZN(_19403_));
 AOI22_X1 _25498_ (.A1(\core.keymem.key_mem[2][10] ),
    .A2(_16858_),
    .B1(_16948_),
    .B2(\core.keymem.key_mem[5][10] ),
    .ZN(_19404_));
 AOI22_X1 _25499_ (.A1(\core.keymem.key_mem[14][10] ),
    .A2(_16436_),
    .B1(_16523_),
    .B2(\core.keymem.key_mem[1][10] ),
    .ZN(_19405_));
 AOI22_X1 _25500_ (.A1(\core.keymem.key_mem[9][10] ),
    .A2(_16461_),
    .B1(_16504_),
    .B2(\core.keymem.key_mem[11][10] ),
    .ZN(_19406_));
 AOI22_X1 _25501_ (.A1(\core.keymem.key_mem[7][10] ),
    .A2(_16954_),
    .B1(_16396_),
    .B2(\core.keymem.key_mem[12][10] ),
    .ZN(_19407_));
 NAND4_X1 _25502_ (.A1(_19404_),
    .A2(_19405_),
    .A3(_19406_),
    .A4(_19407_),
    .ZN(_19408_));
 OR4_X2 _25503_ (.A1(_17013_),
    .A2(_19400_),
    .A3(_19403_),
    .A4(_19408_),
    .ZN(_19409_));
 INV_X1 _25504_ (.A(_00235_),
    .ZN(_19410_));
 OAI21_X4 _25505_ (.A(_19409_),
    .B1(_17533_),
    .B2(_19410_),
    .ZN(_19411_));
 XOR2_X2 _25506_ (.A(\core.dec_block.block_w3_reg[10] ),
    .B(_19411_),
    .Z(_19412_));
 XNOR2_X2 _25507_ (.A(_18942_),
    .B(_19412_),
    .ZN(_19413_));
 XNOR2_X2 _25508_ (.A(_19224_),
    .B(_19413_),
    .ZN(_19414_));
 XNOR2_X1 _25509_ (.A(_18921_),
    .B(_19226_),
    .ZN(_19415_));
 XNOR2_X1 _25510_ (.A(_18884_),
    .B(_19027_),
    .ZN(_19416_));
 XNOR2_X1 _25511_ (.A(_19415_),
    .B(_19416_),
    .ZN(_19417_));
 AOI222_X2 _25512_ (.A1(\core.keymem.key_mem[4][26] ),
    .A2(_16457_),
    .B1(_16424_),
    .B2(\core.keymem.key_mem[2][26] ),
    .C1(_16998_),
    .C2(\core.keymem.key_mem[14][26] ),
    .ZN(_19418_));
 AOI22_X1 _25513_ (.A1(\core.keymem.key_mem[8][26] ),
    .A2(_17666_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][26] ),
    .ZN(_19419_));
 AOI22_X1 _25514_ (.A1(\core.keymem.key_mem[1][26] ),
    .A2(_16525_),
    .B1(_16509_),
    .B2(\core.keymem.key_mem[5][26] ),
    .ZN(_19420_));
 NAND3_X1 _25515_ (.A1(_19418_),
    .A2(_19419_),
    .A3(_19420_),
    .ZN(_19421_));
 AOI22_X1 _25516_ (.A1(\core.keymem.key_mem[10][26] ),
    .A2(_17715_),
    .B1(_16506_),
    .B2(\core.keymem.key_mem[11][26] ),
    .ZN(_19422_));
 AOI22_X1 _25517_ (.A1(\core.keymem.key_mem[7][26] ),
    .A2(_16512_),
    .B1(_16448_),
    .B2(\core.keymem.key_mem[6][26] ),
    .ZN(_19423_));
 AOI22_X1 _25518_ (.A1(\core.keymem.key_mem[9][26] ),
    .A2(_16536_),
    .B1(_16398_),
    .B2(\core.keymem.key_mem[12][26] ),
    .ZN(_19424_));
 AOI21_X1 _25519_ (.A(_16982_),
    .B1(_16866_),
    .B2(\core.keymem.key_mem[3][26] ),
    .ZN(_19425_));
 NAND4_X1 _25520_ (.A1(_19422_),
    .A2(_19423_),
    .A3(_19424_),
    .A4(_19425_),
    .ZN(_19426_));
 NOR2_X2 _25521_ (.A1(_19421_),
    .A2(_19426_),
    .ZN(_19427_));
 AOI21_X4 _25522_ (.A(_19427_),
    .B1(_16497_),
    .B2(_00299_),
    .ZN(_19428_));
 XNOR2_X2 _25523_ (.A(\core.dec_block.block_w3_reg[26] ),
    .B(_19428_),
    .ZN(_19429_));
 XNOR2_X2 _25524_ (.A(_19246_),
    .B(_19429_),
    .ZN(_19430_));
 AOI21_X1 _25525_ (.A(_16544_),
    .B1(_16461_),
    .B2(\core.keymem.key_mem[9][31] ),
    .ZN(_19431_));
 AOI22_X1 _25526_ (.A1(\core.keymem.key_mem[6][31] ),
    .A2(_16519_),
    .B1(_16450_),
    .B2(\core.keymem.key_mem[8][31] ),
    .ZN(_19432_));
 AOI22_X1 _25527_ (.A1(\core.keymem.key_mem[11][31] ),
    .A2(_16504_),
    .B1(_16466_),
    .B2(\core.keymem.key_mem[5][31] ),
    .ZN(_19433_));
 AOI22_X1 _25528_ (.A1(\core.keymem.key_mem[12][31] ),
    .A2(_16396_),
    .B1(_16470_),
    .B2(\core.keymem.key_mem[13][31] ),
    .ZN(_19434_));
 AND4_X2 _25529_ (.A1(_19431_),
    .A2(_19432_),
    .A3(_19433_),
    .A4(_19434_),
    .ZN(_19435_));
 AOI222_X2 _25530_ (.A1(\core.keymem.key_mem[2][31] ),
    .A2(_16858_),
    .B1(_16864_),
    .B2(\core.keymem.key_mem[3][31] ),
    .C1(\core.keymem.key_mem[10][31] ),
    .C2(_16430_),
    .ZN(_19436_));
 AOI22_X1 _25531_ (.A1(\core.keymem.key_mem[4][31] ),
    .A2(_16946_),
    .B1(_16523_),
    .B2(\core.keymem.key_mem[1][31] ),
    .ZN(_19437_));
 AOI22_X1 _25532_ (.A1(\core.keymem.key_mem[14][31] ),
    .A2(_16436_),
    .B1(_16954_),
    .B2(\core.keymem.key_mem[7][31] ),
    .ZN(_19438_));
 AND3_X2 _25533_ (.A1(_19436_),
    .A2(_19437_),
    .A3(_19438_),
    .ZN(_19439_));
 AOI22_X4 _25534_ (.A1(_00297_),
    .A2(_17013_),
    .B1(_19435_),
    .B2(_19439_),
    .ZN(_19440_));
 XNOR2_X2 _25535_ (.A(\core.dec_block.block_w3_reg[31] ),
    .B(_19440_),
    .ZN(_19441_));
 XNOR2_X2 _25536_ (.A(_19430_),
    .B(_19441_),
    .ZN(_19442_));
 XNOR2_X1 _25537_ (.A(_19417_),
    .B(_19442_),
    .ZN(_19443_));
 XNOR2_X2 _25538_ (.A(_19414_),
    .B(_19443_),
    .ZN(_19444_));
 XNOR2_X2 _25539_ (.A(\core.dec_block.block_w3_reg[17] ),
    .B(_19210_),
    .ZN(_19445_));
 XNOR2_X2 _25540_ (.A(_19274_),
    .B(_19445_),
    .ZN(_19446_));
 AOI22_X1 _25541_ (.A1(\core.keymem.key_mem[2][2] ),
    .A2(_17786_),
    .B1(_16525_),
    .B2(\core.keymem.key_mem[1][2] ),
    .ZN(_19447_));
 AOI22_X1 _25542_ (.A1(\core.keymem.key_mem[9][2] ),
    .A2(_17668_),
    .B1(_16539_),
    .B2(\core.keymem.key_mem[12][2] ),
    .ZN(_19448_));
 AOI22_X1 _25543_ (.A1(\core.keymem.key_mem[8][2] ),
    .A2(_17666_),
    .B1(_16506_),
    .B2(\core.keymem.key_mem[11][2] ),
    .ZN(_19449_));
 AOI22_X1 _25544_ (.A1(\core.keymem.key_mem[7][2] ),
    .A2(_17084_),
    .B1(_16448_),
    .B2(\core.keymem.key_mem[6][2] ),
    .ZN(_19450_));
 NAND4_X1 _25545_ (.A1(_19447_),
    .A2(_19448_),
    .A3(_19449_),
    .A4(_19450_),
    .ZN(_19451_));
 AOI22_X1 _25546_ (.A1(\core.keymem.key_mem[4][2] ),
    .A2(_17713_),
    .B1(_16866_),
    .B2(\core.keymem.key_mem[3][2] ),
    .ZN(_19452_));
 AOI22_X1 _25547_ (.A1(\core.keymem.key_mem[5][2] ),
    .A2(_16509_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][2] ),
    .ZN(_19453_));
 AOI22_X1 _25548_ (.A1(\core.keymem.key_mem[14][2] ),
    .A2(_17719_),
    .B1(_17715_),
    .B2(\core.keymem.key_mem[10][2] ),
    .ZN(_19454_));
 NAND3_X1 _25549_ (.A1(_19452_),
    .A2(_19453_),
    .A3(_19454_),
    .ZN(_19455_));
 NOR3_X2 _25550_ (.A1(_16547_),
    .A2(_19451_),
    .A3(_19455_),
    .ZN(_19456_));
 AOI21_X4 _25551_ (.A(_19456_),
    .B1(_16548_),
    .B2(_00195_),
    .ZN(_19457_));
 XNOR2_X2 _25552_ (.A(\core.dec_block.block_w3_reg[2] ),
    .B(_19457_),
    .ZN(_19458_));
 XOR2_X1 _25553_ (.A(_19446_),
    .B(_19458_),
    .Z(_19459_));
 XNOR2_X1 _25554_ (.A(_19444_),
    .B(_19459_),
    .ZN(_19460_));
 AOI21_X1 _25555_ (.A(_19398_),
    .B1(_19460_),
    .B2(_19031_),
    .ZN(_19461_));
 AOI21_X1 _25556_ (.A(_19305_),
    .B1(_19371_),
    .B2(_19461_),
    .ZN(_00576_));
 INV_X1 _25557_ (.A(\core.dec_block.block_w0_reg[19] ),
    .ZN(_19462_));
 OAI22_X1 _25558_ (.A1(_18684_),
    .A2(_18640_),
    .B1(_19317_),
    .B2(_18643_),
    .ZN(_19463_));
 AOI22_X2 _25559_ (.A1(_18815_),
    .A2(_18783_),
    .B1(_19463_),
    .B2(_18634_),
    .ZN(_19464_));
 NOR2_X1 _25560_ (.A1(_18700_),
    .A2(_19464_),
    .ZN(_19465_));
 OAI22_X4 _25561_ (.A1(_18820_),
    .A2(_19135_),
    .B1(_19139_),
    .B2(_19134_),
    .ZN(_19466_));
 AOI21_X1 _25562_ (.A(_18794_),
    .B1(_18776_),
    .B2(_19144_),
    .ZN(_19467_));
 AOI221_X1 _25563_ (.A(_19467_),
    .B1(_18774_),
    .B2(_18712_),
    .C1(_18662_),
    .C2(_18740_),
    .ZN(_19468_));
 OAI21_X1 _25564_ (.A(_19468_),
    .B1(_18687_),
    .B2(_18689_),
    .ZN(_19469_));
 NOR4_X1 _25565_ (.A1(_19349_),
    .A2(_19465_),
    .A3(_19466_),
    .A4(_19469_),
    .ZN(_19470_));
 NOR3_X1 _25566_ (.A1(_18715_),
    .A2(_18758_),
    .A3(_18736_),
    .ZN(_19471_));
 NOR3_X1 _25567_ (.A1(_18805_),
    .A2(_18676_),
    .A3(_18722_),
    .ZN(_19472_));
 NOR3_X1 _25568_ (.A1(_18789_),
    .A2(_19471_),
    .A3(_19472_),
    .ZN(_19473_));
 NOR4_X2 _25569_ (.A1(_18763_),
    .A2(_18741_),
    .A3(_18676_),
    .A4(_19045_),
    .ZN(_19474_));
 NOR2_X1 _25570_ (.A1(_19034_),
    .A2(_18581_),
    .ZN(_19475_));
 NAND3_X1 _25571_ (.A1(_18631_),
    .A2(_18609_),
    .A3(_18752_),
    .ZN(_19476_));
 OAI21_X1 _25572_ (.A(_19476_),
    .B1(_18633_),
    .B2(_18643_),
    .ZN(_19477_));
 OAI22_X2 _25573_ (.A1(_18722_),
    .A2(_18797_),
    .B1(_19076_),
    .B2(_18723_),
    .ZN(_19478_));
 AOI221_X2 _25574_ (.A(_19474_),
    .B1(_19475_),
    .B2(_19477_),
    .C1(_18655_),
    .C2(_19478_),
    .ZN(_19479_));
 AOI21_X1 _25575_ (.A(_19473_),
    .B1(_19479_),
    .B2(_18789_),
    .ZN(_19480_));
 NAND2_X1 _25576_ (.A1(_18573_),
    .A2(_18623_),
    .ZN(_19481_));
 OR3_X1 _25577_ (.A1(_18788_),
    .A2(_19481_),
    .A3(_18672_),
    .ZN(_19482_));
 OAI21_X1 _25578_ (.A(_18823_),
    .B1(_18666_),
    .B2(_18716_),
    .ZN(_19483_));
 NAND2_X1 _25579_ (.A1(_18715_),
    .A2(_18686_),
    .ZN(_19484_));
 OAI21_X1 _25580_ (.A(_19484_),
    .B1(_18820_),
    .B2(_18716_),
    .ZN(_19485_));
 OAI21_X1 _25581_ (.A(_19483_),
    .B1(_19485_),
    .B2(_18823_),
    .ZN(_19486_));
 OAI21_X1 _25582_ (.A(_19482_),
    .B1(_19486_),
    .B2(_18659_),
    .ZN(_19487_));
 AOI21_X1 _25583_ (.A(_19480_),
    .B1(_19487_),
    .B2(_18700_),
    .ZN(_19488_));
 NAND2_X1 _25584_ (.A1(_19470_),
    .A2(_19488_),
    .ZN(_19489_));
 NOR2_X1 _25585_ (.A1(_18699_),
    .A2(_19134_),
    .ZN(_19490_));
 OAI21_X1 _25586_ (.A(_18659_),
    .B1(_19071_),
    .B2(_19490_),
    .ZN(_19491_));
 MUX2_X1 _25587_ (.A(_18662_),
    .B(_18680_),
    .S(_18620_),
    .Z(_19492_));
 AOI221_X2 _25588_ (.A(_18673_),
    .B1(_18840_),
    .B2(_18703_),
    .C1(_19492_),
    .C2(_18805_),
    .ZN(_19493_));
 NAND3_X1 _25589_ (.A1(_18817_),
    .A2(_19491_),
    .A3(_19493_),
    .ZN(_19494_));
 NAND3_X1 _25590_ (.A1(_18807_),
    .A2(_18703_),
    .A3(_18783_),
    .ZN(_19495_));
 NAND2_X1 _25591_ (.A1(_18698_),
    .A2(_18842_),
    .ZN(_19496_));
 AOI22_X1 _25592_ (.A1(_18789_),
    .A2(_18712_),
    .B1(_19357_),
    .B2(_18686_),
    .ZN(_19497_));
 OAI221_X1 _25593_ (.A(_19495_),
    .B1(_19496_),
    .B2(_19052_),
    .C1(_18716_),
    .C2(_19497_),
    .ZN(_19498_));
 OAI21_X1 _25594_ (.A(_19494_),
    .B1(_19498_),
    .B2(_18817_),
    .ZN(_19499_));
 NOR2_X1 _25595_ (.A1(_18651_),
    .A2(_18776_),
    .ZN(_19500_));
 OAI33_X1 _25596_ (.A1(_18674_),
    .A2(_18681_),
    .A3(_18732_),
    .B1(_19093_),
    .B2(_18638_),
    .B3(_18675_),
    .ZN(_19501_));
 NOR3_X1 _25597_ (.A1(_18730_),
    .A2(_19500_),
    .A3(_19501_),
    .ZN(_19502_));
 NOR3_X1 _25598_ (.A1(_18648_),
    .A2(_18639_),
    .A3(_18671_),
    .ZN(_19503_));
 AOI21_X1 _25599_ (.A(_19503_),
    .B1(_18774_),
    .B2(_18662_),
    .ZN(_19504_));
 OAI21_X1 _25600_ (.A(_19502_),
    .B1(_19504_),
    .B2(_18654_),
    .ZN(_19505_));
 OAI21_X1 _25601_ (.A(_18832_),
    .B1(_18636_),
    .B2(_19035_),
    .ZN(_19506_));
 OAI21_X1 _25602_ (.A(_19506_),
    .B1(_18766_),
    .B2(_18832_),
    .ZN(_19507_));
 NAND2_X1 _25603_ (.A1(_18717_),
    .A2(_19507_),
    .ZN(_19508_));
 NOR3_X1 _25604_ (.A1(_18782_),
    .A2(_18808_),
    .A3(_19134_),
    .ZN(_19509_));
 OAI222_X2 _25605_ (.A1(_18749_),
    .A2(_19094_),
    .B1(_19150_),
    .B2(_18801_),
    .C1(_18692_),
    .C2(_19317_),
    .ZN(_19510_));
 AOI21_X1 _25606_ (.A(_18598_),
    .B1(_19363_),
    .B2(_19150_),
    .ZN(_19511_));
 OR2_X1 _25607_ (.A1(_19510_),
    .A2(_19511_),
    .ZN(_19512_));
 OAI21_X1 _25608_ (.A(_18736_),
    .B1(_18778_),
    .B2(_18686_),
    .ZN(_19513_));
 AOI21_X1 _25609_ (.A(_19040_),
    .B1(_18696_),
    .B2(_19513_),
    .ZN(_19514_));
 NOR3_X1 _25610_ (.A1(_19509_),
    .A2(_19512_),
    .A3(_19514_),
    .ZN(_19515_));
 NAND3_X1 _25611_ (.A1(_19078_),
    .A2(_19508_),
    .A3(_19515_),
    .ZN(_19516_));
 NOR3_X1 _25612_ (.A1(_19167_),
    .A2(_19505_),
    .A3(_19516_),
    .ZN(_19517_));
 NAND2_X1 _25613_ (.A1(_19499_),
    .A2(_19517_),
    .ZN(_19518_));
 NOR3_X4 _25614_ (.A1(_18847_),
    .A2(_19489_),
    .A3(_19518_),
    .ZN(_19519_));
 AOI22_X1 _25615_ (.A1(\core.keymem.key_mem[3][115] ),
    .A2(_16387_),
    .B1(_16463_),
    .B2(\core.keymem.key_mem[9][115] ),
    .ZN(_19520_));
 AOI22_X1 _25616_ (.A1(\core.keymem.key_mem[2][115] ),
    .A2(_16994_),
    .B1(_17781_),
    .B2(\core.keymem.key_mem[8][115] ),
    .ZN(_19521_));
 AOI22_X1 _25617_ (.A1(\core.keymem.key_mem[10][115] ),
    .A2(_16433_),
    .B1(_17768_),
    .B2(\core.keymem.key_mem[11][115] ),
    .ZN(_19522_));
 AOI22_X1 _25618_ (.A1(\core.keymem.key_mem[4][115] ),
    .A2(_18232_),
    .B1(_17001_),
    .B2(\core.keymem.key_mem[12][115] ),
    .ZN(_19523_));
 NAND4_X1 _25619_ (.A1(_19520_),
    .A2(_19521_),
    .A3(_19522_),
    .A4(_19523_),
    .ZN(_19524_));
 AOI22_X1 _25620_ (.A1(\core.keymem.key_mem[14][115] ),
    .A2(_16502_),
    .B1(_16991_),
    .B2(\core.keymem.key_mem[6][115] ),
    .ZN(_19525_));
 AOI22_X1 _25621_ (.A1(\core.keymem.key_mem[7][115] ),
    .A2(_16408_),
    .B1(_16417_),
    .B2(\core.keymem.key_mem[1][115] ),
    .ZN(_19526_));
 AOI22_X1 _25622_ (.A1(\core.keymem.key_mem[5][115] ),
    .A2(_17675_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][115] ),
    .ZN(_19527_));
 NAND3_X1 _25623_ (.A1(_19525_),
    .A2(_19526_),
    .A3(_19527_),
    .ZN(_19528_));
 NOR2_X1 _25624_ (.A1(_19524_),
    .A2(_19528_),
    .ZN(_19529_));
 MUX2_X2 _25625_ (.A(_00203_),
    .B(_19529_),
    .S(_16489_),
    .Z(_03286_));
 XNOR2_X2 _25626_ (.A(_19462_),
    .B(_03286_),
    .ZN(_03287_));
 AOI22_X1 _25627_ (.A1(\core.keymem.key_mem[10][19] ),
    .A2(_16433_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][19] ),
    .ZN(_03288_));
 AOI22_X1 _25628_ (.A1(\core.keymem.key_mem[7][19] ),
    .A2(_17789_),
    .B1(_17003_),
    .B2(\core.keymem.key_mem[1][19] ),
    .ZN(_03289_));
 AOI22_X1 _25629_ (.A1(\core.keymem.key_mem[9][19] ),
    .A2(_17914_),
    .B1(_17008_),
    .B2(\core.keymem.key_mem[11][19] ),
    .ZN(_03290_));
 AOI22_X1 _25630_ (.A1(\core.keymem.key_mem[2][19] ),
    .A2(_17786_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][19] ),
    .ZN(_03291_));
 NAND4_X1 _25631_ (.A1(_03288_),
    .A2(_03289_),
    .A3(_03290_),
    .A4(_03291_),
    .ZN(_03292_));
 AOI22_X1 _25632_ (.A1(\core.keymem.key_mem[14][19] ),
    .A2(_16439_),
    .B1(_17683_),
    .B2(\core.keymem.key_mem[3][19] ),
    .ZN(_03293_));
 AOI22_X1 _25633_ (.A1(\core.keymem.key_mem[4][19] ),
    .A2(_18232_),
    .B1(_17781_),
    .B2(\core.keymem.key_mem[8][19] ),
    .ZN(_03294_));
 AOI22_X1 _25634_ (.A1(\core.keymem.key_mem[6][19] ),
    .A2(_16991_),
    .B1(_17001_),
    .B2(\core.keymem.key_mem[12][19] ),
    .ZN(_03295_));
 NAND3_X1 _25635_ (.A1(_03293_),
    .A2(_03294_),
    .A3(_03295_),
    .ZN(_03296_));
 NOR3_X2 _25636_ (.A1(_16497_),
    .A2(_03292_),
    .A3(_03296_),
    .ZN(_03297_));
 AOI21_X4 _25637_ (.A(_03297_),
    .B1(_16498_),
    .B2(_00281_),
    .ZN(_03298_));
 XNOR2_X1 _25638_ (.A(\block_reg[3][19] ),
    .B(_03298_),
    .ZN(_03299_));
 OAI221_X2 _25639_ (.A(_16364_),
    .B1(_19180_),
    .B2(_03287_),
    .C1(_03299_),
    .C2(_17710_),
    .ZN(_03300_));
 XNOR2_X2 _25640_ (.A(_19004_),
    .B(_19226_),
    .ZN(_03301_));
 XNOR2_X2 _25641_ (.A(_19016_),
    .B(_19260_),
    .ZN(_03302_));
 XNOR2_X1 _25642_ (.A(_18956_),
    .B(_03302_),
    .ZN(_03303_));
 XNOR2_X1 _25643_ (.A(_19285_),
    .B(_19445_),
    .ZN(_03304_));
 AND2_X1 _25644_ (.A1(_00300_),
    .A2(_17014_),
    .ZN(_03305_));
 OAI211_X2 _25645_ (.A(\core.keymem.key_mem[13][27] ),
    .B(_17100_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_03306_));
 OAI211_X2 _25646_ (.A(\core.keymem.key_mem[6][27] ),
    .B(_17101_),
    .C1(_17106_),
    .C2(_17107_),
    .ZN(_03307_));
 NAND3_X1 _25647_ (.A1(\core.keymem.key_mem[2][27] ),
    .A2(_17121_),
    .A3(_17101_),
    .ZN(_03308_));
 OAI211_X2 _25648_ (.A(\core.keymem.key_mem[8][27] ),
    .B(_17057_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_03309_));
 NAND4_X2 _25649_ (.A1(_03306_),
    .A2(_03307_),
    .A3(_03308_),
    .A4(_03309_),
    .ZN(_03310_));
 OAI211_X2 _25650_ (.A(\core.keymem.key_mem[7][27] ),
    .B(_17112_),
    .C1(_17107_),
    .C2(_17106_),
    .ZN(_03311_));
 NAND3_X1 _25651_ (.A1(\core.keymem.key_mem[3][27] ),
    .A2(_17112_),
    .A3(_17121_),
    .ZN(_03312_));
 NAND3_X1 _25652_ (.A1(\core.keymem.key_mem[14][27] ),
    .A2(_17100_),
    .A3(_17101_),
    .ZN(_03313_));
 OAI211_X2 _25653_ (.A(\core.keymem.key_mem[4][27] ),
    .B(_17057_),
    .C1(_17107_),
    .C2(_17106_),
    .ZN(_03314_));
 NAND4_X2 _25654_ (.A1(_03311_),
    .A2(_03312_),
    .A3(_03313_),
    .A4(_03314_),
    .ZN(_03315_));
 OAI211_X2 _25655_ (.A(\core.keymem.key_mem[10][27] ),
    .B(_17050_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_03316_));
 OAI211_X2 _25656_ (.A(\core.keymem.key_mem[11][27] ),
    .B(_17112_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_03317_));
 OAI221_X2 _25657_ (.A(\core.keymem.key_mem[5][27] ),
    .B1(_17114_),
    .B2(_17115_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_03318_));
 OAI221_X2 _25658_ (.A(\core.keymem.key_mem[9][27] ),
    .B1(_17128_),
    .B2(_17129_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_03319_));
 NAND4_X2 _25659_ (.A1(_03316_),
    .A2(_03317_),
    .A3(_03318_),
    .A4(_03319_),
    .ZN(_03320_));
 INV_X1 _25660_ (.A(\core.keymem.key_mem[12][27] ),
    .ZN(_03321_));
 INV_X2 _25661_ (.A(\core.keymem.key_mem[1][27] ),
    .ZN(_03322_));
 OAI22_X4 _25662_ (.A1(_03321_),
    .A2(_17843_),
    .B1(_18545_),
    .B2(_03322_),
    .ZN(_03323_));
 NOR4_X4 _25663_ (.A1(_03310_),
    .A2(_03315_),
    .A3(_03320_),
    .A4(_03323_),
    .ZN(_03324_));
 AOI21_X4 _25664_ (.A(_03305_),
    .B1(_03324_),
    .B2(_16489_),
    .ZN(_03325_));
 XNOR2_X2 _25665_ (.A(\core.dec_block.block_w3_reg[27] ),
    .B(_03325_),
    .ZN(_03326_));
 XNOR2_X2 _25666_ (.A(_19441_),
    .B(_03326_),
    .ZN(_03327_));
 XNOR2_X1 _25667_ (.A(_03304_),
    .B(_03327_),
    .ZN(_03328_));
 XNOR2_X1 _25668_ (.A(_18922_),
    .B(_03328_),
    .ZN(_03329_));
 XNOR2_X1 _25669_ (.A(_03303_),
    .B(_03329_),
    .ZN(_03330_));
 XNOR2_X2 _25670_ (.A(_03301_),
    .B(_03330_),
    .ZN(_03331_));
 XNOR2_X2 _25671_ (.A(\core.dec_block.block_w3_reg[18] ),
    .B(_19396_),
    .ZN(_03332_));
 XNOR2_X2 _25672_ (.A(_18956_),
    .B(_03332_),
    .ZN(_03333_));
 AOI22_X1 _25673_ (.A1(\core.keymem.key_mem[6][11] ),
    .A2(_16520_),
    .B1(_17000_),
    .B2(\core.keymem.key_mem[12][11] ),
    .ZN(_03334_));
 AOI22_X1 _25674_ (.A1(\core.keymem.key_mem[9][11] ),
    .A2(_17522_),
    .B1(_17007_),
    .B2(\core.keymem.key_mem[11][11] ),
    .ZN(_03335_));
 AOI21_X1 _25675_ (.A(_16545_),
    .B1(_16416_),
    .B2(\core.keymem.key_mem[1][11] ),
    .ZN(_03336_));
 AOI22_X1 _25676_ (.A1(\core.keymem.key_mem[3][11] ),
    .A2(_17175_),
    .B1(_17193_),
    .B2(\core.keymem.key_mem[13][11] ),
    .ZN(_03337_));
 AND4_X1 _25677_ (.A1(_03334_),
    .A2(_03335_),
    .A3(_03336_),
    .A4(_03337_),
    .ZN(_03338_));
 AOI222_X2 _25678_ (.A1(\core.keymem.key_mem[4][11] ),
    .A2(_16499_),
    .B1(_16859_),
    .B2(\core.keymem.key_mem[2][11] ),
    .C1(_16437_),
    .C2(\core.keymem.key_mem[14][11] ),
    .ZN(_03339_));
 AOI22_X1 _25679_ (.A1(\core.keymem.key_mem[10][11] ),
    .A2(_16432_),
    .B1(_17004_),
    .B2(\core.keymem.key_mem[5][11] ),
    .ZN(_03340_));
 AOI22_X1 _25680_ (.A1(\core.keymem.key_mem[7][11] ),
    .A2(_16407_),
    .B1(_17506_),
    .B2(\core.keymem.key_mem[8][11] ),
    .ZN(_03341_));
 AND3_X1 _25681_ (.A1(_03339_),
    .A2(_03340_),
    .A3(_03341_),
    .ZN(_03342_));
 AOI22_X4 _25682_ (.A1(_00241_),
    .A2(_16852_),
    .B1(_03338_),
    .B2(_03342_),
    .ZN(_03343_));
 XNOR2_X2 _25683_ (.A(_17216_),
    .B(_03343_),
    .ZN(_03344_));
 XNOR2_X1 _25684_ (.A(_03333_),
    .B(_03344_),
    .ZN(_03345_));
 AOI222_X2 _25685_ (.A1(\core.keymem.key_mem[3][3] ),
    .A2(_16987_),
    .B1(_16525_),
    .B2(\core.keymem.key_mem[1][3] ),
    .C1(_16539_),
    .C2(\core.keymem.key_mem[12][3] ),
    .ZN(_03346_));
 AOI22_X2 _25686_ (.A1(\core.keymem.key_mem[4][3] ),
    .A2(_18232_),
    .B1(_16994_),
    .B2(\core.keymem.key_mem[2][3] ),
    .ZN(_03347_));
 AOI22_X2 _25687_ (.A1(\core.keymem.key_mem[10][3] ),
    .A2(_16433_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][3] ),
    .ZN(_03348_));
 NAND3_X2 _25688_ (.A1(_03346_),
    .A2(_03347_),
    .A3(_03348_),
    .ZN(_03349_));
 AOI22_X1 _25689_ (.A1(\core.keymem.key_mem[6][3] ),
    .A2(_16991_),
    .B1(_17768_),
    .B2(\core.keymem.key_mem[11][3] ),
    .ZN(_03350_));
 AOI22_X2 _25690_ (.A1(\core.keymem.key_mem[14][3] ),
    .A2(_16999_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][3] ),
    .ZN(_03351_));
 AOI22_X2 _25691_ (.A1(\core.keymem.key_mem[8][3] ),
    .A2(_17781_),
    .B1(_17914_),
    .B2(\core.keymem.key_mem[9][3] ),
    .ZN(_03352_));
 AOI21_X1 _25692_ (.A(_16871_),
    .B1(_16408_),
    .B2(\core.keymem.key_mem[7][3] ),
    .ZN(_03353_));
 NAND4_X2 _25693_ (.A1(_03350_),
    .A2(_03351_),
    .A3(_03352_),
    .A4(_03353_),
    .ZN(_03354_));
 NOR2_X4 _25694_ (.A1(_03349_),
    .A2(_03354_),
    .ZN(_03355_));
 AND2_X1 _25695_ (.A1(_00201_),
    .A2(_16852_),
    .ZN(_03356_));
 NOR2_X4 _25696_ (.A1(_03355_),
    .A2(_03356_),
    .ZN(_03357_));
 XNOR2_X2 _25697_ (.A(\core.dec_block.block_w3_reg[3] ),
    .B(_03357_),
    .ZN(_03358_));
 XOR2_X1 _25698_ (.A(_19027_),
    .B(_03358_),
    .Z(_03359_));
 XNOR2_X1 _25699_ (.A(_19412_),
    .B(_03359_),
    .ZN(_03360_));
 XNOR2_X1 _25700_ (.A(_18897_),
    .B(_03360_),
    .ZN(_03361_));
 XNOR2_X1 _25701_ (.A(_03345_),
    .B(_03361_),
    .ZN(_03362_));
 XNOR2_X1 _25702_ (.A(_03331_),
    .B(_03362_),
    .ZN(_03363_));
 AOI21_X1 _25703_ (.A(_03300_),
    .B1(_03363_),
    .B2(_18332_),
    .ZN(_03364_));
 AOI22_X1 _25704_ (.A1(_19462_),
    .A2(_17744_),
    .B1(_19519_),
    .B2(_03364_),
    .ZN(_00577_));
 INV_X1 _25705_ (.A(\core.dec_block.block_w0_reg[1] ),
    .ZN(_03365_));
 NAND2_X4 _25706_ (.A1(_16644_),
    .A2(_16580_),
    .ZN(_03366_));
 MUX2_X1 _25707_ (.A(_16670_),
    .B(_03366_),
    .S(_16623_),
    .Z(_03367_));
 NOR3_X1 _25708_ (.A1(_16669_),
    .A2(_16668_),
    .A3(_03367_),
    .ZN(_03368_));
 NAND3_X1 _25709_ (.A1(_16623_),
    .A2(_16669_),
    .A3(_03366_),
    .ZN(_03369_));
 OAI21_X1 _25710_ (.A(_03369_),
    .B1(_16669_),
    .B2(_16648_),
    .ZN(_03370_));
 AOI21_X1 _25711_ (.A(_03368_),
    .B1(_03370_),
    .B2(_16628_),
    .ZN(_03371_));
 AOI21_X1 _25712_ (.A(_16747_),
    .B1(_16790_),
    .B2(_16675_),
    .ZN(_03372_));
 OAI22_X2 _25713_ (.A1(_16808_),
    .A2(_03371_),
    .B1(_03372_),
    .B2(_16715_),
    .ZN(_03373_));
 AOI22_X2 _25714_ (.A1(_16638_),
    .A2(_16704_),
    .B1(_03373_),
    .B2(_16754_),
    .ZN(_03374_));
 NAND2_X1 _25715_ (.A1(_16650_),
    .A2(_16775_),
    .ZN(_03375_));
 OAI221_X1 _25716_ (.A(_16698_),
    .B1(_16631_),
    .B2(_16741_),
    .C1(_03375_),
    .C2(_16796_),
    .ZN(_03376_));
 OAI21_X1 _25717_ (.A(_16732_),
    .B1(_16676_),
    .B2(_16662_),
    .ZN(_03377_));
 OAI21_X1 _25718_ (.A(_03376_),
    .B1(_03377_),
    .B2(_16754_),
    .ZN(_03378_));
 OAI21_X2 _25719_ (.A(_03374_),
    .B1(_03378_),
    .B2(_16655_),
    .ZN(_03379_));
 NAND3_X1 _25720_ (.A1(_16666_),
    .A2(_16828_),
    .A3(_03366_),
    .ZN(_03380_));
 NAND2_X2 _25721_ (.A1(_16632_),
    .A2(_16626_),
    .ZN(_03381_));
 NAND2_X4 _25722_ (.A1(_16661_),
    .A2(_16679_),
    .ZN(_03382_));
 OAI221_X1 _25723_ (.A(_03380_),
    .B1(_03381_),
    .B2(_03382_),
    .C1(_16687_),
    .C2(_16725_),
    .ZN(_03383_));
 OAI22_X1 _25724_ (.A1(_16657_),
    .A2(_16609_),
    .B1(_16710_),
    .B2(_03382_),
    .ZN(_03384_));
 AOI21_X1 _25725_ (.A(_03383_),
    .B1(_03384_),
    .B2(_16782_),
    .ZN(_03385_));
 NAND2_X4 _25726_ (.A1(_16675_),
    .A2(_16575_),
    .ZN(_03386_));
 OAI21_X1 _25727_ (.A(_03386_),
    .B1(_16759_),
    .B2(_16808_),
    .ZN(_03387_));
 NAND3_X1 _25728_ (.A1(_16810_),
    .A2(_16628_),
    .A3(_03387_),
    .ZN(_03388_));
 AOI21_X1 _25729_ (.A(_16623_),
    .B1(_16662_),
    .B2(_16693_),
    .ZN(_03389_));
 AOI21_X1 _25730_ (.A(_03389_),
    .B1(_16647_),
    .B2(_16650_),
    .ZN(_03390_));
 OAI221_X2 _25731_ (.A(_03388_),
    .B1(_03390_),
    .B2(_16634_),
    .C1(_16725_),
    .C2(_16800_),
    .ZN(_03391_));
 OAI21_X1 _25732_ (.A(_16785_),
    .B1(_16689_),
    .B2(_16703_),
    .ZN(_03392_));
 OAI21_X1 _25733_ (.A(_16679_),
    .B1(_16608_),
    .B2(_16623_),
    .ZN(_03393_));
 AOI21_X1 _25734_ (.A(_16636_),
    .B1(_16668_),
    .B2(_16761_),
    .ZN(_03394_));
 OAI33_X1 _25735_ (.A1(_16675_),
    .A2(_16631_),
    .A3(_03392_),
    .B1(_03393_),
    .B2(_03394_),
    .B3(_16625_),
    .ZN(_03395_));
 OAI21_X1 _25736_ (.A(_16725_),
    .B1(_16781_),
    .B2(_16684_),
    .ZN(_03396_));
 NAND2_X2 _25737_ (.A1(_16689_),
    .A2(_16575_),
    .ZN(_03397_));
 NAND2_X1 _25738_ (.A1(_16781_),
    .A2(_03397_),
    .ZN(_03398_));
 AOI21_X2 _25739_ (.A(_03395_),
    .B1(_03396_),
    .B2(_03398_),
    .ZN(_03399_));
 MUX2_X1 _25740_ (.A(_16669_),
    .B(_16618_),
    .S(_16623_),
    .Z(_03400_));
 NAND3_X1 _25741_ (.A1(_16634_),
    .A2(_16683_),
    .A3(_03400_),
    .ZN(_03401_));
 NOR2_X2 _25742_ (.A1(_16649_),
    .A2(_16658_),
    .ZN(_03402_));
 NOR3_X1 _25743_ (.A1(_16625_),
    .A2(_16617_),
    .A3(_16817_),
    .ZN(_03403_));
 OAI21_X1 _25744_ (.A(_16635_),
    .B1(_03402_),
    .B2(_03403_),
    .ZN(_03404_));
 NOR2_X1 _25745_ (.A1(_16699_),
    .A2(_03366_),
    .ZN(_03405_));
 OAI21_X1 _25746_ (.A(_16686_),
    .B1(_16790_),
    .B2(_03405_),
    .ZN(_03406_));
 NAND4_X1 _25747_ (.A1(_03399_),
    .A2(_03401_),
    .A3(_03404_),
    .A4(_03406_),
    .ZN(_03407_));
 AOI221_X2 _25748_ (.A(_16592_),
    .B1(_16596_),
    .B2(_17329_),
    .C1(_16608_),
    .C2(_16614_),
    .ZN(_03408_));
 MUX2_X1 _25749_ (.A(_16606_),
    .B(_16681_),
    .S(_16620_),
    .Z(_03409_));
 AOI221_X2 _25750_ (.A(_03408_),
    .B1(_16666_),
    .B2(_16668_),
    .C1(_16657_),
    .C2(_03409_),
    .ZN(_03410_));
 NOR2_X1 _25751_ (.A1(_16587_),
    .A2(_03410_),
    .ZN(_03411_));
 NOR3_X1 _25752_ (.A1(_03391_),
    .A2(_03407_),
    .A3(_03411_),
    .ZN(_03412_));
 NAND3_X1 _25753_ (.A1(_16653_),
    .A2(_03385_),
    .A3(_03412_),
    .ZN(_03413_));
 NOR2_X1 _25754_ (.A1(_16593_),
    .A2(_16668_),
    .ZN(_03414_));
 OAI21_X1 _25755_ (.A(_16658_),
    .B1(_16612_),
    .B2(_16648_),
    .ZN(_03415_));
 AOI21_X1 _25756_ (.A(_03414_),
    .B1(_03415_),
    .B2(_16770_),
    .ZN(_03416_));
 NAND2_X1 _25757_ (.A1(_16669_),
    .A2(_16742_),
    .ZN(_03417_));
 NOR2_X1 _25758_ (.A1(_16670_),
    .A2(_16816_),
    .ZN(_03418_));
 NAND3_X1 _25759_ (.A1(_16657_),
    .A2(_16636_),
    .A3(_16821_),
    .ZN(_03419_));
 OAI21_X1 _25760_ (.A(_03419_),
    .B1(_16817_),
    .B2(_16821_),
    .ZN(_03420_));
 AOI221_X2 _25761_ (.A(_16648_),
    .B1(_03417_),
    .B2(_03418_),
    .C1(_03420_),
    .C2(_16617_),
    .ZN(_03421_));
 NOR2_X1 _25762_ (.A1(_16587_),
    .A2(_16646_),
    .ZN(_03422_));
 MUX2_X1 _25763_ (.A(_16620_),
    .B(_16668_),
    .S(_03422_),
    .Z(_03423_));
 AOI221_X1 _25764_ (.A(_16635_),
    .B1(_16617_),
    .B2(_16636_),
    .C1(_03423_),
    .C2(_16669_),
    .ZN(_03424_));
 OAI22_X1 _25765_ (.A1(_16636_),
    .A2(_03416_),
    .B1(_03421_),
    .B2(_03424_),
    .ZN(_03425_));
 AND2_X1 _25766_ (.A1(_16664_),
    .A2(_03425_),
    .ZN(_03426_));
 OAI33_X1 _25767_ (.A1(_16663_),
    .A2(_16682_),
    .A3(_16825_),
    .B1(_03379_),
    .B2(_03413_),
    .B3(_03426_),
    .ZN(_03427_));
 AOI21_X1 _25768_ (.A(_16659_),
    .B1(_16677_),
    .B2(_16760_),
    .ZN(_03428_));
 NOR3_X1 _25769_ (.A1(_16682_),
    .A2(_16740_),
    .A3(_03428_),
    .ZN(_03429_));
 NOR2_X1 _25770_ (.A1(_16681_),
    .A2(_16647_),
    .ZN(_03430_));
 OAI21_X1 _25771_ (.A(_03430_),
    .B1(_16717_),
    .B2(_16613_),
    .ZN(_03431_));
 NAND3_X1 _25772_ (.A1(_16796_),
    .A2(_16630_),
    .A3(_03382_),
    .ZN(_03432_));
 OAI21_X1 _25773_ (.A(_03432_),
    .B1(_16831_),
    .B2(_16745_),
    .ZN(_03433_));
 OAI221_X2 _25774_ (.A(_03431_),
    .B1(_03433_),
    .B2(_03397_),
    .C1(_16826_),
    .C2(_16699_),
    .ZN(_03434_));
 NAND2_X1 _25775_ (.A1(_16625_),
    .A2(_16761_),
    .ZN(_03435_));
 OAI21_X1 _25776_ (.A(_03435_),
    .B1(_16691_),
    .B2(_16634_),
    .ZN(_03436_));
 NAND3_X1 _25777_ (.A1(_16715_),
    .A2(_16821_),
    .A3(_03436_),
    .ZN(_03437_));
 NAND3_X1 _25778_ (.A1(_16770_),
    .A2(_16701_),
    .A3(_16782_),
    .ZN(_03438_));
 AOI21_X1 _25779_ (.A(_16769_),
    .B1(_03437_),
    .B2(_03438_),
    .ZN(_03439_));
 NAND2_X1 _25780_ (.A1(_16635_),
    .A2(_03366_),
    .ZN(_03440_));
 OAI21_X1 _25781_ (.A(_16647_),
    .B1(_16700_),
    .B2(_16650_),
    .ZN(_03441_));
 AOI222_X2 _25782_ (.A1(_16651_),
    .A2(_16725_),
    .B1(_03440_),
    .B2(_16634_),
    .C1(_16715_),
    .C2(_03441_),
    .ZN(_03442_));
 AOI21_X1 _25783_ (.A(_16659_),
    .B1(_16764_),
    .B2(_16790_),
    .ZN(_03443_));
 OAI22_X1 _25784_ (.A1(_16793_),
    .A2(_16736_),
    .B1(_03397_),
    .B2(_03443_),
    .ZN(_03444_));
 NOR3_X1 _25785_ (.A1(_03439_),
    .A2(_03442_),
    .A3(_03444_),
    .ZN(_03445_));
 NAND2_X1 _25786_ (.A1(_16625_),
    .A2(_16632_),
    .ZN(_03446_));
 NOR2_X2 _25787_ (.A1(_16635_),
    .A2(_16675_),
    .ZN(_03447_));
 OAI33_X1 _25788_ (.A1(_16753_),
    .A2(_16738_),
    .A3(_03446_),
    .B1(_03447_),
    .B2(_16685_),
    .B3(_16634_),
    .ZN(_03448_));
 NOR2_X2 _25789_ (.A1(_16635_),
    .A2(_16644_),
    .ZN(_03449_));
 OAI33_X1 _25790_ (.A1(_16715_),
    .A2(_16593_),
    .A3(_16637_),
    .B1(_16844_),
    .B2(_03449_),
    .B3(_16705_),
    .ZN(_03450_));
 AOI22_X2 _25791_ (.A1(_16798_),
    .A2(_03448_),
    .B1(_03450_),
    .B2(_16664_),
    .ZN(_03451_));
 NOR3_X1 _25792_ (.A1(_16662_),
    .A2(_16722_),
    .A3(_16800_),
    .ZN(_03452_));
 AND2_X1 _25793_ (.A1(_16746_),
    .A2(_16758_),
    .ZN(_03453_));
 AOI221_X2 _25794_ (.A(_03452_),
    .B1(_03453_),
    .B2(_16722_),
    .C1(_16704_),
    .C2(_16831_),
    .ZN(_03454_));
 NOR2_X1 _25795_ (.A1(_16823_),
    .A2(_03397_),
    .ZN(_03455_));
 OAI22_X2 _25796_ (.A1(_16692_),
    .A2(_16738_),
    .B1(_03381_),
    .B2(_16694_),
    .ZN(_03456_));
 AOI21_X2 _25797_ (.A(_03455_),
    .B1(_03456_),
    .B2(_16798_),
    .ZN(_03457_));
 NAND4_X1 _25798_ (.A1(_03445_),
    .A2(_03451_),
    .A3(_03454_),
    .A4(_03457_),
    .ZN(_03458_));
 NOR4_X1 _25799_ (.A1(_16720_),
    .A2(_03429_),
    .A3(_03434_),
    .A4(_03458_),
    .ZN(_03459_));
 NOR3_X1 _25800_ (.A1(_16655_),
    .A2(_16754_),
    .A3(_16685_),
    .ZN(_03460_));
 NAND2_X1 _25801_ (.A1(_16796_),
    .A2(_16708_),
    .ZN(_03461_));
 AOI21_X1 _25802_ (.A(_16794_),
    .B1(_16680_),
    .B2(_03461_),
    .ZN(_03462_));
 AOI21_X1 _25803_ (.A(_03462_),
    .B1(_16743_),
    .B2(_16655_),
    .ZN(_03463_));
 NOR2_X1 _25804_ (.A1(_16714_),
    .A2(_03463_),
    .ZN(_03464_));
 OAI21_X1 _25805_ (.A(_16799_),
    .B1(_03460_),
    .B2(_03464_),
    .ZN(_03465_));
 BUF_X4 _25806_ (.A(_16753_),
    .Z(_03466_));
 NOR3_X1 _25807_ (.A1(_16798_),
    .A2(_16745_),
    .A3(_16728_),
    .ZN(_03467_));
 AOI21_X1 _25808_ (.A(_16677_),
    .B1(_16680_),
    .B2(_16776_),
    .ZN(_03468_));
 OAI21_X1 _25809_ (.A(_16714_),
    .B1(_03467_),
    .B2(_03468_),
    .ZN(_03469_));
 NAND2_X4 _25810_ (.A1(_16606_),
    .A2(_16646_),
    .ZN(_03470_));
 OAI21_X1 _25811_ (.A(_03469_),
    .B1(_03470_),
    .B2(_16776_),
    .ZN(_03471_));
 NAND2_X1 _25812_ (.A1(_03466_),
    .A2(_03471_),
    .ZN(_03472_));
 NOR3_X1 _25813_ (.A1(_16810_),
    .A2(_16821_),
    .A3(_16736_),
    .ZN(_03473_));
 NOR4_X1 _25814_ (.A1(_16657_),
    .A2(_16770_),
    .A3(_16682_),
    .A4(_16691_),
    .ZN(_03474_));
 OAI21_X1 _25815_ (.A(_16636_),
    .B1(_03473_),
    .B2(_03474_),
    .ZN(_03475_));
 NOR2_X2 _25816_ (.A1(_16681_),
    .A2(_16690_),
    .ZN(_03476_));
 NAND3_X1 _25817_ (.A1(_16810_),
    .A2(_16628_),
    .A3(_03476_),
    .ZN(_03477_));
 AOI21_X1 _25818_ (.A(_16587_),
    .B1(_03475_),
    .B2(_03477_),
    .ZN(_03478_));
 NAND2_X4 _25819_ (.A1(_16741_),
    .A2(_16782_),
    .ZN(_03479_));
 OAI22_X1 _25820_ (.A1(_16694_),
    .A2(_03479_),
    .B1(_03381_),
    .B2(_16769_),
    .ZN(_03480_));
 OAI33_X1 _25821_ (.A1(_16656_),
    .A2(_16740_),
    .A3(_16732_),
    .B1(_03435_),
    .B2(_16707_),
    .B3(_16609_),
    .ZN(_03481_));
 AOI21_X1 _25822_ (.A(_03480_),
    .B1(_03481_),
    .B2(_16767_),
    .ZN(_03482_));
 NOR2_X1 _25823_ (.A1(_16798_),
    .A2(_16841_),
    .ZN(_03483_));
 AOI22_X1 _25824_ (.A1(_16760_),
    .A2(_16761_),
    .B1(_03483_),
    .B2(_16677_),
    .ZN(_03484_));
 OAI21_X1 _25825_ (.A(_03482_),
    .B1(_03484_),
    .B2(_16785_),
    .ZN(_03485_));
 OAI22_X1 _25826_ (.A1(_16764_),
    .A2(_16694_),
    .B1(_16741_),
    .B2(_16844_),
    .ZN(_03486_));
 NAND2_X1 _25827_ (.A1(_16666_),
    .A2(_03486_),
    .ZN(_03487_));
 NOR2_X2 _25828_ (.A1(_16705_),
    .A2(_16630_),
    .ZN(_03488_));
 NOR2_X1 _25829_ (.A1(_03405_),
    .A2(_03488_),
    .ZN(_03489_));
 AOI22_X1 _25830_ (.A1(_16796_),
    .A2(_16613_),
    .B1(_16740_),
    .B2(_16828_),
    .ZN(_03490_));
 OAI221_X2 _25831_ (.A(_03487_),
    .B1(_03489_),
    .B2(_16785_),
    .C1(_03490_),
    .C2(_16682_),
    .ZN(_03491_));
 AOI21_X1 _25832_ (.A(_16686_),
    .B1(_16626_),
    .B2(_16737_),
    .ZN(_03492_));
 OAI33_X1 _25833_ (.A1(_16663_),
    .A2(_16667_),
    .A3(_16692_),
    .B1(_03492_),
    .B2(_16609_),
    .B3(_16658_),
    .ZN(_03493_));
 AOI21_X2 _25834_ (.A(_03491_),
    .B1(_03493_),
    .B2(_16803_),
    .ZN(_03494_));
 NAND2_X1 _25835_ (.A1(_03385_),
    .A2(_03494_),
    .ZN(_03495_));
 NOR3_X1 _25836_ (.A1(_03478_),
    .A2(_03485_),
    .A3(_03495_),
    .ZN(_03496_));
 NAND4_X2 _25837_ (.A1(_03459_),
    .A2(_03465_),
    .A3(_03472_),
    .A4(_03496_),
    .ZN(_03497_));
 OAI21_X4 _25838_ (.A(_18416_),
    .B1(_03427_),
    .B2(_03497_),
    .ZN(_03498_));
 AOI22_X1 _25839_ (.A1(\core.keymem.key_mem[3][97] ),
    .A2(_16987_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][97] ),
    .ZN(_03499_));
 AOI22_X1 _25840_ (.A1(\core.keymem.key_mem[11][97] ),
    .A2(_17008_),
    .B1(_16509_),
    .B2(\core.keymem.key_mem[5][97] ),
    .ZN(_03500_));
 AOI22_X1 _25841_ (.A1(\core.keymem.key_mem[6][97] ),
    .A2(_16521_),
    .B1(_16529_),
    .B2(\core.keymem.key_mem[8][97] ),
    .ZN(_03501_));
 AOI22_X1 _25842_ (.A1(\core.keymem.key_mem[14][97] ),
    .A2(_17719_),
    .B1(_16539_),
    .B2(\core.keymem.key_mem[12][97] ),
    .ZN(_03502_));
 NAND4_X1 _25843_ (.A1(_03499_),
    .A2(_03500_),
    .A3(_03501_),
    .A4(_03502_),
    .ZN(_03503_));
 AOI22_X1 _25844_ (.A1(\core.keymem.key_mem[7][97] ),
    .A2(_17789_),
    .B1(_16525_),
    .B2(\core.keymem.key_mem[1][97] ),
    .ZN(_03504_));
 AOI22_X1 _25845_ (.A1(\core.keymem.key_mem[9][97] ),
    .A2(_17914_),
    .B1(_17715_),
    .B2(\core.keymem.key_mem[10][97] ),
    .ZN(_03505_));
 AOI22_X1 _25846_ (.A1(\core.keymem.key_mem[4][97] ),
    .A2(_17713_),
    .B1(_16860_),
    .B2(\core.keymem.key_mem[2][97] ),
    .ZN(_03506_));
 NAND3_X1 _25847_ (.A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .ZN(_03507_));
 NOR2_X1 _25848_ (.A1(_03503_),
    .A2(_03507_),
    .ZN(_03508_));
 MUX2_X2 _25849_ (.A(_00194_),
    .B(_03508_),
    .S(_17533_),
    .Z(_03509_));
 XNOR2_X2 _25850_ (.A(_03365_),
    .B(_03509_),
    .ZN(_03510_));
 AOI22_X1 _25851_ (.A1(\core.keymem.key_mem[3][65] ),
    .A2(_17175_),
    .B1(_17000_),
    .B2(\core.keymem.key_mem[12][65] ),
    .ZN(_03511_));
 AOI21_X1 _25852_ (.A(_16494_),
    .B1(_16407_),
    .B2(\core.keymem.key_mem[7][65] ),
    .ZN(_03512_));
 AOI22_X1 _25853_ (.A1(\core.keymem.key_mem[14][65] ),
    .A2(_16998_),
    .B1(_17007_),
    .B2(\core.keymem.key_mem[11][65] ),
    .ZN(_03513_));
 AOI22_X1 _25854_ (.A1(\core.keymem.key_mem[4][65] ),
    .A2(_16499_),
    .B1(_16988_),
    .B2(\core.keymem.key_mem[10][65] ),
    .ZN(_03514_));
 AND4_X2 _25855_ (.A1(_03511_),
    .A2(_03512_),
    .A3(_03513_),
    .A4(_03514_),
    .ZN(_03515_));
 AOI222_X2 _25856_ (.A1(\core.keymem.key_mem[6][65] ),
    .A2(_16520_),
    .B1(_16423_),
    .B2(\core.keymem.key_mem[2][65] ),
    .C1(_16415_),
    .C2(\core.keymem.key_mem[1][65] ),
    .ZN(_03516_));
 AOI22_X1 _25857_ (.A1(\core.keymem.key_mem[8][65] ),
    .A2(_16452_),
    .B1(_16472_),
    .B2(\core.keymem.key_mem[13][65] ),
    .ZN(_03517_));
 AOI22_X1 _25858_ (.A1(\core.keymem.key_mem[9][65] ),
    .A2(_17522_),
    .B1(_17004_),
    .B2(\core.keymem.key_mem[5][65] ),
    .ZN(_03518_));
 AND3_X2 _25859_ (.A1(_03516_),
    .A2(_03517_),
    .A3(_03518_),
    .ZN(_03519_));
 AOI22_X4 _25860_ (.A1(_00233_),
    .A2(_16872_),
    .B1(_03515_),
    .B2(_03519_),
    .ZN(_03520_));
 XNOR2_X1 _25861_ (.A(\block_reg[1][1] ),
    .B(_03520_),
    .ZN(_03521_));
 OAI221_X1 _25862_ (.A(_16364_),
    .B1(_19180_),
    .B2(_03510_),
    .C1(_03521_),
    .C2(_17710_),
    .ZN(_03522_));
 XNOR2_X2 _25863_ (.A(_17079_),
    .B(_17198_),
    .ZN(_03523_));
 INV_X1 _25864_ (.A(\core.dec_block.block_w1_reg[0] ),
    .ZN(_03524_));
 XNOR2_X2 _25865_ (.A(_03524_),
    .B(_16490_),
    .ZN(_03525_));
 XNOR2_X1 _25866_ (.A(_17097_),
    .B(_03525_),
    .ZN(_03526_));
 XNOR2_X2 _25867_ (.A(_03523_),
    .B(_03526_),
    .ZN(_03527_));
 NAND3_X1 _25868_ (.A1(\core.keymem.key_mem[4][94] ),
    .A2(_17057_),
    .A3(_16967_),
    .ZN(_03528_));
 NAND3_X1 _25869_ (.A1(\core.keymem.key_mem[14][94] ),
    .A2(_17016_),
    .A3(_17055_),
    .ZN(_03529_));
 AOI21_X2 _25870_ (.A(_17043_),
    .B1(_03528_),
    .B2(_03529_),
    .ZN(_03530_));
 AOI22_X1 _25871_ (.A1(\core.keymem.key_mem[6][94] ),
    .A2(_17648_),
    .B1(_16467_),
    .B2(\core.keymem.key_mem[5][94] ),
    .ZN(_03531_));
 AOI22_X2 _25872_ (.A1(\core.keymem.key_mem[3][94] ),
    .A2(_16385_),
    .B1(_16441_),
    .B2(\core.keymem.key_mem[11][94] ),
    .ZN(_03532_));
 AOI22_X2 _25873_ (.A1(\core.keymem.key_mem[7][94] ),
    .A2(_16406_),
    .B1(_16514_),
    .B2(\core.keymem.key_mem[10][94] ),
    .ZN(_03533_));
 AOI22_X2 _25874_ (.A1(\core.keymem.key_mem[8][94] ),
    .A2(_16451_),
    .B1(_16397_),
    .B2(\core.keymem.key_mem[12][94] ),
    .ZN(_03534_));
 NAND4_X2 _25875_ (.A1(_03531_),
    .A2(_03532_),
    .A3(_03533_),
    .A4(_03534_),
    .ZN(_03535_));
 AOI22_X1 _25876_ (.A1(\core.keymem.key_mem[9][94] ),
    .A2(_16535_),
    .B1(_16854_),
    .B2(\core.keymem.key_mem[1][94] ),
    .ZN(_03536_));
 AOI22_X1 _25877_ (.A1(\core.keymem.key_mem[2][94] ),
    .A2(_16859_),
    .B1(_16531_),
    .B2(\core.keymem.key_mem[13][94] ),
    .ZN(_03537_));
 NAND2_X1 _25878_ (.A1(_03536_),
    .A2(_03537_),
    .ZN(_03538_));
 NOR4_X4 _25879_ (.A1(_16546_),
    .A2(_03530_),
    .A3(_03535_),
    .A4(_03538_),
    .ZN(_03539_));
 AOI21_X4 _25880_ (.A(_03539_),
    .B1(_16547_),
    .B2(_00216_),
    .ZN(_03540_));
 XNOR2_X2 _25881_ (.A(\core.dec_block.block_w1_reg[30] ),
    .B(_03540_),
    .ZN(_03541_));
 XNOR2_X2 _25882_ (.A(_17169_),
    .B(_03541_),
    .ZN(_03542_));
 AOI22_X1 _25883_ (.A1(\core.keymem.key_mem[7][89] ),
    .A2(_17084_),
    .B1(_16529_),
    .B2(\core.keymem.key_mem[8][89] ),
    .ZN(_03543_));
 AOI22_X1 _25884_ (.A1(\core.keymem.key_mem[14][89] ),
    .A2(_17719_),
    .B1(_16860_),
    .B2(\core.keymem.key_mem[2][89] ),
    .ZN(_03544_));
 AOI22_X1 _25885_ (.A1(\core.keymem.key_mem[3][89] ),
    .A2(_16386_),
    .B1(_16515_),
    .B2(\core.keymem.key_mem[10][89] ),
    .ZN(_03545_));
 AOI21_X1 _25886_ (.A(_16982_),
    .B1(_16539_),
    .B2(\core.keymem.key_mem[12][89] ),
    .ZN(_03546_));
 NAND4_X1 _25887_ (.A1(_03543_),
    .A2(_03544_),
    .A3(_03545_),
    .A4(_03546_),
    .ZN(_03547_));
 MUX2_X1 _25888_ (.A(\core.keymem.key_mem[5][89] ),
    .B(\core.keymem.key_mem[13][89] ),
    .S(_17054_),
    .Z(_03548_));
 AOI22_X1 _25889_ (.A1(\core.keymem.key_mem[9][89] ),
    .A2(_17067_),
    .B1(_17051_),
    .B2(_03548_),
    .ZN(_03549_));
 NOR2_X1 _25890_ (.A1(_16880_),
    .A2(_03549_),
    .ZN(_03550_));
 AOI22_X1 _25891_ (.A1(\core.keymem.key_mem[4][89] ),
    .A2(_16457_),
    .B1(_16855_),
    .B2(\core.keymem.key_mem[1][89] ),
    .ZN(_03551_));
 AOI22_X1 _25892_ (.A1(\core.keymem.key_mem[6][89] ),
    .A2(_16448_),
    .B1(_16442_),
    .B2(\core.keymem.key_mem[11][89] ),
    .ZN(_03552_));
 NAND2_X1 _25893_ (.A1(_03551_),
    .A2(_03552_),
    .ZN(_03553_));
 NOR3_X2 _25894_ (.A1(_03547_),
    .A2(_03550_),
    .A3(_03553_),
    .ZN(_03554_));
 AOI21_X4 _25895_ (.A(_03554_),
    .B1(_16497_),
    .B2(_00229_),
    .ZN(_03555_));
 XNOR2_X2 _25896_ (.A(\core.dec_block.block_w1_reg[25] ),
    .B(_03555_),
    .ZN(_03556_));
 XNOR2_X1 _25897_ (.A(_03542_),
    .B(_03556_),
    .ZN(_03557_));
 XNOR2_X2 _25898_ (.A(_03527_),
    .B(_03557_),
    .ZN(_03558_));
 MUX2_X1 _25899_ (.A(\core.keymem.key_mem[3][73] ),
    .B(\core.keymem.key_mem[11][73] ),
    .S(_16972_),
    .Z(_03559_));
 NOR2_X1 _25900_ (.A1(_16378_),
    .A2(_16960_),
    .ZN(_03560_));
 AOI22_X2 _25901_ (.A1(\core.keymem.key_mem[14][73] ),
    .A2(_16436_),
    .B1(_03559_),
    .B2(_03560_),
    .ZN(_03561_));
 AOI22_X2 _25902_ (.A1(\core.keymem.key_mem[13][73] ),
    .A2(_16881_),
    .B1(_17067_),
    .B2(\core.keymem.key_mem[9][73] ),
    .ZN(_03562_));
 AOI222_X2 _25903_ (.A1(\core.keymem.key_mem[6][73] ),
    .A2(_16906_),
    .B1(_16964_),
    .B2(\core.keymem.key_mem[5][73] ),
    .C1(\core.keymem.key_mem[4][73] ),
    .C2(_16483_),
    .ZN(_03563_));
 OAI221_X2 _25904_ (.A(_03561_),
    .B1(_03562_),
    .B2(_16880_),
    .C1(_17042_),
    .C2(_03563_),
    .ZN(_03564_));
 AOI22_X1 _25905_ (.A1(\core.keymem.key_mem[2][73] ),
    .A2(_17025_),
    .B1(_16964_),
    .B2(\core.keymem.key_mem[1][73] ),
    .ZN(_03565_));
 NAND2_X1 _25906_ (.A1(_16902_),
    .A2(_03565_),
    .ZN(_03566_));
 NAND3_X1 _25907_ (.A1(\core.keymem.key_mem[8][73] ),
    .A2(_16484_),
    .A3(_16958_),
    .ZN(_03567_));
 AOI21_X1 _25908_ (.A(_16958_),
    .B1(_16481_),
    .B2(\core.keymem.key_mem[7][73] ),
    .ZN(_03568_));
 OAI21_X1 _25909_ (.A(_03567_),
    .B1(_03568_),
    .B2(_17054_),
    .ZN(_03569_));
 NAND3_X1 _25910_ (.A1(\core.keymem.key_mem[10][73] ),
    .A2(_16907_),
    .A3(_16958_),
    .ZN(_03570_));
 NAND3_X1 _25911_ (.A1(\core.keymem.key_mem[12][73] ),
    .A2(_16931_),
    .A3(_16961_),
    .ZN(_03571_));
 NAND2_X1 _25912_ (.A1(_03570_),
    .A2(_03571_),
    .ZN(_03572_));
 AOI221_X2 _25913_ (.A(_03564_),
    .B1(_03566_),
    .B2(_03569_),
    .C1(_03572_),
    .C2(_17055_),
    .ZN(_03573_));
 MUX2_X2 _25914_ (.A(_00234_),
    .B(_03573_),
    .S(_16488_),
    .Z(_03574_));
 XOR2_X2 _25915_ (.A(\core.dec_block.block_w1_reg[9] ),
    .B(_03574_),
    .Z(_03575_));
 XNOR2_X2 _25916_ (.A(_17062_),
    .B(_03575_),
    .ZN(_03576_));
 AOI222_X2 _25917_ (.A1(\core.keymem.key_mem[3][78] ),
    .A2(_16864_),
    .B1(_16460_),
    .B2(\core.keymem.key_mem[9][78] ),
    .C1(\core.keymem.key_mem[10][78] ),
    .C2(_16430_),
    .ZN(_03577_));
 AOI22_X1 _25918_ (.A1(\core.keymem.key_mem[4][78] ),
    .A2(_16946_),
    .B1(_16396_),
    .B2(\core.keymem.key_mem[12][78] ),
    .ZN(_03578_));
 AOI22_X1 _25919_ (.A1(\core.keymem.key_mem[6][78] ),
    .A2(_16447_),
    .B1(_16523_),
    .B2(\core.keymem.key_mem[1][78] ),
    .ZN(_03579_));
 AND3_X1 _25920_ (.A1(_03577_),
    .A2(_03578_),
    .A3(_03579_),
    .ZN(_03580_));
 INV_X1 _25921_ (.A(\core.keymem.key_mem[2][78] ),
    .ZN(_03581_));
 INV_X1 _25922_ (.A(\core.keymem.key_mem[8][78] ),
    .ZN(_03582_));
 OAI22_X4 _25923_ (.A1(_03581_),
    .A2(_17886_),
    .B1(_17134_),
    .B2(_03582_),
    .ZN(_03583_));
 INV_X1 _25924_ (.A(\core.keymem.key_mem[7][78] ),
    .ZN(_03584_));
 OAI21_X2 _25925_ (.A(_16481_),
    .B1(_16926_),
    .B2(_16928_),
    .ZN(_03585_));
 INV_X1 _25926_ (.A(\core.keymem.key_mem[11][78] ),
    .ZN(_03586_));
 OAI22_X4 _25927_ (.A1(_03584_),
    .A2(_18544_),
    .B1(_03585_),
    .B2(_03586_),
    .ZN(_03587_));
 NAND2_X1 _25928_ (.A1(\core.keymem.key_mem[14][78] ),
    .A2(_17025_),
    .ZN(_03588_));
 OAI21_X1 _25929_ (.A(\core.keymem.key_mem[13][78] ),
    .B1(_16912_),
    .B2(_16914_),
    .ZN(_03589_));
 AOI21_X2 _25930_ (.A(_16390_),
    .B1(_03588_),
    .B2(_03589_),
    .ZN(_03590_));
 OAI22_X4 _25931_ (.A1(_16895_),
    .A2(_16898_),
    .B1(_16912_),
    .B2(_16914_),
    .ZN(_03591_));
 INV_X1 _25932_ (.A(\core.keymem.key_mem[5][78] ),
    .ZN(_03592_));
 OAI21_X2 _25933_ (.A(_16486_),
    .B1(_03591_),
    .B2(_03592_),
    .ZN(_03593_));
 NOR4_X4 _25934_ (.A1(_03583_),
    .A2(_03587_),
    .A3(_03590_),
    .A4(_03593_),
    .ZN(_03594_));
 AOI22_X4 _25935_ (.A1(_00221_),
    .A2(_17013_),
    .B1(_03580_),
    .B2(_03594_),
    .ZN(_03595_));
 XNOR2_X2 _25936_ (.A(\core.dec_block.block_w1_reg[14] ),
    .B(_03595_),
    .ZN(_03596_));
 XNOR2_X2 _25937_ (.A(_03576_),
    .B(_03596_),
    .ZN(_03597_));
 INV_X1 _25938_ (.A(\core.dec_block.block_w1_reg[17] ),
    .ZN(_03598_));
 OAI211_X2 _25939_ (.A(\core.keymem.key_mem[4][81] ),
    .B(_16921_),
    .C1(_16933_),
    .C2(_16934_),
    .ZN(_03599_));
 OAI211_X2 _25940_ (.A(\core.keymem.key_mem[10][81] ),
    .B(_17025_),
    .C1(_16926_),
    .C2(_16928_),
    .ZN(_03600_));
 MUX2_X1 _25941_ (.A(\core.keymem.key_mem[3][81] ),
    .B(\core.keymem.key_mem[7][81] ),
    .S(_16960_),
    .Z(_03601_));
 NAND3_X1 _25942_ (.A1(_16938_),
    .A2(_16967_),
    .A3(_03601_),
    .ZN(_03602_));
 OAI221_X1 _25943_ (.A(\core.keymem.key_mem[9][81] ),
    .B1(_16884_),
    .B2(_16888_),
    .C1(_16912_),
    .C2(_16914_),
    .ZN(_03603_));
 AND4_X1 _25944_ (.A1(_03599_),
    .A2(_03600_),
    .A3(_03602_),
    .A4(_03603_),
    .ZN(_03604_));
 AOI22_X2 _25945_ (.A1(\core.keymem.key_mem[2][81] ),
    .A2(_17163_),
    .B1(_16964_),
    .B2(\core.keymem.key_mem[1][81] ),
    .ZN(_03605_));
 AOI22_X2 _25946_ (.A1(\core.keymem.key_mem[12][81] ),
    .A2(_16882_),
    .B1(_17067_),
    .B2(\core.keymem.key_mem[8][81] ),
    .ZN(_03606_));
 OAI221_X2 _25947_ (.A(_03604_),
    .B1(_03605_),
    .B2(_16383_),
    .C1(_03606_),
    .C2(_16394_),
    .ZN(_03607_));
 NAND3_X1 _25948_ (.A1(\core.keymem.key_mem[11][81] ),
    .A2(_17048_),
    .A3(_17043_),
    .ZN(_03608_));
 NAND2_X1 _25949_ (.A1(\core.keymem.key_mem[13][81] ),
    .A2(_16961_),
    .ZN(_03609_));
 OAI21_X1 _25950_ (.A(_03608_),
    .B1(_03609_),
    .B2(_16880_),
    .ZN(_03610_));
 NAND3_X1 _25951_ (.A1(\core.keymem.key_mem[14][81] ),
    .A2(_17050_),
    .A3(_17055_),
    .ZN(_03611_));
 AOI22_X1 _25952_ (.A1(\core.keymem.key_mem[6][81] ),
    .A2(_17016_),
    .B1(_16964_),
    .B2(\core.keymem.key_mem[5][81] ),
    .ZN(_03612_));
 OAI21_X1 _25953_ (.A(_03611_),
    .B1(_03612_),
    .B2(_17055_),
    .ZN(_03613_));
 AOI221_X2 _25954_ (.A(_03607_),
    .B1(_03610_),
    .B2(_17055_),
    .C1(_17051_),
    .C2(_03613_),
    .ZN(_03614_));
 MUX2_X2 _25955_ (.A(_00231_),
    .B(_03614_),
    .S(_16489_),
    .Z(_03615_));
 XNOR2_X2 _25956_ (.A(_03598_),
    .B(_03615_),
    .ZN(_03616_));
 AOI21_X1 _25957_ (.A(_16545_),
    .B1(_16949_),
    .B2(\core.keymem.key_mem[5][87] ),
    .ZN(_03617_));
 AOI22_X1 _25958_ (.A1(\core.keymem.key_mem[4][87] ),
    .A2(_16947_),
    .B1(_16998_),
    .B2(\core.keymem.key_mem[14][87] ),
    .ZN(_03618_));
 AOI22_X1 _25959_ (.A1(\core.keymem.key_mem[7][87] ),
    .A2(_17736_),
    .B1(_16520_),
    .B2(\core.keymem.key_mem[6][87] ),
    .ZN(_03619_));
 AOI22_X1 _25960_ (.A1(\core.keymem.key_mem[8][87] ),
    .A2(_17506_),
    .B1(_16416_),
    .B2(\core.keymem.key_mem[1][87] ),
    .ZN(_03620_));
 AND4_X1 _25961_ (.A1(_03617_),
    .A2(_03618_),
    .A3(_03619_),
    .A4(_03620_),
    .ZN(_03621_));
 AOI222_X2 _25962_ (.A1(\core.keymem.key_mem[3][87] ),
    .A2(_17175_),
    .B1(_16505_),
    .B2(\core.keymem.key_mem[11][87] ),
    .C1(\core.keymem.key_mem[13][87] ),
    .C2(_16531_),
    .ZN(_03622_));
 AOI22_X1 _25963_ (.A1(\core.keymem.key_mem[2][87] ),
    .A2(_16424_),
    .B1(_16432_),
    .B2(\core.keymem.key_mem[10][87] ),
    .ZN(_03623_));
 AOI22_X1 _25964_ (.A1(\core.keymem.key_mem[9][87] ),
    .A2(_16462_),
    .B1(_16398_),
    .B2(\core.keymem.key_mem[12][87] ),
    .ZN(_03624_));
 AND3_X1 _25965_ (.A1(_03622_),
    .A2(_03623_),
    .A3(_03624_),
    .ZN(_03625_));
 AOI22_X4 _25966_ (.A1(_00237_),
    .A2(_16852_),
    .B1(_03621_),
    .B2(_03625_),
    .ZN(_03626_));
 XNOR2_X2 _25967_ (.A(_18577_),
    .B(_03626_),
    .ZN(_03627_));
 XNOR2_X2 _25968_ (.A(_16943_),
    .B(_03627_),
    .ZN(_03628_));
 XOR2_X1 _25969_ (.A(_03616_),
    .B(_03628_),
    .Z(_03629_));
 XNOR2_X1 _25970_ (.A(_03597_),
    .B(_03629_),
    .ZN(_03630_));
 XNOR2_X2 _25971_ (.A(_03558_),
    .B(_03630_),
    .ZN(_03631_));
 AOI21_X1 _25972_ (.A(_03522_),
    .B1(_03631_),
    .B2(_18332_),
    .ZN(_03632_));
 AOI22_X1 _25973_ (.A1(_03365_),
    .A2(_17744_),
    .B1(_03498_),
    .B2(_03632_),
    .ZN(_00578_));
 NOR2_X1 _25974_ (.A1(\core.dec_block.block_w0_reg[20] ),
    .A2(_18330_),
    .ZN(_03633_));
 AOI21_X1 _25975_ (.A(_19358_),
    .B1(_18712_),
    .B2(_18745_),
    .ZN(_03634_));
 NAND2_X1 _25976_ (.A1(_18698_),
    .A2(_03634_),
    .ZN(_03635_));
 OAI21_X1 _25977_ (.A(_03635_),
    .B1(_19098_),
    .B2(_18698_),
    .ZN(_03636_));
 OAI221_X1 _25978_ (.A(_18788_),
    .B1(_18733_),
    .B2(_19314_),
    .C1(_03636_),
    .C2(_18716_),
    .ZN(_03637_));
 NAND2_X1 _25979_ (.A1(_18763_),
    .A2(_18668_),
    .ZN(_03638_));
 OAI33_X1 _25980_ (.A1(_18805_),
    .A2(_18744_),
    .A3(_18614_),
    .B1(_03638_),
    .B2(_18679_),
    .B3(_18646_),
    .ZN(_03639_));
 OAI21_X1 _25981_ (.A(_03637_),
    .B1(_03639_),
    .B2(_18789_),
    .ZN(_03640_));
 MUX2_X1 _25982_ (.A(_18647_),
    .B(_18652_),
    .S(_18816_),
    .Z(_03641_));
 NAND2_X1 _25983_ (.A1(_18703_),
    .A2(_03641_),
    .ZN(_03642_));
 AOI21_X1 _25984_ (.A(_18655_),
    .B1(_18801_),
    .B2(_19325_),
    .ZN(_03643_));
 AOI21_X1 _25985_ (.A(_03643_),
    .B1(_18652_),
    .B2(_18823_),
    .ZN(_03644_));
 OAI21_X2 _25986_ (.A(_03642_),
    .B1(_03644_),
    .B2(_19040_),
    .ZN(_03645_));
 AOI21_X2 _25987_ (.A(_18740_),
    .B1(_18760_),
    .B2(_19104_),
    .ZN(_03646_));
 AOI21_X1 _25988_ (.A(_03646_),
    .B1(_19134_),
    .B2(_19094_),
    .ZN(_03647_));
 NAND2_X1 _25989_ (.A1(_19160_),
    .A2(_19319_),
    .ZN(_03648_));
 NOR3_X1 _25990_ (.A1(_03645_),
    .A2(_03647_),
    .A3(_03648_),
    .ZN(_03649_));
 AOI21_X1 _25991_ (.A(_18635_),
    .B1(_18725_),
    .B2(_18738_),
    .ZN(_03650_));
 AOI21_X1 _25992_ (.A(_03650_),
    .B1(_18688_),
    .B2(_18695_),
    .ZN(_03651_));
 OAI221_X1 _25993_ (.A(_18817_),
    .B1(_19040_),
    .B2(_19496_),
    .C1(_03651_),
    .C2(_18629_),
    .ZN(_03652_));
 NOR3_X1 _25994_ (.A1(_18738_),
    .A2(_18648_),
    .A3(_18758_),
    .ZN(_03653_));
 AOI21_X1 _25995_ (.A(_03653_),
    .B1(_18768_),
    .B2(_18738_),
    .ZN(_03654_));
 OAI222_X2 _25996_ (.A1(_18722_),
    .A2(_18725_),
    .B1(_19115_),
    .B2(_18782_),
    .C1(_18805_),
    .C2(_03654_),
    .ZN(_03655_));
 OAI21_X1 _25997_ (.A(_03652_),
    .B1(_03655_),
    .B2(_18817_),
    .ZN(_03656_));
 NAND2_X1 _25998_ (.A1(_18715_),
    .A2(_18840_),
    .ZN(_03657_));
 OAI21_X1 _25999_ (.A(_18820_),
    .B1(_18744_),
    .B2(_18723_),
    .ZN(_03658_));
 NAND2_X1 _26000_ (.A1(_18805_),
    .A2(_03658_),
    .ZN(_03659_));
 AOI21_X1 _26001_ (.A(_18770_),
    .B1(_03657_),
    .B2(_03659_),
    .ZN(_03660_));
 NOR2_X1 _26002_ (.A1(_19149_),
    .A2(_03660_),
    .ZN(_03661_));
 AOI22_X2 _26003_ (.A1(_18765_),
    .A2(_19070_),
    .B1(_19355_),
    .B2(_18726_),
    .ZN(_03662_));
 OAI221_X2 _26004_ (.A(_03662_),
    .B1(_18749_),
    .B2(_18672_),
    .C1(_18665_),
    .C2(_19317_),
    .ZN(_03663_));
 NAND2_X1 _26005_ (.A1(_18763_),
    .A2(_18697_),
    .ZN(_03664_));
 OAI33_X1 _26006_ (.A1(_18698_),
    .A2(_18639_),
    .A3(_18672_),
    .B1(_03664_),
    .B2(_18651_),
    .B3(_18620_),
    .ZN(_03665_));
 AOI221_X2 _26007_ (.A(_03663_),
    .B1(_18845_),
    .B2(_18746_),
    .C1(_18816_),
    .C2(_03665_),
    .ZN(_03666_));
 AOI21_X1 _26008_ (.A(_18778_),
    .B1(_18764_),
    .B2(_18623_),
    .ZN(_03667_));
 OAI21_X1 _26009_ (.A(_18642_),
    .B1(_18596_),
    .B2(_18603_),
    .ZN(_03668_));
 MUX2_X1 _26010_ (.A(_18679_),
    .B(_03668_),
    .S(_18612_),
    .Z(_03669_));
 OAI33_X1 _26011_ (.A1(_18668_),
    .A2(_18670_),
    .A3(_03667_),
    .B1(_03669_),
    .B2(_18674_),
    .B3(_18678_),
    .ZN(_03670_));
 OR2_X1 _26012_ (.A1(_18794_),
    .A2(_18705_),
    .ZN(_03671_));
 OAI221_X2 _26013_ (.A(_03671_),
    .B1(_19164_),
    .B2(_19140_),
    .C1(_18672_),
    .C2(_19150_),
    .ZN(_03672_));
 NOR2_X1 _26014_ (.A1(_18573_),
    .A2(_18728_),
    .ZN(_03673_));
 NOR2_X1 _26015_ (.A1(_18661_),
    .A2(_18680_),
    .ZN(_03674_));
 OAI33_X1 _26016_ (.A1(_18624_),
    .A2(_18598_),
    .A3(_03673_),
    .B1(_03674_),
    .B2(_18614_),
    .B3(_18670_),
    .ZN(_03675_));
 NOR3_X1 _26017_ (.A1(_03670_),
    .A2(_03672_),
    .A3(_03675_),
    .ZN(_03676_));
 OAI21_X1 _26018_ (.A(_19168_),
    .B1(_18810_),
    .B2(_18796_),
    .ZN(_03677_));
 NAND3_X1 _26019_ (.A1(_18698_),
    .A2(_18688_),
    .A3(_03677_),
    .ZN(_03678_));
 OAI21_X1 _26020_ (.A(_18653_),
    .B1(_18793_),
    .B2(_19322_),
    .ZN(_03679_));
 AOI21_X1 _26021_ (.A(_18793_),
    .B1(_18653_),
    .B2(_18763_),
    .ZN(_03680_));
 OAI21_X1 _26022_ (.A(_03679_),
    .B1(_03680_),
    .B2(_18620_),
    .ZN(_03681_));
 NAND2_X1 _26023_ (.A1(_18842_),
    .A2(_03681_),
    .ZN(_03682_));
 NAND4_X1 _26024_ (.A1(_19054_),
    .A2(_03676_),
    .A3(_03678_),
    .A4(_03682_),
    .ZN(_03683_));
 NOR3_X1 _26025_ (.A1(_18748_),
    .A2(_19466_),
    .A3(_03683_),
    .ZN(_03684_));
 NAND4_X2 _26026_ (.A1(_03656_),
    .A2(_03661_),
    .A3(_03666_),
    .A4(_03684_),
    .ZN(_03685_));
 NOR2_X1 _26027_ (.A1(_18653_),
    .A2(_18639_),
    .ZN(_03686_));
 AOI21_X1 _26028_ (.A(_18715_),
    .B1(_18770_),
    .B2(_19131_),
    .ZN(_03687_));
 AOI221_X1 _26029_ (.A(_18698_),
    .B1(_18842_),
    .B2(_03686_),
    .C1(_03687_),
    .C2(_18783_),
    .ZN(_03688_));
 OAI21_X1 _26030_ (.A(_18738_),
    .B1(_18745_),
    .B2(_18758_),
    .ZN(_03689_));
 OAI21_X1 _26031_ (.A(_18715_),
    .B1(_19334_),
    .B2(_03689_),
    .ZN(_03690_));
 NOR2_X1 _26032_ (.A1(_18765_),
    .A2(_19098_),
    .ZN(_03691_));
 OAI22_X1 _26033_ (.A1(_19094_),
    .A2(_18770_),
    .B1(_03690_),
    .B2(_03691_),
    .ZN(_03692_));
 OAI21_X1 _26034_ (.A(_03690_),
    .B1(_18766_),
    .B2(_18808_),
    .ZN(_03693_));
 AOI21_X1 _26035_ (.A(_03692_),
    .B1(_03693_),
    .B2(_18659_),
    .ZN(_03694_));
 AOI21_X1 _26036_ (.A(_03688_),
    .B1(_03694_),
    .B2(_18700_),
    .ZN(_03695_));
 NOR2_X1 _26037_ (.A1(_03685_),
    .A2(_03695_),
    .ZN(_03696_));
 NAND4_X2 _26038_ (.A1(_19344_),
    .A2(_03640_),
    .A3(_03649_),
    .A4(_03696_),
    .ZN(_03697_));
 OAI21_X4 _26039_ (.A(_18416_),
    .B1(_19107_),
    .B2(_03697_),
    .ZN(_03698_));
 INV_X1 _26040_ (.A(\block_reg[3][20] ),
    .ZN(_03699_));
 NAND2_X1 _26041_ (.A1(_00286_),
    .A2(_16852_),
    .ZN(_03700_));
 AOI22_X1 _26042_ (.A1(\core.keymem.key_mem[8][20] ),
    .A2(_17506_),
    .B1(_16988_),
    .B2(\core.keymem.key_mem[10][20] ),
    .ZN(_03701_));
 AOI22_X1 _26043_ (.A1(\core.keymem.key_mem[7][20] ),
    .A2(_17736_),
    .B1(_16859_),
    .B2(\core.keymem.key_mem[2][20] ),
    .ZN(_03702_));
 AOI22_X1 _26044_ (.A1(\core.keymem.key_mem[3][20] ),
    .A2(_16986_),
    .B1(_16854_),
    .B2(\core.keymem.key_mem[1][20] ),
    .ZN(_03703_));
 AOI22_X1 _26045_ (.A1(\core.keymem.key_mem[6][20] ),
    .A2(_17648_),
    .B1(_16467_),
    .B2(\core.keymem.key_mem[5][20] ),
    .ZN(_03704_));
 AND4_X1 _26046_ (.A1(_03701_),
    .A2(_03702_),
    .A3(_03703_),
    .A4(_03704_),
    .ZN(_03705_));
 AOI22_X2 _26047_ (.A1(\core.keymem.key_mem[9][20] ),
    .A2(_17914_),
    .B1(_17720_),
    .B2(\core.keymem.key_mem[12][20] ),
    .ZN(_03706_));
 AOI22_X2 _26048_ (.A1(\core.keymem.key_mem[4][20] ),
    .A2(_16500_),
    .B1(_17008_),
    .B2(\core.keymem.key_mem[11][20] ),
    .ZN(_03707_));
 AOI22_X4 _26049_ (.A1(\core.keymem.key_mem[14][20] ),
    .A2(_16999_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][20] ),
    .ZN(_03708_));
 NAND4_X4 _26050_ (.A1(_03705_),
    .A2(_03706_),
    .A3(_03707_),
    .A4(_03708_),
    .ZN(_03709_));
 OAI21_X4 _26051_ (.A(_03700_),
    .B1(_03709_),
    .B2(_16547_),
    .ZN(_03710_));
 XNOR2_X1 _26052_ (.A(_03699_),
    .B(_03710_),
    .ZN(_03711_));
 AOI222_X2 _26053_ (.A1(\core.keymem.key_mem[14][116] ),
    .A2(_17581_),
    .B1(_17086_),
    .B2(\core.keymem.key_mem[2][116] ),
    .C1(_17771_),
    .C2(\core.keymem.key_mem[13][116] ),
    .ZN(_03712_));
 AOI22_X2 _26054_ (.A1(\core.keymem.key_mem[6][116] ),
    .A2(_16522_),
    .B1(_17765_),
    .B2(\core.keymem.key_mem[8][116] ),
    .ZN(_03713_));
 AOI22_X2 _26055_ (.A1(\core.keymem.key_mem[10][116] ),
    .A2(_17082_),
    .B1(_17769_),
    .B2(\core.keymem.key_mem[11][116] ),
    .ZN(_03714_));
 NAND3_X2 _26056_ (.A1(_03712_),
    .A2(_03713_),
    .A3(_03714_),
    .ZN(_03715_));
 AOI22_X1 _26057_ (.A1(\core.keymem.key_mem[12][116] ),
    .A2(_17093_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][116] ),
    .ZN(_03716_));
 AOI22_X2 _26058_ (.A1(\core.keymem.key_mem[4][116] ),
    .A2(_16501_),
    .B1(_16510_),
    .B2(\core.keymem.key_mem[5][116] ),
    .ZN(_03717_));
 AOI22_X2 _26059_ (.A1(\core.keymem.key_mem[3][116] ),
    .A2(_17091_),
    .B1(_17585_),
    .B2(\core.keymem.key_mem[9][116] ),
    .ZN(_03718_));
 AOI21_X2 _26060_ (.A(_16547_),
    .B1(_17085_),
    .B2(\core.keymem.key_mem[7][116] ),
    .ZN(_03719_));
 NAND4_X2 _26061_ (.A1(_03716_),
    .A2(_03717_),
    .A3(_03718_),
    .A4(_03719_),
    .ZN(_03720_));
 NOR2_X4 _26062_ (.A1(_03715_),
    .A2(_03720_),
    .ZN(_03721_));
 AND2_X2 _26063_ (.A1(_00208_),
    .A2(_16498_),
    .ZN(_03722_));
 NOR2_X4 _26064_ (.A1(_03721_),
    .A2(_03722_),
    .ZN(_03723_));
 XNOR2_X2 _26065_ (.A(\core.dec_block.block_w0_reg[20] ),
    .B(_03723_),
    .ZN(_03724_));
 OAI221_X2 _26066_ (.A(_18329_),
    .B1(_18466_),
    .B2(_03711_),
    .C1(_03724_),
    .C2(_18479_),
    .ZN(_03725_));
 XNOR2_X1 _26067_ (.A(_19247_),
    .B(_03304_),
    .ZN(_03726_));
 XNOR2_X2 _26068_ (.A(_18923_),
    .B(_03726_),
    .ZN(_03727_));
 AOI222_X2 _26069_ (.A1(\core.keymem.key_mem[6][28] ),
    .A2(_17648_),
    .B1(_16854_),
    .B2(\core.keymem.key_mem[1][28] ),
    .C1(_16531_),
    .C2(\core.keymem.key_mem[13][28] ),
    .ZN(_03728_));
 AOI22_X2 _26070_ (.A1(\core.keymem.key_mem[9][28] ),
    .A2(_17522_),
    .B1(_16432_),
    .B2(\core.keymem.key_mem[10][28] ),
    .ZN(_03729_));
 AOI22_X2 _26071_ (.A1(\core.keymem.key_mem[12][28] ),
    .A2(_17000_),
    .B1(_17007_),
    .B2(\core.keymem.key_mem[11][28] ),
    .ZN(_03730_));
 NAND3_X2 _26072_ (.A1(_03728_),
    .A2(_03729_),
    .A3(_03730_),
    .ZN(_03731_));
 AOI22_X2 _26073_ (.A1(\core.keymem.key_mem[14][28] ),
    .A2(_16998_),
    .B1(_16986_),
    .B2(\core.keymem.key_mem[3][28] ),
    .ZN(_03732_));
 AOI22_X2 _26074_ (.A1(\core.keymem.key_mem[2][28] ),
    .A2(_16993_),
    .B1(_16528_),
    .B2(\core.keymem.key_mem[8][28] ),
    .ZN(_03733_));
 AOI22_X2 _26075_ (.A1(\core.keymem.key_mem[7][28] ),
    .A2(_17736_),
    .B1(_16467_),
    .B2(\core.keymem.key_mem[5][28] ),
    .ZN(_03734_));
 AOI21_X1 _26076_ (.A(_16494_),
    .B1(_16499_),
    .B2(\core.keymem.key_mem[4][28] ),
    .ZN(_03735_));
 NAND4_X2 _26077_ (.A1(_03732_),
    .A2(_03733_),
    .A3(_03734_),
    .A4(_03735_),
    .ZN(_03736_));
 NOR2_X4 _26078_ (.A1(_03731_),
    .A2(_03736_),
    .ZN(_03737_));
 AOI21_X4 _26079_ (.A(_03737_),
    .B1(_16872_),
    .B2(_00301_),
    .ZN(_03738_));
 XNOR2_X2 _26080_ (.A(\core.dec_block.block_w3_reg[28] ),
    .B(_03738_),
    .ZN(_03739_));
 XNOR2_X1 _26081_ (.A(_19299_),
    .B(_03739_),
    .ZN(_03740_));
 XNOR2_X1 _26082_ (.A(_03727_),
    .B(_03740_),
    .ZN(_03741_));
 XNOR2_X2 _26083_ (.A(_19260_),
    .B(_19458_),
    .ZN(_03742_));
 XNOR2_X2 _26084_ (.A(_18884_),
    .B(_03742_),
    .ZN(_03743_));
 XNOR2_X1 _26085_ (.A(_18921_),
    .B(_19274_),
    .ZN(_03744_));
 XNOR2_X1 _26086_ (.A(_03333_),
    .B(_03744_),
    .ZN(_03745_));
 XOR2_X1 _26087_ (.A(_03743_),
    .B(_03745_),
    .Z(_03746_));
 XNOR2_X1 _26088_ (.A(_03741_),
    .B(_03746_),
    .ZN(_03747_));
 AOI222_X2 _26089_ (.A1(\core.keymem.key_mem[14][4] ),
    .A2(_17719_),
    .B1(_16424_),
    .B2(\core.keymem.key_mem[2][4] ),
    .C1(_16452_),
    .C2(\core.keymem.key_mem[8][4] ),
    .ZN(_03748_));
 AOI22_X2 _26090_ (.A1(\core.keymem.key_mem[1][4] ),
    .A2(_17003_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][4] ),
    .ZN(_03749_));
 AOI22_X2 _26091_ (.A1(\core.keymem.key_mem[9][4] ),
    .A2(_17914_),
    .B1(_17008_),
    .B2(\core.keymem.key_mem[11][4] ),
    .ZN(_03750_));
 NAND3_X2 _26092_ (.A1(_03748_),
    .A2(_03749_),
    .A3(_03750_),
    .ZN(_03751_));
 AOI22_X2 _26093_ (.A1(\core.keymem.key_mem[10][4] ),
    .A2(_16989_),
    .B1(_17720_),
    .B2(\core.keymem.key_mem[12][4] ),
    .ZN(_03752_));
 AOI22_X2 _26094_ (.A1(\core.keymem.key_mem[6][4] ),
    .A2(_17695_),
    .B1(_16866_),
    .B2(\core.keymem.key_mem[3][4] ),
    .ZN(_03753_));
 AOI22_X2 _26095_ (.A1(\core.keymem.key_mem[7][4] ),
    .A2(_17084_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][4] ),
    .ZN(_03754_));
 AOI21_X1 _26096_ (.A(_16495_),
    .B1(_17713_),
    .B2(\core.keymem.key_mem[4][4] ),
    .ZN(_03755_));
 NAND4_X2 _26097_ (.A1(_03752_),
    .A2(_03753_),
    .A3(_03754_),
    .A4(_03755_),
    .ZN(_03756_));
 NOR2_X4 _26098_ (.A1(_03751_),
    .A2(_03756_),
    .ZN(_03757_));
 AND2_X2 _26099_ (.A1(_00206_),
    .A2(_17014_),
    .ZN(_03758_));
 NOR2_X4 _26100_ (.A1(_03757_),
    .A2(_03758_),
    .ZN(_03759_));
 XNOR2_X2 _26101_ (.A(\core.dec_block.block_w3_reg[4] ),
    .B(_03759_),
    .ZN(_03760_));
 XNOR2_X2 _26102_ (.A(_19225_),
    .B(_03760_),
    .ZN(_03761_));
 XNOR2_X2 _26103_ (.A(\core.dec_block.block_w3_reg[19] ),
    .B(_03298_),
    .ZN(_03762_));
 XNOR2_X2 _26104_ (.A(_18956_),
    .B(_03762_),
    .ZN(_03763_));
 NAND2_X1 _26105_ (.A1(_00246_),
    .A2(_17183_),
    .ZN(_03764_));
 AOI22_X1 _26106_ (.A1(\core.keymem.key_mem[10][12] ),
    .A2(_17715_),
    .B1(_16532_),
    .B2(\core.keymem.key_mem[13][12] ),
    .ZN(_03765_));
 AOI22_X1 _26107_ (.A1(\core.keymem.key_mem[9][12] ),
    .A2(_16462_),
    .B1(_16416_),
    .B2(\core.keymem.key_mem[1][12] ),
    .ZN(_03766_));
 AOI22_X1 _26108_ (.A1(\core.keymem.key_mem[4][12] ),
    .A2(_16947_),
    .B1(_16407_),
    .B2(\core.keymem.key_mem[7][12] ),
    .ZN(_03767_));
 AOI22_X1 _26109_ (.A1(\core.keymem.key_mem[14][12] ),
    .A2(_16438_),
    .B1(_16386_),
    .B2(\core.keymem.key_mem[3][12] ),
    .ZN(_03768_));
 AND4_X1 _26110_ (.A1(_03765_),
    .A2(_03766_),
    .A3(_03767_),
    .A4(_03768_),
    .ZN(_03769_));
 AOI22_X2 _26111_ (.A1(\core.keymem.key_mem[6][12] ),
    .A2(_16449_),
    .B1(_16443_),
    .B2(\core.keymem.key_mem[11][12] ),
    .ZN(_03770_));
 AOI22_X2 _26112_ (.A1(\core.keymem.key_mem[2][12] ),
    .A2(_16425_),
    .B1(_16469_),
    .B2(\core.keymem.key_mem[5][12] ),
    .ZN(_03771_));
 AOI22_X2 _26113_ (.A1(\core.keymem.key_mem[8][12] ),
    .A2(_16530_),
    .B1(_16540_),
    .B2(\core.keymem.key_mem[12][12] ),
    .ZN(_03772_));
 NAND4_X4 _26114_ (.A1(_03769_),
    .A2(_03770_),
    .A3(_03771_),
    .A4(_03772_),
    .ZN(_03773_));
 OAI21_X4 _26115_ (.A(_03764_),
    .B1(_03773_),
    .B2(_16873_),
    .ZN(_03774_));
 XOR2_X2 _26116_ (.A(\core.dec_block.block_w3_reg[12] ),
    .B(_03774_),
    .Z(_03775_));
 XNOR2_X2 _26117_ (.A(_18942_),
    .B(_03344_),
    .ZN(_03776_));
 XNOR2_X1 _26118_ (.A(_03775_),
    .B(_03776_),
    .ZN(_03777_));
 XNOR2_X1 _26119_ (.A(_03763_),
    .B(_03777_),
    .ZN(_03778_));
 XNOR2_X1 _26120_ (.A(_03761_),
    .B(_03778_),
    .ZN(_03779_));
 XNOR2_X1 _26121_ (.A(_03747_),
    .B(_03779_),
    .ZN(_03780_));
 AOI21_X1 _26122_ (.A(_03725_),
    .B1(_03780_),
    .B2(_19031_),
    .ZN(_03781_));
 AOI21_X1 _26123_ (.A(_03633_),
    .B1(_03698_),
    .B2(_03781_),
    .ZN(_00579_));
 NOR2_X1 _26124_ (.A1(\core.dec_block.block_w0_reg[21] ),
    .A2(_18330_),
    .ZN(_03782_));
 XNOR2_X2 _26125_ (.A(_19260_),
    .B(_03358_),
    .ZN(_03783_));
 XOR2_X2 _26126_ (.A(_19442_),
    .B(_03783_),
    .Z(_03784_));
 XNOR2_X1 _26127_ (.A(_19002_),
    .B(_03762_),
    .ZN(_03785_));
 XNOR2_X1 _26128_ (.A(_18921_),
    .B(_03332_),
    .ZN(_03786_));
 XNOR2_X1 _26129_ (.A(_03785_),
    .B(_03786_),
    .ZN(_03787_));
 XNOR2_X1 _26130_ (.A(_03784_),
    .B(_03787_),
    .ZN(_03788_));
 XNOR2_X2 _26131_ (.A(_18970_),
    .B(_19414_),
    .ZN(_03789_));
 XOR2_X2 _26132_ (.A(\core.dec_block.block_w3_reg[20] ),
    .B(_03710_),
    .Z(_03790_));
 XNOR2_X2 _26133_ (.A(_18897_),
    .B(_03742_),
    .ZN(_03791_));
 XNOR2_X1 _26134_ (.A(_03790_),
    .B(_03791_),
    .ZN(_03792_));
 XNOR2_X2 _26135_ (.A(_03789_),
    .B(_03792_),
    .ZN(_03793_));
 XNOR2_X1 _26136_ (.A(_03788_),
    .B(_03793_),
    .ZN(_03794_));
 XNOR2_X1 _26137_ (.A(_03775_),
    .B(_03794_),
    .ZN(_03795_));
 NAND2_X1 _26138_ (.A1(_18333_),
    .A2(_03795_),
    .ZN(_03796_));
 OAI221_X2 _26139_ (.A(_18789_),
    .B1(_18676_),
    .B2(_19094_),
    .C1(_18769_),
    .C2(_18694_),
    .ZN(_03797_));
 OAI33_X1 _26140_ (.A1(_18700_),
    .A2(_19314_),
    .A3(_19134_),
    .B1(_19322_),
    .B2(_18598_),
    .B3(_18817_),
    .ZN(_03798_));
 OAI21_X1 _26141_ (.A(_03797_),
    .B1(_03798_),
    .B2(_18789_),
    .ZN(_03799_));
 NAND3_X1 _26142_ (.A1(_18788_),
    .A2(_18744_),
    .A3(_18672_),
    .ZN(_03800_));
 OAI21_X1 _26143_ (.A(_03800_),
    .B1(_18708_),
    .B2(_18788_),
    .ZN(_03801_));
 OAI21_X1 _26144_ (.A(_19043_),
    .B1(_03801_),
    .B2(_19314_),
    .ZN(_03802_));
 NOR2_X1 _26145_ (.A1(_19176_),
    .A2(_03802_),
    .ZN(_03803_));
 NAND3_X1 _26146_ (.A1(_18788_),
    .A2(_18699_),
    .A3(_18711_),
    .ZN(_03804_));
 NAND3_X1 _26147_ (.A1(_18832_),
    .A2(_18609_),
    .A3(_18768_),
    .ZN(_03805_));
 AOI21_X1 _26148_ (.A(_18716_),
    .B1(_03804_),
    .B2(_03805_),
    .ZN(_03806_));
 OAI22_X1 _26149_ (.A1(_18696_),
    .A2(_18705_),
    .B1(_19144_),
    .B2(_18744_),
    .ZN(_03807_));
 OAI21_X1 _26150_ (.A(_18722_),
    .B1(_18796_),
    .B2(_18665_),
    .ZN(_03808_));
 OAI21_X1 _26151_ (.A(_19134_),
    .B1(_18676_),
    .B2(_18665_),
    .ZN(_03809_));
 AOI22_X1 _26152_ (.A1(_19142_),
    .A2(_03808_),
    .B1(_03809_),
    .B2(_18703_),
    .ZN(_03810_));
 NOR3_X1 _26153_ (.A1(_18741_),
    .A2(_18670_),
    .A3(_18736_),
    .ZN(_03811_));
 AOI21_X1 _26154_ (.A(_03811_),
    .B1(_19307_),
    .B2(_18793_),
    .ZN(_03812_));
 OAI21_X1 _26155_ (.A(_03810_),
    .B1(_03812_),
    .B2(_18635_),
    .ZN(_03813_));
 NOR4_X1 _26156_ (.A1(_18724_),
    .A2(_03806_),
    .A3(_03807_),
    .A4(_03813_),
    .ZN(_03814_));
 OAI22_X1 _26157_ (.A1(_18710_),
    .A2(_19363_),
    .B1(_19317_),
    .B2(_18631_),
    .ZN(_03815_));
 AOI21_X1 _26158_ (.A(_19469_),
    .B1(_03815_),
    .B2(_18650_),
    .ZN(_03816_));
 NOR2_X1 _26159_ (.A1(_18653_),
    .A2(_18819_),
    .ZN(_03817_));
 AOI21_X1 _26160_ (.A(_03817_),
    .B1(_19322_),
    .B2(_18768_),
    .ZN(_03818_));
 NOR2_X1 _26161_ (.A1(_18832_),
    .A2(_03818_),
    .ZN(_03819_));
 OAI21_X1 _26162_ (.A(_18726_),
    .B1(_18677_),
    .B2(_18682_),
    .ZN(_03820_));
 OAI221_X2 _26163_ (.A(_03820_),
    .B1(_19135_),
    .B2(_18733_),
    .C1(_18666_),
    .C2(_18705_),
    .ZN(_03821_));
 AOI21_X1 _26164_ (.A(_18765_),
    .B1(_19104_),
    .B2(_18668_),
    .ZN(_03822_));
 OAI22_X2 _26165_ (.A1(_19094_),
    .A2(_19136_),
    .B1(_03822_),
    .B2(_19052_),
    .ZN(_03823_));
 NOR4_X1 _26166_ (.A1(_18734_),
    .A2(_03819_),
    .A3(_03821_),
    .A4(_03823_),
    .ZN(_03824_));
 AND4_X1 _26167_ (.A1(_03803_),
    .A2(_03814_),
    .A3(_03816_),
    .A4(_03824_),
    .ZN(_03825_));
 OAI21_X1 _26168_ (.A(_18699_),
    .B1(_18651_),
    .B2(_18808_),
    .ZN(_03826_));
 OAI221_X1 _26169_ (.A(_18815_),
    .B1(_18699_),
    .B2(_18712_),
    .C1(_19334_),
    .C2(_03826_),
    .ZN(_03827_));
 OAI21_X1 _26170_ (.A(_18719_),
    .B1(_18681_),
    .B2(_18832_),
    .ZN(_03828_));
 AOI22_X1 _26171_ (.A1(_18789_),
    .A2(_19155_),
    .B1(_18680_),
    .B2(_03828_),
    .ZN(_03829_));
 OAI21_X1 _26172_ (.A(_03827_),
    .B1(_03829_),
    .B2(_18716_),
    .ZN(_03830_));
 OAI21_X1 _26173_ (.A(_18746_),
    .B1(_19098_),
    .B2(_03817_),
    .ZN(_03831_));
 MUX2_X1 _26174_ (.A(_18573_),
    .B(_19481_),
    .S(_18750_),
    .Z(_03832_));
 NOR3_X1 _26175_ (.A1(_18738_),
    .A2(_18741_),
    .A3(_03832_),
    .ZN(_03833_));
 XNOR2_X1 _26176_ (.A(_18626_),
    .B(_18750_),
    .ZN(_03834_));
 NOR3_X1 _26177_ (.A1(_18621_),
    .A2(_18629_),
    .A3(_03834_),
    .ZN(_03835_));
 OAI21_X1 _26178_ (.A(_18634_),
    .B1(_03833_),
    .B2(_03835_),
    .ZN(_03836_));
 NAND4_X1 _26179_ (.A1(_18621_),
    .A2(_18805_),
    .A3(_18654_),
    .A4(_18780_),
    .ZN(_03837_));
 OAI21_X1 _26180_ (.A(_19076_),
    .B1(_18744_),
    .B2(_18715_),
    .ZN(_03838_));
 NAND3_X1 _26181_ (.A1(_18832_),
    .A2(_18816_),
    .A3(_03838_),
    .ZN(_03839_));
 NAND4_X1 _26182_ (.A1(_03831_),
    .A2(_03836_),
    .A3(_03837_),
    .A4(_03839_),
    .ZN(_03840_));
 MUX2_X1 _26183_ (.A(_18665_),
    .B(_18743_),
    .S(_18620_),
    .Z(_03841_));
 OAI22_X1 _26184_ (.A1(_19040_),
    .A2(_18733_),
    .B1(_03841_),
    .B2(_19481_),
    .ZN(_03842_));
 MUX2_X1 _26185_ (.A(_03840_),
    .B(_03842_),
    .S(_18700_),
    .Z(_03843_));
 NOR3_X2 _26186_ (.A1(_03645_),
    .A2(_03830_),
    .A3(_03843_),
    .ZN(_03844_));
 NAND4_X4 _26187_ (.A1(_19369_),
    .A2(_03799_),
    .A3(_03825_),
    .A4(_03844_),
    .ZN(_03845_));
 XNOR2_X1 _26188_ (.A(\block_reg[3][21] ),
    .B(_18908_),
    .ZN(_03846_));
 AOI22_X1 _26189_ (.A1(\core.keymem.key_mem[10][117] ),
    .A2(_16430_),
    .B1(_16414_),
    .B2(\core.keymem.key_mem[1][117] ),
    .ZN(_03847_));
 AOI21_X1 _26190_ (.A(_16493_),
    .B1(_16405_),
    .B2(\core.keymem.key_mem[7][117] ),
    .ZN(_03848_));
 AOI22_X1 _26191_ (.A1(\core.keymem.key_mem[3][117] ),
    .A2(_16384_),
    .B1(_16460_),
    .B2(\core.keymem.key_mem[9][117] ),
    .ZN(_03849_));
 AOI22_X2 _26192_ (.A1(\core.keymem.key_mem[14][117] ),
    .A2(_16435_),
    .B1(_16395_),
    .B2(\core.keymem.key_mem[12][117] ),
    .ZN(_03850_));
 AND4_X2 _26193_ (.A1(_03847_),
    .A2(_03848_),
    .A3(_03849_),
    .A4(_03850_),
    .ZN(_03851_));
 AOI222_X2 _26194_ (.A1(\core.keymem.key_mem[6][117] ),
    .A2(_16446_),
    .B1(_16422_),
    .B2(\core.keymem.key_mem[2][117] ),
    .C1(_16450_),
    .C2(\core.keymem.key_mem[8][117] ),
    .ZN(_03852_));
 AOI22_X1 _26195_ (.A1(\core.keymem.key_mem[11][117] ),
    .A2(_16504_),
    .B1(_16470_),
    .B2(\core.keymem.key_mem[13][117] ),
    .ZN(_03853_));
 AOI22_X1 _26196_ (.A1(\core.keymem.key_mem[4][117] ),
    .A2(_16455_),
    .B1(_16466_),
    .B2(\core.keymem.key_mem[5][117] ),
    .ZN(_03854_));
 AND3_X2 _26197_ (.A1(_03852_),
    .A2(_03853_),
    .A3(_03854_),
    .ZN(_03855_));
 AOI22_X4 _26198_ (.A1(_00178_),
    .A2(_16545_),
    .B1(_03851_),
    .B2(_03855_),
    .ZN(_03856_));
 XNOR2_X2 _26199_ (.A(\core.dec_block.block_w0_reg[21] ),
    .B(_03856_),
    .ZN(_03857_));
 BUF_X4 _26200_ (.A(_16555_),
    .Z(_03858_));
 OAI221_X2 _26201_ (.A(_18329_),
    .B1(_18553_),
    .B2(_03846_),
    .C1(_03857_),
    .C2(_03858_),
    .ZN(_03859_));
 NOR2_X1 _26202_ (.A1(_03845_),
    .A2(_03859_),
    .ZN(_03860_));
 AOI21_X1 _26203_ (.A(_03782_),
    .B1(_03796_),
    .B2(_03860_),
    .ZN(_00580_));
 NOR2_X1 _26204_ (.A1(\core.dec_block.block_w0_reg[22] ),
    .A2(_18330_),
    .ZN(_03861_));
 NOR3_X1 _26205_ (.A1(_18808_),
    .A2(_18723_),
    .A3(_18820_),
    .ZN(_03862_));
 AOI21_X1 _26206_ (.A(_03862_),
    .B1(_19490_),
    .B2(_18817_),
    .ZN(_03863_));
 MUX2_X1 _26207_ (.A(_18723_),
    .B(_18668_),
    .S(_18738_),
    .Z(_03864_));
 AOI21_X1 _26208_ (.A(_18803_),
    .B1(_03864_),
    .B2(_18647_),
    .ZN(_03865_));
 OAI22_X1 _26209_ (.A1(_18782_),
    .A2(_03863_),
    .B1(_03865_),
    .B2(_18716_),
    .ZN(_03866_));
 NOR3_X1 _26210_ (.A1(_18658_),
    .A2(_18816_),
    .A3(_19347_),
    .ZN(_03867_));
 NAND2_X1 _26211_ (.A1(_18774_),
    .A2(_19358_),
    .ZN(_03868_));
 OAI21_X1 _26212_ (.A(_19135_),
    .B1(_19144_),
    .B2(_18743_),
    .ZN(_03869_));
 OAI21_X1 _26213_ (.A(_03869_),
    .B1(_18768_),
    .B2(_18686_),
    .ZN(_03870_));
 AOI222_X2 _26214_ (.A1(_18628_),
    .A2(_18842_),
    .B1(_18726_),
    .B2(_19053_),
    .C1(_18682_),
    .C2(_18779_),
    .ZN(_03871_));
 NAND3_X1 _26215_ (.A1(_03868_),
    .A2(_03870_),
    .A3(_03871_),
    .ZN(_03872_));
 OR4_X1 _26216_ (.A1(_19330_),
    .A2(_03867_),
    .A3(_19505_),
    .A4(_03872_),
    .ZN(_03873_));
 NOR4_X1 _26217_ (.A1(_18813_),
    .A2(_03823_),
    .A3(_03866_),
    .A4(_03873_),
    .ZN(_03874_));
 NAND2_X1 _26218_ (.A1(_19102_),
    .A2(_03874_),
    .ZN(_03875_));
 OAI33_X1 _26219_ (.A1(_18782_),
    .A2(_18684_),
    .A3(_18706_),
    .B1(_18681_),
    .B2(_18758_),
    .B3(_18621_),
    .ZN(_03876_));
 OAI21_X1 _26220_ (.A(_18776_),
    .B1(_18749_),
    .B2(_18598_),
    .ZN(_03877_));
 NAND2_X1 _26221_ (.A1(_18820_),
    .A2(_18598_),
    .ZN(_03878_));
 NOR2_X1 _26222_ (.A1(_18581_),
    .A2(_18640_),
    .ZN(_03879_));
 OAI21_X1 _26223_ (.A(_18633_),
    .B1(_18653_),
    .B2(_18697_),
    .ZN(_03880_));
 OAI21_X1 _26224_ (.A(_03880_),
    .B1(_18694_),
    .B2(_18750_),
    .ZN(_03881_));
 NOR2_X1 _26225_ (.A1(_18631_),
    .A2(_18654_),
    .ZN(_03882_));
 OAI33_X1 _26226_ (.A1(_18643_),
    .A2(_18585_),
    .A3(_18655_),
    .B1(_03881_),
    .B2(_03882_),
    .B3(_18741_),
    .ZN(_03883_));
 AOI221_X2 _26227_ (.A(_03876_),
    .B1(_03877_),
    .B2(_03878_),
    .C1(_03879_),
    .C2(_03883_),
    .ZN(_03884_));
 INV_X1 _26228_ (.A(_03640_),
    .ZN(_03885_));
 MUX2_X1 _26229_ (.A(_18692_),
    .B(_19094_),
    .S(_19034_),
    .Z(_03886_));
 OAI221_X1 _26230_ (.A(_18700_),
    .B1(_18672_),
    .B2(_19317_),
    .C1(_03886_),
    .C2(_18770_),
    .ZN(_03887_));
 MUX2_X1 _26231_ (.A(_18647_),
    .B(_18783_),
    .S(_18763_),
    .Z(_03888_));
 AOI22_X1 _26232_ (.A1(_18636_),
    .A2(_18703_),
    .B1(_03888_),
    .B2(_18832_),
    .ZN(_03889_));
 OAI221_X1 _26233_ (.A(_18807_),
    .B1(_18744_),
    .B2(_18782_),
    .C1(_03889_),
    .C2(_18823_),
    .ZN(_03890_));
 AOI21_X1 _26234_ (.A(_03885_),
    .B1(_03887_),
    .B2(_03890_),
    .ZN(_03891_));
 NAND4_X2 _26235_ (.A1(_19090_),
    .A2(_19158_),
    .A3(_03884_),
    .A4(_03891_),
    .ZN(_03892_));
 OAI21_X4 _26236_ (.A(_18416_),
    .B1(_03875_),
    .B2(_03892_),
    .ZN(_03893_));
 AND2_X1 _26237_ (.A1(_00179_),
    .A2(_16982_),
    .ZN(_03894_));
 OAI21_X1 _26238_ (.A(\core.keymem.key_mem[6][118] ),
    .B1(_17146_),
    .B2(_17622_),
    .ZN(_03895_));
 OAI21_X1 _26239_ (.A(\core.keymem.key_mem[10][118] ),
    .B1(_16886_),
    .B2(_16890_),
    .ZN(_03896_));
 AOI21_X2 _26240_ (.A(_16968_),
    .B1(_03895_),
    .B2(_03896_),
    .ZN(_03897_));
 OAI221_X2 _26241_ (.A(\core.keymem.key_mem[5][118] ),
    .B1(_16908_),
    .B2(_16917_),
    .C1(_16913_),
    .C2(_16915_),
    .ZN(_03898_));
 NAND3_X1 _26242_ (.A1(\core.keymem.key_mem[12][118] ),
    .A2(_17099_),
    .A3(_17028_),
    .ZN(_03899_));
 NAND3_X1 _26243_ (.A1(\core.keymem.key_mem[3][118] ),
    .A2(_17074_),
    .A3(_16902_),
    .ZN(_03900_));
 NAND3_X1 _26244_ (.A1(\core.keymem.key_mem[14][118] ),
    .A2(_17099_),
    .A3(_17163_),
    .ZN(_03901_));
 NAND4_X2 _26245_ (.A1(_03898_),
    .A2(_03899_),
    .A3(_03900_),
    .A4(_03901_),
    .ZN(_03902_));
 OAI221_X2 _26246_ (.A(\core.keymem.key_mem[9][118] ),
    .B1(_16885_),
    .B2(_16889_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_03903_));
 NAND3_X1 _26247_ (.A1(\core.keymem.key_mem[2][118] ),
    .A2(_16902_),
    .A3(_17163_),
    .ZN(_03904_));
 OAI211_X2 _26248_ (.A(\core.keymem.key_mem[13][118] ),
    .B(_16919_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_03905_));
 OAI211_X2 _26249_ (.A(\core.keymem.key_mem[8][118] ),
    .B(_16931_),
    .C1(_16927_),
    .C2(_16929_),
    .ZN(_03906_));
 NAND4_X2 _26250_ (.A1(_03903_),
    .A2(_03904_),
    .A3(_03905_),
    .A4(_03906_),
    .ZN(_03907_));
 OAI211_X2 _26251_ (.A(\core.keymem.key_mem[1][118] ),
    .B(_16902_),
    .C1(_16913_),
    .C2(_16915_),
    .ZN(_03908_));
 OAI211_X2 _26252_ (.A(\core.keymem.key_mem[7][118] ),
    .B(_16901_),
    .C1(_16896_),
    .C2(_16899_),
    .ZN(_03909_));
 OAI211_X2 _26253_ (.A(\core.keymem.key_mem[4][118] ),
    .B(_16931_),
    .C1(_16908_),
    .C2(_16917_),
    .ZN(_03910_));
 OAI211_X2 _26254_ (.A(\core.keymem.key_mem[11][118] ),
    .B(_16901_),
    .C1(_16922_),
    .C2(_16923_),
    .ZN(_03911_));
 NAND4_X2 _26255_ (.A1(_03908_),
    .A2(_03909_),
    .A3(_03910_),
    .A4(_03911_),
    .ZN(_03912_));
 NOR4_X4 _26256_ (.A1(_03897_),
    .A2(_03902_),
    .A3(_03907_),
    .A4(_03912_),
    .ZN(_03913_));
 AOI21_X4 _26257_ (.A(_03894_),
    .B1(_03913_),
    .B2(_16488_),
    .ZN(_03914_));
 XNOR2_X2 _26258_ (.A(\core.dec_block.block_w0_reg[22] ),
    .B(_03914_),
    .ZN(_03915_));
 XOR2_X2 _26259_ (.A(\block_reg[3][22] ),
    .B(_18920_),
    .Z(_03916_));
 OAI221_X2 _26260_ (.A(_18329_),
    .B1(_17741_),
    .B2(_03915_),
    .C1(_03916_),
    .C2(_18553_),
    .ZN(_03917_));
 XNOR2_X2 _26261_ (.A(_03326_),
    .B(_03783_),
    .ZN(_03918_));
 XNOR2_X2 _26262_ (.A(_03762_),
    .B(_03776_),
    .ZN(_03919_));
 XOR2_X1 _26263_ (.A(_03918_),
    .B(_03919_),
    .Z(_03920_));
 XNOR2_X2 _26264_ (.A(_03760_),
    .B(_03790_),
    .ZN(_03921_));
 XNOR2_X1 _26265_ (.A(_18884_),
    .B(_18956_),
    .ZN(_03922_));
 XNOR2_X1 _26266_ (.A(_19441_),
    .B(_03922_),
    .ZN(_03923_));
 XNOR2_X1 _26267_ (.A(_03921_),
    .B(_03923_),
    .ZN(_03924_));
 XNOR2_X2 _26268_ (.A(_18909_),
    .B(_19246_),
    .ZN(_03925_));
 XNOR2_X2 _26269_ (.A(_19225_),
    .B(_03925_),
    .ZN(_03926_));
 XNOR2_X1 _26270_ (.A(_03924_),
    .B(_03926_),
    .ZN(_03927_));
 XNOR2_X1 _26271_ (.A(_03920_),
    .B(_03927_),
    .ZN(_03928_));
 AOI21_X1 _26272_ (.A(_03917_),
    .B1(_03928_),
    .B2(_19031_),
    .ZN(_03929_));
 AOI21_X1 _26273_ (.A(_03861_),
    .B1(_03893_),
    .B2(_03929_),
    .ZN(_00581_));
 AOI22_X1 _26274_ (.A1(_18685_),
    .A2(_18793_),
    .B1(_19322_),
    .B2(_19071_),
    .ZN(_03930_));
 NOR3_X1 _26275_ (.A1(_18658_),
    .A2(_18796_),
    .A3(_03930_),
    .ZN(_03931_));
 OAI33_X1 _26276_ (.A1(_18621_),
    .A2(_18741_),
    .A3(_18635_),
    .B1(_18598_),
    .B2(_18697_),
    .B3(_18674_),
    .ZN(_03932_));
 OAI22_X1 _26277_ (.A1(_18782_),
    .A2(_18666_),
    .B1(_18689_),
    .B2(_19168_),
    .ZN(_03933_));
 AOI221_X1 _26278_ (.A(_03931_),
    .B1(_03932_),
    .B2(_18816_),
    .C1(_03933_),
    .C2(_18699_),
    .ZN(_03934_));
 NOR3_X1 _26279_ (.A1(_18780_),
    .A2(_18711_),
    .A3(_19104_),
    .ZN(_03935_));
 OAI221_X1 _26280_ (.A(_03671_),
    .B1(_03935_),
    .B2(_19113_),
    .C1(_19317_),
    .C2(_18801_),
    .ZN(_03936_));
 AOI21_X1 _26281_ (.A(_18785_),
    .B1(_03936_),
    .B2(_18700_),
    .ZN(_03937_));
 NAND2_X1 _26282_ (.A1(_18768_),
    .A2(_19132_),
    .ZN(_03938_));
 AOI21_X1 _26283_ (.A(_18653_),
    .B1(_18810_),
    .B2(_18709_),
    .ZN(_03939_));
 AOI21_X1 _26284_ (.A(_03939_),
    .B1(_18719_),
    .B2(_18779_),
    .ZN(_03940_));
 OAI221_X2 _26285_ (.A(_03938_),
    .B1(_03940_),
    .B2(_18640_),
    .C1(_18770_),
    .C2(_03886_),
    .ZN(_03941_));
 NOR4_X1 _26286_ (.A1(_18734_),
    .A2(_03819_),
    .A3(_03821_),
    .A4(_03941_),
    .ZN(_03942_));
 AND4_X1 _26287_ (.A1(_03666_),
    .A2(_03934_),
    .A3(_03937_),
    .A4(_03942_),
    .ZN(_03943_));
 AND2_X1 _26288_ (.A1(_19314_),
    .A2(_19357_),
    .ZN(_03944_));
 AOI22_X2 _26289_ (.A1(_18682_),
    .A2(_18712_),
    .B1(_18765_),
    .B2(_03944_),
    .ZN(_03945_));
 OAI221_X2 _26290_ (.A(_03945_),
    .B1(_19135_),
    .B2(_18666_),
    .C1(_18782_),
    .C2(_18696_),
    .ZN(_03946_));
 NOR2_X1 _26291_ (.A1(_18808_),
    .A2(_19040_),
    .ZN(_03947_));
 OAI21_X1 _26292_ (.A(_18708_),
    .B1(_18774_),
    .B2(_03947_),
    .ZN(_03948_));
 OAI221_X2 _26293_ (.A(_03948_),
    .B1(_18733_),
    .B2(_19364_),
    .C1(_18747_),
    .C2(_18810_),
    .ZN(_03949_));
 NOR4_X2 _26294_ (.A1(_19312_),
    .A2(_19512_),
    .A3(_03946_),
    .A4(_03949_),
    .ZN(_03950_));
 OAI21_X1 _26295_ (.A(_18693_),
    .B1(_18719_),
    .B2(_19094_),
    .ZN(_03951_));
 NAND2_X1 _26296_ (.A1(_18806_),
    .A2(_19104_),
    .ZN(_03952_));
 AOI21_X1 _26297_ (.A(_18719_),
    .B1(_19484_),
    .B2(_03952_),
    .ZN(_03953_));
 AOI221_X2 _26298_ (.A(_19041_),
    .B1(_03951_),
    .B2(_18703_),
    .C1(_03953_),
    .C2(_18659_),
    .ZN(_03954_));
 NAND4_X4 _26299_ (.A1(_03884_),
    .A2(_03943_),
    .A3(_03950_),
    .A4(_03954_),
    .ZN(_03955_));
 INV_X1 _26300_ (.A(\block_reg[3][23] ),
    .ZN(_03956_));
 XNOR2_X2 _26301_ (.A(_03956_),
    .B(_18955_),
    .ZN(_03957_));
 AOI21_X1 _26302_ (.A(_16367_),
    .B1(_16371_),
    .B2(_03957_),
    .ZN(_03958_));
 XNOR2_X2 _26303_ (.A(_03775_),
    .B(_03921_),
    .ZN(_03959_));
 XNOR2_X1 _26304_ (.A(_19262_),
    .B(_03959_),
    .ZN(_03960_));
 XNOR2_X2 _26305_ (.A(_19441_),
    .B(_03739_),
    .ZN(_03961_));
 XNOR2_X2 _26306_ (.A(_19224_),
    .B(_03961_),
    .ZN(_03962_));
 XNOR2_X2 _26307_ (.A(_18922_),
    .B(_03962_),
    .ZN(_03963_));
 XNOR2_X2 _26308_ (.A(_03960_),
    .B(_03963_),
    .ZN(_03964_));
 NAND2_X1 _26309_ (.A1(_00190_),
    .A2(_16871_),
    .ZN(_03965_));
 AOI222_X2 _26310_ (.A1(\core.keymem.key_mem[10][119] ),
    .A2(_16514_),
    .B1(_16441_),
    .B2(\core.keymem.key_mem[11][119] ),
    .C1(\core.keymem.key_mem[13][119] ),
    .C2(_16471_),
    .ZN(_03966_));
 AOI22_X2 _26311_ (.A1(\core.keymem.key_mem[4][119] ),
    .A2(_16499_),
    .B1(_16524_),
    .B2(\core.keymem.key_mem[1][119] ),
    .ZN(_03967_));
 AOI22_X2 _26312_ (.A1(\core.keymem.key_mem[7][119] ),
    .A2(_17736_),
    .B1(_16528_),
    .B2(\core.keymem.key_mem[8][119] ),
    .ZN(_03968_));
 NAND3_X2 _26313_ (.A1(_03966_),
    .A2(_03967_),
    .A3(_03968_),
    .ZN(_03969_));
 AOI21_X1 _26314_ (.A(_16494_),
    .B1(_16993_),
    .B2(\core.keymem.key_mem[2][119] ),
    .ZN(_03970_));
 AOI22_X2 _26315_ (.A1(\core.keymem.key_mem[14][119] ),
    .A2(_17191_),
    .B1(_16865_),
    .B2(\core.keymem.key_mem[3][119] ),
    .ZN(_03971_));
 AOI22_X2 _26316_ (.A1(\core.keymem.key_mem[9][119] ),
    .A2(_16535_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][119] ),
    .ZN(_03972_));
 AOI22_X2 _26317_ (.A1(\core.keymem.key_mem[6][119] ),
    .A2(_17648_),
    .B1(_16467_),
    .B2(\core.keymem.key_mem[5][119] ),
    .ZN(_03973_));
 NAND4_X2 _26318_ (.A1(_03970_),
    .A2(_03971_),
    .A3(_03972_),
    .A4(_03973_),
    .ZN(_03974_));
 OAI21_X4 _26319_ (.A(_03965_),
    .B1(_03969_),
    .B2(_03974_),
    .ZN(_03975_));
 XOR2_X2 _26320_ (.A(_18574_),
    .B(_03975_),
    .Z(_03976_));
 OAI221_X1 _26321_ (.A(_03958_),
    .B1(_03964_),
    .B2(_17203_),
    .C1(_16556_),
    .C2(_03976_),
    .ZN(_03977_));
 OAI22_X1 _26322_ (.A1(_18574_),
    .A2(_16366_),
    .B1(_03955_),
    .B2(_03977_),
    .ZN(_03978_));
 INV_X1 _26323_ (.A(_03978_),
    .ZN(_00582_));
 NOR2_X1 _26324_ (.A1(\core.dec_block.block_w0_reg[24] ),
    .A2(_18330_),
    .ZN(_03979_));
 NAND2_X1 _26325_ (.A1(_16357_),
    .A2(\core.dec_block.block_w0_reg[26] ),
    .ZN(_03980_));
 AOI222_X2 _26326_ (.A1(\core.dec_block.block_w2_reg[26] ),
    .A2(_16566_),
    .B1(_16266_),
    .B2(\core.dec_block.block_w3_reg[26] ),
    .C1(_16568_),
    .C2(\core.dec_block.block_w1_reg[26] ),
    .ZN(_03981_));
 OAI21_X4 _26327_ (.A(_03980_),
    .B1(_03981_),
    .B2(_16584_),
    .ZN(_03982_));
 NAND2_X4 _26328_ (.A1(_16560_),
    .A2(_03982_),
    .ZN(_03983_));
 NAND2_X1 _26329_ (.A1(_16357_),
    .A2(\core.dec_block.block_w0_reg[27] ),
    .ZN(_03984_));
 AOI222_X2 _26330_ (.A1(\core.dec_block.block_w2_reg[27] ),
    .A2(_16565_),
    .B1(_16266_),
    .B2(\core.dec_block.block_w3_reg[27] ),
    .C1(_16568_),
    .C2(\core.dec_block.block_w1_reg[27] ),
    .ZN(_03985_));
 OAI21_X4 _26331_ (.A(_03984_),
    .B1(_03985_),
    .B2(_16357_),
    .ZN(_03986_));
 AND2_X2 _26332_ (.A1(_16562_),
    .A2(_03986_),
    .ZN(_03987_));
 NOR2_X2 _26333_ (.A1(_03983_),
    .A2(_03987_),
    .ZN(_03988_));
 BUF_X4 _26334_ (.A(_03988_),
    .Z(_03989_));
 NAND2_X1 _26335_ (.A1(_18566_),
    .A2(\core.dec_block.block_w0_reg[25] ),
    .ZN(_03990_));
 AOI222_X2 _26336_ (.A1(\core.dec_block.block_w2_reg[25] ),
    .A2(_18569_),
    .B1(_16268_),
    .B2(\core.dec_block.block_w3_reg[25] ),
    .C1(_18568_),
    .C2(\core.dec_block.block_w1_reg[25] ),
    .ZN(_03991_));
 OAI21_X4 _26337_ (.A(_03990_),
    .B1(_03991_),
    .B2(_16359_),
    .ZN(_03992_));
 AND2_X2 _26338_ (.A1(_16622_),
    .A2(_03992_),
    .ZN(_03993_));
 BUF_X4 _26339_ (.A(_03993_),
    .Z(_03994_));
 BUF_X4 _26340_ (.A(_03994_),
    .Z(_03995_));
 CLKBUF_X3 _26341_ (.A(_03995_),
    .Z(_03996_));
 NAND2_X1 _26342_ (.A1(\core.dec_block.block_w0_reg[24] ),
    .A2(_16358_),
    .ZN(_03997_));
 AOI222_X2 _26343_ (.A1(\core.dec_block.block_w2_reg[24] ),
    .A2(_16566_),
    .B1(_16267_),
    .B2(\core.dec_block.block_w3_reg[24] ),
    .C1(_16569_),
    .C2(\core.dec_block.block_w1_reg[24] ),
    .ZN(_03998_));
 OAI21_X4 _26344_ (.A(_03997_),
    .B1(_03998_),
    .B2(_18566_),
    .ZN(_03999_));
 NAND2_X4 _26345_ (.A1(_16622_),
    .A2(_03999_),
    .ZN(_04000_));
 BUF_X4 _26346_ (.A(_04000_),
    .Z(_04001_));
 BUF_X4 _26347_ (.A(_04001_),
    .Z(_04002_));
 BUF_X2 _26348_ (.A(\core.dec_block.block_w0_reg[31] ),
    .Z(_04003_));
 NAND2_X1 _26349_ (.A1(_04003_),
    .A2(_16584_),
    .ZN(_04004_));
 AOI222_X2 _26350_ (.A1(\core.dec_block.block_w2_reg[31] ),
    .A2(_16566_),
    .B1(_16267_),
    .B2(\core.dec_block.block_w3_reg[31] ),
    .C1(_16569_),
    .C2(\core.dec_block.block_w1_reg[31] ),
    .ZN(_04005_));
 OAI21_X2 _26351_ (.A(_04004_),
    .B1(_04005_),
    .B2(_16358_),
    .ZN(_04006_));
 AND2_X1 _26352_ (.A1(_16561_),
    .A2(_04006_),
    .ZN(_04007_));
 BUF_X4 _26353_ (.A(_04007_),
    .Z(_04008_));
 NAND2_X1 _26354_ (.A1(_16584_),
    .A2(\core.dec_block.block_w0_reg[30] ),
    .ZN(_04009_));
 AOI222_X2 _26355_ (.A1(\core.dec_block.block_w2_reg[30] ),
    .A2(_16566_),
    .B1(_16267_),
    .B2(\core.dec_block.block_w3_reg[30] ),
    .C1(_16569_),
    .C2(\core.dec_block.block_w1_reg[30] ),
    .ZN(_04010_));
 OAI21_X2 _26356_ (.A(_04009_),
    .B1(_04010_),
    .B2(_16584_),
    .ZN(_04011_));
 AND2_X1 _26357_ (.A1(_16561_),
    .A2(_04011_),
    .ZN(_04012_));
 BUF_X4 _26358_ (.A(_04012_),
    .Z(_04013_));
 NAND2_X4 _26359_ (.A1(_04008_),
    .A2(_04013_),
    .ZN(_04014_));
 NAND2_X1 _26360_ (.A1(\core.dec_block.block_w0_reg[29] ),
    .A2(_16357_),
    .ZN(_04015_));
 AOI222_X2 _26361_ (.A1(\core.dec_block.block_w2_reg[29] ),
    .A2(_16565_),
    .B1(_16266_),
    .B2(\core.dec_block.block_w3_reg[29] ),
    .C1(_16568_),
    .C2(\core.dec_block.block_w1_reg[29] ),
    .ZN(_04016_));
 OAI21_X2 _26362_ (.A(_04015_),
    .B1(_04016_),
    .B2(_16584_),
    .ZN(_04017_));
 AND2_X1 _26363_ (.A1(_16561_),
    .A2(_04017_),
    .ZN(_04018_));
 BUF_X4 _26364_ (.A(_04018_),
    .Z(_04019_));
 NAND2_X1 _26365_ (.A1(_16356_),
    .A2(\core.dec_block.block_w0_reg[28] ),
    .ZN(_04020_));
 AOI222_X2 _26366_ (.A1(\core.dec_block.block_w2_reg[28] ),
    .A2(_16565_),
    .B1(_16265_),
    .B2(\core.dec_block.block_w3_reg[28] ),
    .C1(_16568_),
    .C2(\core.dec_block.block_w1_reg[28] ),
    .ZN(_04021_));
 OAI21_X2 _26367_ (.A(_04020_),
    .B1(_04021_),
    .B2(_16356_),
    .ZN(_04022_));
 NAND2_X4 _26368_ (.A1(_16562_),
    .A2(_04022_),
    .ZN(_04023_));
 NAND2_X4 _26369_ (.A1(_04019_),
    .A2(_04023_),
    .ZN(_04024_));
 NOR2_X4 _26370_ (.A1(_04014_),
    .A2(_04024_),
    .ZN(_04025_));
 NAND3_X1 _26371_ (.A1(_03996_),
    .A2(_04002_),
    .A3(_04025_),
    .ZN(_04026_));
 AND2_X1 _26372_ (.A1(_16562_),
    .A2(_03999_),
    .ZN(_04027_));
 BUF_X4 _26373_ (.A(_04027_),
    .Z(_04028_));
 BUF_X4 _26374_ (.A(_04028_),
    .Z(_04029_));
 BUF_X4 _26375_ (.A(_04029_),
    .Z(_04030_));
 AND2_X1 _26376_ (.A1(_16559_),
    .A2(_04022_),
    .ZN(_04031_));
 BUF_X4 _26377_ (.A(_04031_),
    .Z(_04032_));
 NAND2_X4 _26378_ (.A1(_04019_),
    .A2(_04032_),
    .ZN(_04033_));
 NOR2_X4 _26379_ (.A1(_04014_),
    .A2(_04033_),
    .ZN(_04034_));
 NAND2_X1 _26380_ (.A1(_04030_),
    .A2(_04034_),
    .ZN(_04035_));
 OAI21_X1 _26381_ (.A(_04026_),
    .B1(_04035_),
    .B2(_03996_),
    .ZN(_04036_));
 NAND2_X1 _26382_ (.A1(_03989_),
    .A2(_04036_),
    .ZN(_04037_));
 AND2_X1 _26383_ (.A1(_16576_),
    .A2(_03982_),
    .ZN(_04038_));
 BUF_X4 _26384_ (.A(_04038_),
    .Z(_04039_));
 NAND2_X2 _26385_ (.A1(_16560_),
    .A2(_03986_),
    .ZN(_04040_));
 BUF_X4 _26386_ (.A(_04040_),
    .Z(_04041_));
 NAND2_X4 _26387_ (.A1(_04039_),
    .A2(_04041_),
    .ZN(_04042_));
 BUF_X4 _26388_ (.A(_04042_),
    .Z(_04043_));
 NAND2_X4 _26389_ (.A1(_16622_),
    .A2(_03992_),
    .ZN(_04044_));
 BUF_X4 _26390_ (.A(_04044_),
    .Z(_04045_));
 BUF_X4 _26391_ (.A(_04045_),
    .Z(_04046_));
 BUF_X4 _26392_ (.A(_04046_),
    .Z(_04047_));
 BUF_X4 _26393_ (.A(_04030_),
    .Z(_04048_));
 NAND2_X2 _26394_ (.A1(_16560_),
    .A2(_04017_),
    .ZN(_04049_));
 BUF_X4 _26395_ (.A(_04049_),
    .Z(_04050_));
 NOR2_X4 _26396_ (.A1(_04050_),
    .A2(_04023_),
    .ZN(_04051_));
 NAND2_X2 _26397_ (.A1(_16561_),
    .A2(_04011_),
    .ZN(_04052_));
 BUF_X4 _26398_ (.A(_04052_),
    .Z(_04053_));
 NOR2_X4 _26399_ (.A1(_04008_),
    .A2(_04053_),
    .ZN(_04054_));
 NAND2_X4 _26400_ (.A1(_04051_),
    .A2(_04054_),
    .ZN(_04055_));
 NOR4_X2 _26401_ (.A1(_04043_),
    .A2(_04047_),
    .A3(_04048_),
    .A4(_04055_),
    .ZN(_04056_));
 BUF_X4 _26402_ (.A(_03983_),
    .Z(_04057_));
 BUF_X4 _26403_ (.A(_04057_),
    .Z(_04058_));
 BUF_X4 _26404_ (.A(_04041_),
    .Z(_04059_));
 NAND2_X2 _26405_ (.A1(_04059_),
    .A2(_04030_),
    .ZN(_04060_));
 BUF_X4 _26406_ (.A(_04055_),
    .Z(_04061_));
 NOR2_X4 _26407_ (.A1(_04019_),
    .A2(_04032_),
    .ZN(_04062_));
 NAND2_X4 _26408_ (.A1(_16562_),
    .A2(_04006_),
    .ZN(_04063_));
 NOR2_X4 _26409_ (.A1(_04063_),
    .A2(_04013_),
    .ZN(_04064_));
 NAND2_X4 _26410_ (.A1(_04062_),
    .A2(_04064_),
    .ZN(_04065_));
 NAND2_X1 _26411_ (.A1(_04058_),
    .A2(_04001_),
    .ZN(_04066_));
 OAI33_X1 _26412_ (.A1(_04058_),
    .A2(_04060_),
    .A3(_04061_),
    .B1(_04065_),
    .B2(_04066_),
    .B3(_04059_),
    .ZN(_04067_));
 BUF_X4 _26413_ (.A(_04046_),
    .Z(_04068_));
 BUF_X4 _26414_ (.A(_03987_),
    .Z(_04069_));
 BUF_X4 _26415_ (.A(_04069_),
    .Z(_04070_));
 BUF_X4 _26416_ (.A(_04070_),
    .Z(_04071_));
 CLKBUF_X3 _26417_ (.A(_04071_),
    .Z(_04072_));
 BUF_X4 _26418_ (.A(_04039_),
    .Z(_04073_));
 BUF_X4 _26419_ (.A(_04073_),
    .Z(_04074_));
 NOR2_X4 _26420_ (.A1(_04063_),
    .A2(_04052_),
    .ZN(_04075_));
 NOR2_X4 _26421_ (.A1(_04019_),
    .A2(_04023_),
    .ZN(_04076_));
 NAND2_X4 _26422_ (.A1(_04075_),
    .A2(_04076_),
    .ZN(_04077_));
 NOR2_X2 _26423_ (.A1(_04074_),
    .A2(_04077_),
    .ZN(_04078_));
 NAND2_X1 _26424_ (.A1(_04048_),
    .A2(_04078_),
    .ZN(_04079_));
 NAND2_X4 _26425_ (.A1(_04050_),
    .A2(_04023_),
    .ZN(_04080_));
 NAND2_X4 _26426_ (.A1(_04063_),
    .A2(_04013_),
    .ZN(_04081_));
 NOR2_X1 _26427_ (.A1(_04080_),
    .A2(_04081_),
    .ZN(_04082_));
 CLKBUF_X3 _26428_ (.A(_04082_),
    .Z(_04083_));
 BUF_X4 _26429_ (.A(_04073_),
    .Z(_04084_));
 AOI21_X1 _26430_ (.A(_04078_),
    .B1(_04083_),
    .B2(_04084_),
    .ZN(_04085_));
 BUF_X4 _26431_ (.A(_03995_),
    .Z(_04086_));
 OAI21_X1 _26432_ (.A(_04079_),
    .B1(_04085_),
    .B2(_04086_),
    .ZN(_04087_));
 AOI221_X2 _26433_ (.A(_04056_),
    .B1(_04067_),
    .B2(_04068_),
    .C1(_04072_),
    .C2(_04087_),
    .ZN(_04088_));
 NAND2_X1 _26434_ (.A1(_04037_),
    .A2(_04088_),
    .ZN(_04089_));
 NOR2_X4 _26435_ (.A1(_04039_),
    .A2(_03987_),
    .ZN(_04090_));
 BUF_X4 _26436_ (.A(_04090_),
    .Z(_04091_));
 NAND2_X1 _26437_ (.A1(_03996_),
    .A2(_04025_),
    .ZN(_04092_));
 NAND2_X4 _26438_ (.A1(_04063_),
    .A2(_04053_),
    .ZN(_04093_));
 NOR2_X4 _26439_ (.A1(_04080_),
    .A2(_04093_),
    .ZN(_04094_));
 NAND2_X1 _26440_ (.A1(_04030_),
    .A2(_04094_),
    .ZN(_04095_));
 OAI21_X1 _26441_ (.A(_04092_),
    .B1(_04095_),
    .B2(_03996_),
    .ZN(_04096_));
 NAND2_X1 _26442_ (.A1(_04091_),
    .A2(_04096_),
    .ZN(_04097_));
 NOR2_X4 _26443_ (.A1(_04050_),
    .A2(_04032_),
    .ZN(_04098_));
 NAND2_X1 _26444_ (.A1(_04098_),
    .A2(_04064_),
    .ZN(_04099_));
 NOR2_X1 _26445_ (.A1(_04069_),
    .A2(_04099_),
    .ZN(_04100_));
 NOR2_X4 _26446_ (.A1(_04041_),
    .A2(_03994_),
    .ZN(_04101_));
 AOI21_X1 _26447_ (.A(_04100_),
    .B1(_04101_),
    .B2(_04034_),
    .ZN(_04102_));
 NOR2_X2 _26448_ (.A1(_04058_),
    .A2(_04102_),
    .ZN(_04103_));
 NAND2_X2 _26449_ (.A1(_04076_),
    .A2(_04064_),
    .ZN(_04104_));
 NOR2_X4 _26450_ (.A1(_04008_),
    .A2(_04013_),
    .ZN(_04105_));
 NAND2_X1 _26451_ (.A1(_04098_),
    .A2(_04105_),
    .ZN(_04106_));
 BUF_X4 _26452_ (.A(_04106_),
    .Z(_04107_));
 OAI21_X1 _26453_ (.A(_04104_),
    .B1(_04107_),
    .B2(_04045_),
    .ZN(_04108_));
 NOR2_X2 _26454_ (.A1(_04024_),
    .A2(_04081_),
    .ZN(_04109_));
 BUF_X4 _26455_ (.A(_04109_),
    .Z(_04110_));
 NAND2_X4 _26456_ (.A1(_04057_),
    .A2(_04069_),
    .ZN(_04111_));
 NAND2_X2 _26457_ (.A1(_03993_),
    .A2(_04028_),
    .ZN(_04112_));
 NOR2_X2 _26458_ (.A1(_04111_),
    .A2(_04112_),
    .ZN(_04113_));
 AOI221_X2 _26459_ (.A(_04103_),
    .B1(_04108_),
    .B2(_03989_),
    .C1(_04110_),
    .C2(_04113_),
    .ZN(_04114_));
 CLKBUF_X3 _26460_ (.A(_04059_),
    .Z(_04115_));
 NOR4_X1 _26461_ (.A1(_04057_),
    .A2(_04063_),
    .A3(_04053_),
    .A4(_04032_),
    .ZN(_04116_));
 CLKBUF_X3 _26462_ (.A(_04023_),
    .Z(_04117_));
 NAND4_X1 _26463_ (.A1(_04057_),
    .A2(_03994_),
    .A3(_04053_),
    .A4(_04117_),
    .ZN(_04118_));
 XNOR2_X1 _26464_ (.A(_04073_),
    .B(_04013_),
    .ZN(_04119_));
 OAI21_X1 _26465_ (.A(_04118_),
    .B1(_04119_),
    .B2(_04117_),
    .ZN(_04120_));
 BUF_X2 _26466_ (.A(_04063_),
    .Z(_04121_));
 AOI21_X1 _26467_ (.A(_04116_),
    .B1(_04120_),
    .B2(_04121_),
    .ZN(_04122_));
 OR3_X1 _26468_ (.A1(_04115_),
    .A2(_04050_),
    .A3(_04122_),
    .ZN(_04123_));
 NAND3_X2 _26469_ (.A1(_04097_),
    .A2(_04114_),
    .A3(_04123_),
    .ZN(_04124_));
 NAND2_X4 _26470_ (.A1(_04044_),
    .A2(_04028_),
    .ZN(_04125_));
 NAND2_X2 _26471_ (.A1(_04051_),
    .A2(_04105_),
    .ZN(_04126_));
 BUF_X4 _26472_ (.A(_04126_),
    .Z(_04127_));
 NAND2_X2 _26473_ (.A1(_03993_),
    .A2(_04000_),
    .ZN(_04128_));
 BUF_X4 _26474_ (.A(_04128_),
    .Z(_04129_));
 NAND2_X4 _26475_ (.A1(_04051_),
    .A2(_04064_),
    .ZN(_04130_));
 OAI22_X2 _26476_ (.A1(_04125_),
    .A2(_04127_),
    .B1(_04129_),
    .B2(_04130_),
    .ZN(_04131_));
 BUF_X4 _26477_ (.A(_03996_),
    .Z(_04132_));
 NOR2_X2 _26478_ (.A1(_04001_),
    .A2(_04130_),
    .ZN(_04133_));
 AOI21_X1 _26479_ (.A(_04100_),
    .B1(_04133_),
    .B2(_04071_),
    .ZN(_04134_));
 NAND2_X4 _26480_ (.A1(_04008_),
    .A2(_04053_),
    .ZN(_04135_));
 NOR2_X1 _26481_ (.A1(_04024_),
    .A2(_04135_),
    .ZN(_04136_));
 CLKBUF_X3 _26482_ (.A(_04136_),
    .Z(_04137_));
 NOR2_X1 _26483_ (.A1(_04033_),
    .A2(_04135_),
    .ZN(_04138_));
 CLKBUF_X3 _26484_ (.A(_04138_),
    .Z(_04139_));
 AOI21_X1 _26485_ (.A(_04137_),
    .B1(_04139_),
    .B2(_04086_),
    .ZN(_04140_));
 OAI22_X2 _26486_ (.A1(_04132_),
    .A2(_04134_),
    .B1(_04140_),
    .B2(_04060_),
    .ZN(_04141_));
 BUF_X4 _26487_ (.A(_04058_),
    .Z(_04142_));
 BUF_X4 _26488_ (.A(_04142_),
    .Z(_04143_));
 AOI22_X2 _26489_ (.A1(_03989_),
    .A2(_04131_),
    .B1(_04141_),
    .B2(_04143_),
    .ZN(_04144_));
 NAND2_X1 _26490_ (.A1(_04075_),
    .A2(_04062_),
    .ZN(_04145_));
 NAND2_X2 _26491_ (.A1(_04125_),
    .A2(_04128_),
    .ZN(_04146_));
 NOR3_X1 _26492_ (.A1(_04057_),
    .A2(_04145_),
    .A3(_04146_),
    .ZN(_04147_));
 NAND2_X4 _26493_ (.A1(_04075_),
    .A2(_04098_),
    .ZN(_04148_));
 NOR2_X1 _26494_ (.A1(_03993_),
    .A2(_04000_),
    .ZN(_04149_));
 NOR2_X4 _26495_ (.A1(_04044_),
    .A2(_04028_),
    .ZN(_04150_));
 NOR2_X2 _26496_ (.A1(_04149_),
    .A2(_04150_),
    .ZN(_04151_));
 NOR3_X1 _26497_ (.A1(_04074_),
    .A2(_04148_),
    .A3(_04151_),
    .ZN(_04152_));
 OAI21_X1 _26498_ (.A(_04070_),
    .B1(_04147_),
    .B2(_04152_),
    .ZN(_04153_));
 NAND2_X4 _26499_ (.A1(_04049_),
    .A2(_04032_),
    .ZN(_04154_));
 NOR2_X1 _26500_ (.A1(_04154_),
    .A2(_04093_),
    .ZN(_04155_));
 CLKBUF_X3 _26501_ (.A(_04155_),
    .Z(_04156_));
 NOR2_X4 _26502_ (.A1(_04014_),
    .A2(_04080_),
    .ZN(_04157_));
 AOI21_X1 _26503_ (.A(_04156_),
    .B1(_04157_),
    .B2(_04146_),
    .ZN(_04158_));
 OAI21_X1 _26504_ (.A(_04153_),
    .B1(_04158_),
    .B2(_04043_),
    .ZN(_04159_));
 NAND2_X4 _26505_ (.A1(_03983_),
    .A2(_04041_),
    .ZN(_04160_));
 NOR2_X2 _26506_ (.A1(_04160_),
    .A2(_04128_),
    .ZN(_04161_));
 NOR2_X4 _26507_ (.A1(_03993_),
    .A2(_04160_),
    .ZN(_04162_));
 AOI221_X2 _26508_ (.A(_04159_),
    .B1(_04161_),
    .B2(_04110_),
    .C1(_04034_),
    .C2(_04162_),
    .ZN(_04163_));
 NAND2_X4 _26509_ (.A1(_04041_),
    .A2(_03994_),
    .ZN(_04164_));
 NAND2_X2 _26510_ (.A1(_04030_),
    .A2(_04157_),
    .ZN(_04165_));
 NOR2_X4 _26511_ (.A1(_04154_),
    .A2(_04081_),
    .ZN(_04166_));
 NAND2_X1 _26512_ (.A1(_04074_),
    .A2(_04166_),
    .ZN(_04167_));
 NOR2_X1 _26513_ (.A1(_04069_),
    .A2(_04029_),
    .ZN(_04168_));
 NAND2_X4 _26514_ (.A1(_04069_),
    .A2(_04028_),
    .ZN(_04169_));
 AOI21_X1 _26515_ (.A(_04168_),
    .B1(_04169_),
    .B2(_04046_),
    .ZN(_04170_));
 OAI22_X2 _26516_ (.A1(_04164_),
    .A2(_04165_),
    .B1(_04167_),
    .B2(_04170_),
    .ZN(_04171_));
 NOR2_X1 _26517_ (.A1(_04045_),
    .A2(_04160_),
    .ZN(_04172_));
 NAND2_X2 _26518_ (.A1(_04076_),
    .A2(_04105_),
    .ZN(_04173_));
 BUF_X4 _26519_ (.A(_04173_),
    .Z(_04174_));
 OAI21_X1 _26520_ (.A(_04077_),
    .B1(_04174_),
    .B2(_04030_),
    .ZN(_04175_));
 NAND2_X4 _26521_ (.A1(_04062_),
    .A2(_04105_),
    .ZN(_04176_));
 NOR2_X1 _26522_ (.A1(_04034_),
    .A2(_04137_),
    .ZN(_04177_));
 OAI221_X2 _26523_ (.A(_04035_),
    .B1(_04176_),
    .B2(_04030_),
    .C1(_04177_),
    .C2(_03996_),
    .ZN(_04178_));
 NOR2_X4 _26524_ (.A1(_04039_),
    .A2(_04041_),
    .ZN(_04179_));
 AOI221_X2 _26525_ (.A(_04171_),
    .B1(_04172_),
    .B2(_04175_),
    .C1(_04178_),
    .C2(_04179_),
    .ZN(_04180_));
 CLKBUF_X3 _26526_ (.A(_04048_),
    .Z(_04181_));
 BUF_X4 _26527_ (.A(_04111_),
    .Z(_04182_));
 NOR2_X1 _26528_ (.A1(_04046_),
    .A2(_04174_),
    .ZN(_04183_));
 AOI21_X1 _26529_ (.A(_04183_),
    .B1(_04157_),
    .B2(_04068_),
    .ZN(_04184_));
 NOR3_X1 _26530_ (.A1(_04181_),
    .A2(_04182_),
    .A3(_04184_),
    .ZN(_04185_));
 NOR2_X4 _26531_ (.A1(_04024_),
    .A2(_04093_),
    .ZN(_04186_));
 NAND2_X2 _26532_ (.A1(_04039_),
    .A2(_04186_),
    .ZN(_04187_));
 CLKBUF_X3 _26533_ (.A(_04149_),
    .Z(_04188_));
 NAND2_X1 _26534_ (.A1(_04041_),
    .A2(_04188_),
    .ZN(_04189_));
 OAI33_X1 _26535_ (.A1(_04041_),
    .A2(_04129_),
    .A3(_04187_),
    .B1(_04189_),
    .B2(_04065_),
    .B3(_04073_),
    .ZN(_04190_));
 BUF_X4 _26536_ (.A(_03995_),
    .Z(_04191_));
 BUF_X4 _26537_ (.A(_04077_),
    .Z(_04192_));
 BUF_X4 _26538_ (.A(_04104_),
    .Z(_04193_));
 OAI33_X1 _26539_ (.A1(_04043_),
    .A2(_04191_),
    .A3(_04192_),
    .B1(_04193_),
    .B2(_04151_),
    .B3(_04115_),
    .ZN(_04194_));
 NOR3_X2 _26540_ (.A1(_04185_),
    .A2(_04190_),
    .A3(_04194_),
    .ZN(_04195_));
 NAND4_X2 _26541_ (.A1(_04144_),
    .A2(_04163_),
    .A3(_04180_),
    .A4(_04195_),
    .ZN(_04196_));
 BUF_X4 _26542_ (.A(_04068_),
    .Z(_04197_));
 BUF_X4 _26543_ (.A(_04059_),
    .Z(_04198_));
 NOR3_X1 _26544_ (.A1(_04143_),
    .A2(_04198_),
    .A3(_04192_),
    .ZN(_04199_));
 NOR2_X2 _26545_ (.A1(_04080_),
    .A2(_04135_),
    .ZN(_04200_));
 NAND2_X1 _26546_ (.A1(_04073_),
    .A2(_04200_),
    .ZN(_04201_));
 AOI21_X2 _26547_ (.A(_04002_),
    .B1(_04077_),
    .B2(_04174_),
    .ZN(_04202_));
 OAI21_X1 _26548_ (.A(_04142_),
    .B1(_04157_),
    .B2(_04202_),
    .ZN(_04203_));
 AOI21_X1 _26549_ (.A(_04072_),
    .B1(_04201_),
    .B2(_04203_),
    .ZN(_04204_));
 OAI21_X1 _26550_ (.A(_04197_),
    .B1(_04199_),
    .B2(_04204_),
    .ZN(_04205_));
 NOR2_X4 _26551_ (.A1(_03983_),
    .A2(_04040_),
    .ZN(_04206_));
 BUF_X4 _26552_ (.A(_04206_),
    .Z(_04207_));
 NOR2_X1 _26553_ (.A1(_04008_),
    .A2(_04019_),
    .ZN(_04208_));
 NOR2_X1 _26554_ (.A1(_04150_),
    .A2(_04208_),
    .ZN(_04209_));
 OAI21_X1 _26555_ (.A(_04209_),
    .B1(_04121_),
    .B2(_04086_),
    .ZN(_04210_));
 NOR3_X1 _26556_ (.A1(_04053_),
    .A2(_04117_),
    .A3(_04210_),
    .ZN(_04211_));
 CLKBUF_X3 _26557_ (.A(_04013_),
    .Z(_04212_));
 NOR2_X1 _26558_ (.A1(_04002_),
    .A2(_04121_),
    .ZN(_04213_));
 AOI21_X1 _26559_ (.A(_04208_),
    .B1(_04213_),
    .B2(_04086_),
    .ZN(_04214_));
 NOR3_X1 _26560_ (.A1(_04212_),
    .A2(_04032_),
    .A3(_04214_),
    .ZN(_04215_));
 OAI21_X1 _26561_ (.A(_04207_),
    .B1(_04211_),
    .B2(_04215_),
    .ZN(_04216_));
 NOR3_X1 _26562_ (.A1(_04084_),
    .A2(_04001_),
    .A3(_04126_),
    .ZN(_04217_));
 AOI21_X1 _26563_ (.A(_04217_),
    .B1(_04183_),
    .B2(_04084_),
    .ZN(_04218_));
 NOR2_X2 _26564_ (.A1(_04042_),
    .A2(_04112_),
    .ZN(_04219_));
 INV_X1 _26565_ (.A(_04219_),
    .ZN(_04220_));
 NOR2_X2 _26566_ (.A1(_04044_),
    .A2(_04000_),
    .ZN(_04221_));
 NAND2_X2 _26567_ (.A1(_04179_),
    .A2(_04221_),
    .ZN(_04222_));
 BUF_X4 _26568_ (.A(_04145_),
    .Z(_04223_));
 OAI222_X2 _26569_ (.A1(_04198_),
    .A2(_04218_),
    .B1(_04220_),
    .B2(_04192_),
    .C1(_04222_),
    .C2(_04223_),
    .ZN(_04224_));
 NOR2_X1 _26570_ (.A1(_04000_),
    .A2(_04160_),
    .ZN(_04225_));
 NAND2_X1 _26571_ (.A1(_04186_),
    .A2(_04225_),
    .ZN(_04226_));
 NAND3_X1 _26572_ (.A1(_04048_),
    .A2(_04166_),
    .A3(_04207_),
    .ZN(_04227_));
 AOI21_X1 _26573_ (.A(_04191_),
    .B1(_04226_),
    .B2(_04227_),
    .ZN(_04228_));
 BUF_X4 _26574_ (.A(_04001_),
    .Z(_04229_));
 NAND4_X1 _26575_ (.A1(_04191_),
    .A2(_04229_),
    .A3(_04166_),
    .A4(_04207_),
    .ZN(_04230_));
 INV_X1 _26576_ (.A(_04230_),
    .ZN(_04231_));
 NOR3_X2 _26577_ (.A1(_04224_),
    .A2(_04228_),
    .A3(_04231_),
    .ZN(_04232_));
 XNOR2_X2 _26578_ (.A(_04039_),
    .B(_04029_),
    .ZN(_04233_));
 NOR3_X4 _26579_ (.A1(_04176_),
    .A2(_04164_),
    .A3(_04233_),
    .ZN(_04234_));
 OAI33_X1 _26580_ (.A1(_04160_),
    .A2(_04126_),
    .A3(_04128_),
    .B1(_04164_),
    .B2(_04073_),
    .B3(_04065_),
    .ZN(_04235_));
 NOR2_X1 _26581_ (.A1(_04234_),
    .A2(_04235_),
    .ZN(_04236_));
 NAND2_X4 _26582_ (.A1(_04076_),
    .A2(_04054_),
    .ZN(_04237_));
 NOR2_X1 _26583_ (.A1(_04074_),
    .A2(_04237_),
    .ZN(_04238_));
 NOR2_X1 _26584_ (.A1(_03995_),
    .A2(_04130_),
    .ZN(_04239_));
 AOI21_X1 _26585_ (.A(_04238_),
    .B1(_04239_),
    .B2(_04074_),
    .ZN(_04240_));
 OAI21_X1 _26586_ (.A(_04236_),
    .B1(_04240_),
    .B2(_04169_),
    .ZN(_04241_));
 NAND2_X1 _26587_ (.A1(_04069_),
    .A2(_04233_),
    .ZN(_04242_));
 OAI22_X2 _26588_ (.A1(_04058_),
    .A2(_04129_),
    .B1(_04242_),
    .B2(_03995_),
    .ZN(_04243_));
 NOR2_X4 _26589_ (.A1(_04033_),
    .A2(_04081_),
    .ZN(_04244_));
 NAND3_X1 _26590_ (.A1(_04048_),
    .A2(_04244_),
    .A3(_04091_),
    .ZN(_04245_));
 BUF_X4 _26591_ (.A(_04200_),
    .Z(_04246_));
 NAND3_X1 _26592_ (.A1(_04002_),
    .A2(_04246_),
    .A3(_04179_),
    .ZN(_04247_));
 NAND2_X1 _26593_ (.A1(_04245_),
    .A2(_04247_),
    .ZN(_04248_));
 AOI221_X2 _26594_ (.A(_04241_),
    .B1(_04243_),
    .B2(_04110_),
    .C1(_04191_),
    .C2(_04248_),
    .ZN(_04249_));
 NAND4_X2 _26595_ (.A1(_04205_),
    .A2(_04216_),
    .A3(_04232_),
    .A4(_04249_),
    .ZN(_04250_));
 NOR4_X4 _26596_ (.A1(_04089_),
    .A2(_04124_),
    .A3(_04196_),
    .A4(_04250_),
    .ZN(_04251_));
 AOI222_X2 _26597_ (.A1(\core.keymem.key_mem[7][120] ),
    .A2(_17084_),
    .B1(_16536_),
    .B2(\core.keymem.key_mem[9][120] ),
    .C1(\core.keymem.key_mem[12][120] ),
    .C2(_16398_),
    .ZN(_04252_));
 AOI22_X1 _26598_ (.A1(\core.keymem.key_mem[14][120] ),
    .A2(_16999_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][120] ),
    .ZN(_04253_));
 AOI22_X1 _26599_ (.A1(\core.keymem.key_mem[4][120] ),
    .A2(_18232_),
    .B1(_17768_),
    .B2(\core.keymem.key_mem[11][120] ),
    .ZN(_04254_));
 NAND3_X1 _26600_ (.A1(_04252_),
    .A2(_04253_),
    .A3(_04254_),
    .ZN(_04255_));
 AOI22_X1 _26601_ (.A1(\core.keymem.key_mem[3][120] ),
    .A2(_16987_),
    .B1(_17003_),
    .B2(\core.keymem.key_mem[1][120] ),
    .ZN(_04256_));
 AOI22_X1 _26602_ (.A1(\core.keymem.key_mem[2][120] ),
    .A2(_17786_),
    .B1(_16989_),
    .B2(\core.keymem.key_mem[10][120] ),
    .ZN(_04257_));
 AOI22_X1 _26603_ (.A1(\core.keymem.key_mem[6][120] ),
    .A2(_16521_),
    .B1(_17666_),
    .B2(\core.keymem.key_mem[8][120] ),
    .ZN(_04258_));
 AOI21_X1 _26604_ (.A(_16495_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][120] ),
    .ZN(_04259_));
 NAND4_X1 _26605_ (.A1(_04256_),
    .A2(_04257_),
    .A3(_04258_),
    .A4(_04259_),
    .ZN(_04260_));
 NOR2_X1 _26606_ (.A1(_04255_),
    .A2(_04260_),
    .ZN(_04261_));
 AOI21_X4 _26607_ (.A(_04261_),
    .B1(_16873_),
    .B2(_00177_),
    .ZN(_04262_));
 XNOR2_X2 _26608_ (.A(\core.dec_block.block_w0_reg[24] ),
    .B(_04262_),
    .ZN(_04263_));
 CLKBUF_X3 _26609_ (.A(_16554_),
    .Z(_04264_));
 XNOR2_X1 _26610_ (.A(\block_reg[0][24] ),
    .B(_04262_),
    .ZN(_04265_));
 BUF_X4 _26611_ (.A(_18552_),
    .Z(_04266_));
 OAI221_X1 _26612_ (.A(_04251_),
    .B1(_04263_),
    .B2(_04264_),
    .C1(_04265_),
    .C2(_04266_),
    .ZN(_04267_));
 AND2_X1 _26613_ (.A1(_00175_),
    .A2(_16545_),
    .ZN(_04268_));
 NAND3_X1 _26614_ (.A1(\core.keymem.key_mem[12][125] ),
    .A2(_17099_),
    .A3(_16893_),
    .ZN(_04269_));
 OAI211_X2 _26615_ (.A(\core.keymem.key_mem[1][125] ),
    .B(_16902_),
    .C1(_16913_),
    .C2(_16915_),
    .ZN(_04270_));
 NAND3_X1 _26616_ (.A1(\core.keymem.key_mem[2][125] ),
    .A2(_16902_),
    .A3(_16907_),
    .ZN(_04271_));
 OAI211_X2 _26617_ (.A(\core.keymem.key_mem[13][125] ),
    .B(_16919_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_04272_));
 NAND4_X2 _26618_ (.A1(_04269_),
    .A2(_04270_),
    .A3(_04271_),
    .A4(_04272_),
    .ZN(_04273_));
 OAI221_X2 _26619_ (.A(\core.keymem.key_mem[5][125] ),
    .B1(_16933_),
    .B2(_16934_),
    .C1(_17018_),
    .C2(_17020_),
    .ZN(_04274_));
 OAI211_X2 _26620_ (.A(\core.keymem.key_mem[7][125] ),
    .B(_16938_),
    .C1(_16933_),
    .C2(_16934_),
    .ZN(_04275_));
 NAND3_X1 _26621_ (.A1(\core.keymem.key_mem[14][125] ),
    .A2(_16881_),
    .A3(_17015_),
    .ZN(_04276_));
 OAI211_X2 _26622_ (.A(\core.keymem.key_mem[4][125] ),
    .B(_16921_),
    .C1(_16933_),
    .C2(_16934_),
    .ZN(_04277_));
 NAND4_X2 _26623_ (.A1(_04274_),
    .A2(_04275_),
    .A3(_04276_),
    .A4(_04277_),
    .ZN(_04278_));
 OAI211_X2 _26624_ (.A(\core.keymem.key_mem[6][125] ),
    .B(_17015_),
    .C1(_16934_),
    .C2(_16933_),
    .ZN(_04279_));
 OAI211_X2 _26625_ (.A(\core.keymem.key_mem[10][125] ),
    .B(_17025_),
    .C1(_16885_),
    .C2(_16889_),
    .ZN(_04280_));
 OAI221_X2 _26626_ (.A(\core.keymem.key_mem[9][125] ),
    .B1(_16926_),
    .B2(_16928_),
    .C1(_17018_),
    .C2(_17020_),
    .ZN(_04281_));
 OAI211_X2 _26627_ (.A(\core.keymem.key_mem[11][125] ),
    .B(_16938_),
    .C1(_16885_),
    .C2(_16889_),
    .ZN(_04282_));
 NAND4_X2 _26628_ (.A1(_04279_),
    .A2(_04280_),
    .A3(_04281_),
    .A4(_04282_),
    .ZN(_04283_));
 INV_X1 _26629_ (.A(\core.keymem.key_mem[8][125] ),
    .ZN(_04284_));
 INV_X1 _26630_ (.A(\core.keymem.key_mem[3][125] ),
    .ZN(_04285_));
 OAI22_X4 _26631_ (.A1(_04284_),
    .A2(_17134_),
    .B1(_17637_),
    .B2(_04285_),
    .ZN(_04286_));
 NOR4_X4 _26632_ (.A1(_04273_),
    .A2(_04278_),
    .A3(_04283_),
    .A4(_04286_),
    .ZN(_04287_));
 AOI21_X4 _26633_ (.A(_04268_),
    .B1(_04287_),
    .B2(_16487_),
    .ZN(_04288_));
 XNOR2_X2 _26634_ (.A(\core.dec_block.block_w0_reg[29] ),
    .B(_04288_),
    .ZN(_04289_));
 INV_X1 _26635_ (.A(\core.dec_block.block_w0_reg[30] ),
    .ZN(_04290_));
 OAI21_X1 _26636_ (.A(\core.keymem.key_mem[9][126] ),
    .B1(_17018_),
    .B2(_17020_),
    .ZN(_04291_));
 NAND2_X1 _26637_ (.A1(\core.keymem.key_mem[11][126] ),
    .A2(_16938_),
    .ZN(_04292_));
 AOI21_X1 _26638_ (.A(_17529_),
    .B1(_04291_),
    .B2(_04292_),
    .ZN(_04293_));
 OAI211_X2 _26639_ (.A(\core.keymem.key_mem[7][126] ),
    .B(_16481_),
    .C1(_16895_),
    .C2(_16898_),
    .ZN(_04294_));
 NAND3_X1 _26640_ (.A1(\core.keymem.key_mem[3][126] ),
    .A2(_16481_),
    .A3(_16969_),
    .ZN(_04295_));
 OAI211_X2 _26641_ (.A(\core.keymem.key_mem[8][126] ),
    .B(_16484_),
    .C1(_16926_),
    .C2(_16928_),
    .ZN(_04296_));
 OAI211_X2 _26642_ (.A(\core.keymem.key_mem[6][126] ),
    .B(_16906_),
    .C1(_16898_),
    .C2(_16895_),
    .ZN(_04297_));
 NAND4_X1 _26643_ (.A1(_04294_),
    .A2(_04295_),
    .A3(_04296_),
    .A4(_04297_),
    .ZN(_04298_));
 OAI211_X2 _26644_ (.A(\core.keymem.key_mem[4][126] ),
    .B(_16484_),
    .C1(_16895_),
    .C2(_16898_),
    .ZN(_04299_));
 OAI211_X2 _26645_ (.A(\core.keymem.key_mem[13][126] ),
    .B(_16478_),
    .C1(_16912_),
    .C2(_16914_),
    .ZN(_04300_));
 OAI211_X2 _26646_ (.A(\core.keymem.key_mem[10][126] ),
    .B(_16906_),
    .C1(_16884_),
    .C2(_16888_),
    .ZN(_04301_));
 NAND3_X1 _26647_ (.A1(\core.keymem.key_mem[14][126] ),
    .A2(_16478_),
    .A3(_16906_),
    .ZN(_04302_));
 NAND4_X1 _26648_ (.A1(_04299_),
    .A2(_04300_),
    .A3(_04301_),
    .A4(_04302_),
    .ZN(_04303_));
 OAI221_X1 _26649_ (.A(\core.keymem.key_mem[5][126] ),
    .B1(_16895_),
    .B2(_16897_),
    .C1(_16912_),
    .C2(_16914_),
    .ZN(_04304_));
 NAND3_X1 _26650_ (.A1(\core.keymem.key_mem[2][126] ),
    .A2(_16485_),
    .A3(_16906_),
    .ZN(_04305_));
 OAI211_X2 _26651_ (.A(\core.keymem.key_mem[1][126] ),
    .B(_16485_),
    .C1(_16912_),
    .C2(_16914_),
    .ZN(_04306_));
 NAND3_X1 _26652_ (.A1(\core.keymem.key_mem[12][126] ),
    .A2(_16478_),
    .A3(_16484_),
    .ZN(_04307_));
 NAND4_X1 _26653_ (.A1(_04304_),
    .A2(_04305_),
    .A3(_04306_),
    .A4(_04307_),
    .ZN(_04308_));
 NOR4_X2 _26654_ (.A1(_04293_),
    .A2(_04298_),
    .A3(_04303_),
    .A4(_04308_),
    .ZN(_04309_));
 MUX2_X2 _26655_ (.A(_00188_),
    .B(_04309_),
    .S(_16487_),
    .Z(_04310_));
 XNOR2_X2 _26656_ (.A(_04290_),
    .B(_04310_),
    .ZN(_04311_));
 XNOR2_X2 _26657_ (.A(_04289_),
    .B(_04311_),
    .ZN(_04312_));
 XNOR2_X2 _26658_ (.A(_18410_),
    .B(_04312_),
    .ZN(_04313_));
 XNOR2_X1 _26659_ (.A(_18478_),
    .B(_04313_),
    .ZN(_04314_));
 XNOR2_X1 _26660_ (.A(_18871_),
    .B(_03857_),
    .ZN(_04315_));
 XNOR2_X2 _26661_ (.A(_03976_),
    .B(_04315_),
    .ZN(_04316_));
 AOI21_X1 _26662_ (.A(_16494_),
    .B1(_17191_),
    .B2(\core.keymem.key_mem[14][104] ),
    .ZN(_04317_));
 AOI22_X1 _26663_ (.A1(\core.keymem.key_mem[4][104] ),
    .A2(_16456_),
    .B1(_17648_),
    .B2(\core.keymem.key_mem[6][104] ),
    .ZN(_04318_));
 AOI22_X1 _26664_ (.A1(\core.keymem.key_mem[9][104] ),
    .A2(_16535_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][104] ),
    .ZN(_04319_));
 AOI22_X1 _26665_ (.A1(\core.keymem.key_mem[3][104] ),
    .A2(_16865_),
    .B1(_16531_),
    .B2(\core.keymem.key_mem[13][104] ),
    .ZN(_04320_));
 AND4_X1 _26666_ (.A1(_04317_),
    .A2(_04318_),
    .A3(_04319_),
    .A4(_04320_),
    .ZN(_04321_));
 AOI222_X2 _26667_ (.A1(\core.keymem.key_mem[7][104] ),
    .A2(_16955_),
    .B1(_16858_),
    .B2(\core.keymem.key_mem[2][104] ),
    .C1(_16948_),
    .C2(\core.keymem.key_mem[5][104] ),
    .ZN(_04322_));
 AOI22_X1 _26668_ (.A1(\core.keymem.key_mem[8][104] ),
    .A2(_16528_),
    .B1(_16514_),
    .B2(\core.keymem.key_mem[10][104] ),
    .ZN(_04323_));
 AOI22_X1 _26669_ (.A1(\core.keymem.key_mem[11][104] ),
    .A2(_16505_),
    .B1(_16854_),
    .B2(\core.keymem.key_mem[1][104] ),
    .ZN(_04324_));
 AND3_X1 _26670_ (.A1(_04322_),
    .A2(_04323_),
    .A3(_04324_),
    .ZN(_04325_));
 AOI22_X4 _26671_ (.A1(_00182_),
    .A2(_16496_),
    .B1(_04321_),
    .B2(_04325_),
    .ZN(_04326_));
 XNOR2_X2 _26672_ (.A(\core.dec_block.block_w0_reg[8] ),
    .B(_04326_),
    .ZN(_04327_));
 AND2_X1 _26673_ (.A1(_00176_),
    .A2(_16982_),
    .ZN(_04328_));
 OAI211_X2 _26674_ (.A(\core.keymem.key_mem[11][127] ),
    .B(_17111_),
    .C1(_16886_),
    .C2(_16890_),
    .ZN(_04329_));
 OAI211_X2 _26675_ (.A(\core.keymem.key_mem[1][127] ),
    .B(_17120_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_04330_));
 OAI211_X2 _26676_ (.A(\core.keymem.key_mem[7][127] ),
    .B(_17074_),
    .C1(_17030_),
    .C2(_17031_),
    .ZN(_04331_));
 OAI211_X2 _26677_ (.A(\core.keymem.key_mem[6][127] ),
    .B(_17026_),
    .C1(_17622_),
    .C2(_17030_),
    .ZN(_04332_));
 NAND4_X2 _26678_ (.A1(_04329_),
    .A2(_04330_),
    .A3(_04331_),
    .A4(_04332_),
    .ZN(_04333_));
 OAI221_X2 _26679_ (.A(\core.keymem.key_mem[5][127] ),
    .B1(_16908_),
    .B2(_16917_),
    .C1(_16913_),
    .C2(_16915_),
    .ZN(_04334_));
 OAI221_X2 _26680_ (.A(\core.keymem.key_mem[9][127] ),
    .B1(_16885_),
    .B2(_16889_),
    .C1(_16913_),
    .C2(_16915_),
    .ZN(_04335_));
 NAND3_X1 _26681_ (.A1(\core.keymem.key_mem[2][127] ),
    .A2(_17827_),
    .A3(_17163_),
    .ZN(_04336_));
 OAI211_X2 _26682_ (.A(\core.keymem.key_mem[4][127] ),
    .B(_16893_),
    .C1(_16896_),
    .C2(_16899_),
    .ZN(_04337_));
 NAND4_X2 _26683_ (.A1(_04334_),
    .A2(_04335_),
    .A3(_04336_),
    .A4(_04337_),
    .ZN(_04338_));
 OAI211_X2 _26684_ (.A(\core.keymem.key_mem[10][127] ),
    .B(_17163_),
    .C1(_17035_),
    .C2(_17036_),
    .ZN(_04339_));
 NAND3_X1 _26685_ (.A1(\core.keymem.key_mem[12][127] ),
    .A2(_17099_),
    .A3(_16893_),
    .ZN(_04340_));
 OAI211_X2 _26686_ (.A(\core.keymem.key_mem[8][127] ),
    .B(_16931_),
    .C1(_16927_),
    .C2(_16929_),
    .ZN(_04341_));
 NAND3_X1 _26687_ (.A1(\core.keymem.key_mem[14][127] ),
    .A2(_16919_),
    .A3(_16907_),
    .ZN(_04342_));
 NAND4_X2 _26688_ (.A1(_04339_),
    .A2(_04340_),
    .A3(_04341_),
    .A4(_04342_),
    .ZN(_04343_));
 INV_X1 _26689_ (.A(\core.keymem.key_mem[3][127] ),
    .ZN(_04344_));
 INV_X1 _26690_ (.A(\core.keymem.key_mem[13][127] ),
    .ZN(_04345_));
 OAI22_X4 _26691_ (.A1(_04344_),
    .A2(_17637_),
    .B1(_17638_),
    .B2(_04345_),
    .ZN(_04346_));
 NOR4_X4 _26692_ (.A1(_04333_),
    .A2(_04338_),
    .A3(_04343_),
    .A4(_04346_),
    .ZN(_04347_));
 AOI21_X4 _26693_ (.A(_04328_),
    .B1(_04347_),
    .B2(_16488_),
    .ZN(_04348_));
 XNOR2_X2 _26694_ (.A(_04003_),
    .B(_04348_),
    .ZN(_04349_));
 XOR2_X1 _26695_ (.A(_04327_),
    .B(_04349_),
    .Z(_04350_));
 AOI22_X1 _26696_ (.A1(\core.keymem.key_mem[1][101] ),
    .A2(_16854_),
    .B1(_16531_),
    .B2(\core.keymem.key_mem[13][101] ),
    .ZN(_04351_));
 AOI22_X1 _26697_ (.A1(\core.keymem.key_mem[8][101] ),
    .A2(_16528_),
    .B1(_16948_),
    .B2(\core.keymem.key_mem[5][101] ),
    .ZN(_04352_));
 AOI22_X1 _26698_ (.A1(\core.keymem.key_mem[7][101] ),
    .A2(_16406_),
    .B1(_16423_),
    .B2(\core.keymem.key_mem[2][101] ),
    .ZN(_04353_));
 AOI21_X1 _26699_ (.A(_16544_),
    .B1(_16538_),
    .B2(\core.keymem.key_mem[12][101] ),
    .ZN(_04354_));
 AND4_X1 _26700_ (.A1(_04351_),
    .A2(_04352_),
    .A3(_04353_),
    .A4(_04354_),
    .ZN(_04355_));
 INV_X1 _26701_ (.A(\core.keymem.key_mem[10][101] ),
    .ZN(_04356_));
 AOI21_X1 _26702_ (.A(_04356_),
    .B1(_16427_),
    .B2(_16429_),
    .ZN(_04357_));
 MUX2_X1 _26703_ (.A(\core.keymem.key_mem[6][101] ),
    .B(\core.keymem.key_mem[14][101] ),
    .S(_16972_),
    .Z(_04358_));
 AND2_X1 _26704_ (.A1(_16961_),
    .A2(_04358_),
    .ZN(_04359_));
 OAI21_X1 _26705_ (.A(_17016_),
    .B1(_04357_),
    .B2(_04359_),
    .ZN(_04360_));
 AOI22_X1 _26706_ (.A1(\core.keymem.key_mem[4][101] ),
    .A2(_16456_),
    .B1(_16441_),
    .B2(\core.keymem.key_mem[11][101] ),
    .ZN(_04361_));
 AOI22_X1 _26707_ (.A1(\core.keymem.key_mem[3][101] ),
    .A2(_16865_),
    .B1(_16461_),
    .B2(\core.keymem.key_mem[9][101] ),
    .ZN(_04362_));
 AND3_X1 _26708_ (.A1(_04360_),
    .A2(_04361_),
    .A3(_04362_),
    .ZN(_04363_));
 AOI22_X4 _26709_ (.A1(_00183_),
    .A2(_16983_),
    .B1(_04355_),
    .B2(_04363_),
    .ZN(_04364_));
 XNOR2_X2 _26710_ (.A(\core.dec_block.block_w0_reg[5] ),
    .B(_04364_),
    .ZN(_04365_));
 XNOR2_X1 _26711_ (.A(_16551_),
    .B(_04365_),
    .ZN(_04366_));
 XNOR2_X1 _26712_ (.A(_04350_),
    .B(_04366_),
    .ZN(_04367_));
 XNOR2_X1 _26713_ (.A(_04316_),
    .B(_04367_),
    .ZN(_04368_));
 XNOR2_X1 _26714_ (.A(_04314_),
    .B(_04368_),
    .ZN(_04369_));
 BUF_X4 _26715_ (.A(_17748_),
    .Z(_04370_));
 AOI21_X1 _26716_ (.A(_04267_),
    .B1(_04369_),
    .B2(_04370_),
    .ZN(_04371_));
 AOI21_X1 _26717_ (.A(_03979_),
    .B1(_04371_),
    .B2(_16366_),
    .ZN(_00583_));
 INV_X1 _26718_ (.A(\core.dec_block.block_w0_reg[25] ),
    .ZN(_04372_));
 AOI22_X1 _26719_ (.A1(_04094_),
    .A2(_04207_),
    .B1(_04225_),
    .B2(_04034_),
    .ZN(_04373_));
 NAND3_X1 _26720_ (.A1(_04181_),
    .A2(_04094_),
    .A3(_04207_),
    .ZN(_04374_));
 AOI21_X1 _26721_ (.A(_04373_),
    .B1(_04374_),
    .B2(_04197_),
    .ZN(_04375_));
 NOR2_X4 _26722_ (.A1(_04033_),
    .A2(_04093_),
    .ZN(_04376_));
 AOI21_X1 _26723_ (.A(_04045_),
    .B1(_04029_),
    .B2(_04155_),
    .ZN(_04377_));
 AOI21_X1 _26724_ (.A(_04377_),
    .B1(_04148_),
    .B2(_04045_),
    .ZN(_04378_));
 MUX2_X1 _26725_ (.A(_04166_),
    .B(_04378_),
    .S(_04058_),
    .Z(_04379_));
 NOR3_X1 _26726_ (.A1(_04071_),
    .A2(_04376_),
    .A3(_04379_),
    .ZN(_04380_));
 BUF_X4 _26727_ (.A(_04099_),
    .Z(_04381_));
 AOI21_X1 _26728_ (.A(_04380_),
    .B1(_04381_),
    .B2(_04072_),
    .ZN(_04382_));
 NOR3_X1 _26729_ (.A1(_04086_),
    .A2(_04053_),
    .A3(_04033_),
    .ZN(_04383_));
 NAND3_X1 _26730_ (.A1(_04212_),
    .A2(_04024_),
    .A3(_04154_),
    .ZN(_04384_));
 OAI21_X1 _26731_ (.A(_04154_),
    .B1(_04024_),
    .B2(_04029_),
    .ZN(_04385_));
 NAND3_X1 _26732_ (.A1(_04046_),
    .A2(_04053_),
    .A3(_04385_),
    .ZN(_04386_));
 AOI21_X1 _26733_ (.A(_04008_),
    .B1(_04384_),
    .B2(_04386_),
    .ZN(_04387_));
 OAI21_X1 _26734_ (.A(_04091_),
    .B1(_04383_),
    .B2(_04387_),
    .ZN(_04388_));
 NAND2_X4 _26735_ (.A1(_04075_),
    .A2(_04051_),
    .ZN(_04389_));
 OAI21_X1 _26736_ (.A(_04042_),
    .B1(_04169_),
    .B2(_04073_),
    .ZN(_04390_));
 NOR3_X1 _26737_ (.A1(_04045_),
    .A2(_04389_),
    .A3(_04390_),
    .ZN(_04391_));
 AOI21_X1 _26738_ (.A(_04082_),
    .B1(_04156_),
    .B2(_04045_),
    .ZN(_04392_));
 OAI21_X1 _26739_ (.A(_04237_),
    .B1(_04392_),
    .B2(_04074_),
    .ZN(_04393_));
 AOI221_X2 _26740_ (.A(_04391_),
    .B1(_04161_),
    .B2(_04186_),
    .C1(_04070_),
    .C2(_04393_),
    .ZN(_04394_));
 NAND2_X1 _26741_ (.A1(_04388_),
    .A2(_04394_),
    .ZN(_04395_));
 NOR3_X1 _26742_ (.A1(_04111_),
    .A2(_04221_),
    .A3(_04127_),
    .ZN(_04396_));
 NAND2_X2 _26743_ (.A1(_04062_),
    .A2(_04054_),
    .ZN(_04397_));
 OAI22_X1 _26744_ (.A1(_04053_),
    .A2(_04033_),
    .B1(_04397_),
    .B2(_04146_),
    .ZN(_04398_));
 AOI21_X2 _26745_ (.A(_04396_),
    .B1(_04398_),
    .B2(_03989_),
    .ZN(_04399_));
 NOR2_X1 _26746_ (.A1(_04052_),
    .A2(_04049_),
    .ZN(_04400_));
 NOR2_X2 _26747_ (.A1(_04012_),
    .A2(_04154_),
    .ZN(_04401_));
 AOI221_X2 _26748_ (.A(_04008_),
    .B1(_04206_),
    .B2(_04400_),
    .C1(_04401_),
    .C2(_04040_),
    .ZN(_04402_));
 NAND2_X1 _26749_ (.A1(_04039_),
    .A2(_04062_),
    .ZN(_04403_));
 AOI221_X2 _26750_ (.A(_04402_),
    .B1(_04403_),
    .B2(_04008_),
    .C1(_04057_),
    .C2(_04128_),
    .ZN(_04404_));
 NAND2_X1 _26751_ (.A1(_04098_),
    .A2(_04054_),
    .ZN(_04405_));
 OAI21_X1 _26752_ (.A(_04405_),
    .B1(_04151_),
    .B2(_04397_),
    .ZN(_04406_));
 NAND2_X2 _26753_ (.A1(_04073_),
    .A2(_04069_),
    .ZN(_04407_));
 NAND2_X4 _26754_ (.A1(_04029_),
    .A2(_04091_),
    .ZN(_04408_));
 BUF_X4 _26755_ (.A(_04405_),
    .Z(_04409_));
 OAI22_X2 _26756_ (.A1(_04397_),
    .A2(_04407_),
    .B1(_04408_),
    .B2(_04409_),
    .ZN(_04410_));
 AOI221_X2 _26757_ (.A(_04404_),
    .B1(_04406_),
    .B2(_03988_),
    .C1(_04410_),
    .C2(_03995_),
    .ZN(_04411_));
 NAND2_X4 _26758_ (.A1(_03988_),
    .A2(_04044_),
    .ZN(_04412_));
 NOR2_X1 _26759_ (.A1(_04106_),
    .A2(_04412_),
    .ZN(_04413_));
 NAND2_X4 _26760_ (.A1(_04090_),
    .A2(_04150_),
    .ZN(_04414_));
 NAND2_X2 _26761_ (.A1(_04045_),
    .A2(_04090_),
    .ZN(_04415_));
 NAND2_X1 _26762_ (.A1(_04414_),
    .A2(_04415_),
    .ZN(_04416_));
 NOR2_X1 _26763_ (.A1(_04057_),
    .A2(_04077_),
    .ZN(_04417_));
 AOI21_X1 _26764_ (.A(_04176_),
    .B1(_04149_),
    .B2(_04057_),
    .ZN(_04418_));
 OR2_X1 _26765_ (.A1(_04417_),
    .A2(_04418_),
    .ZN(_04419_));
 AOI221_X2 _26766_ (.A(_04413_),
    .B1(_04416_),
    .B2(_04109_),
    .C1(_04419_),
    .C2(_04070_),
    .ZN(_04420_));
 NOR2_X2 _26767_ (.A1(_04025_),
    .A2(_04094_),
    .ZN(_04421_));
 OAI21_X4 _26768_ (.A(_04226_),
    .B1(_04421_),
    .B2(_04042_),
    .ZN(_04422_));
 NAND2_X1 _26769_ (.A1(_04013_),
    .A2(_04050_),
    .ZN(_04423_));
 AOI21_X1 _26770_ (.A(_04063_),
    .B1(_04423_),
    .B2(_04041_),
    .ZN(_04424_));
 AOI21_X1 _26771_ (.A(_04050_),
    .B1(_04023_),
    .B2(_04013_),
    .ZN(_04425_));
 OAI221_X2 _26772_ (.A(_04069_),
    .B1(_04013_),
    .B2(_04019_),
    .C1(_04425_),
    .C2(_04073_),
    .ZN(_04426_));
 OAI21_X1 _26773_ (.A(_04160_),
    .B1(_04206_),
    .B2(_04033_),
    .ZN(_04427_));
 AOI221_X2 _26774_ (.A(_04422_),
    .B1(_04424_),
    .B2(_04426_),
    .C1(_04064_),
    .C2(_04427_),
    .ZN(_04428_));
 NAND4_X2 _26775_ (.A1(_04399_),
    .A2(_04411_),
    .A3(_04420_),
    .A4(_04428_),
    .ZN(_04429_));
 NOR4_X2 _26776_ (.A1(_04124_),
    .A2(_04382_),
    .A3(_04395_),
    .A4(_04429_),
    .ZN(_04430_));
 NAND4_X1 _26777_ (.A1(_04229_),
    .A2(_04121_),
    .A3(_04212_),
    .A4(_04117_),
    .ZN(_04431_));
 AOI21_X1 _26778_ (.A(_04075_),
    .B1(_04105_),
    .B2(_03994_),
    .ZN(_04432_));
 NOR3_X1 _26779_ (.A1(_04001_),
    .A2(_04117_),
    .A3(_04432_),
    .ZN(_04433_));
 NAND2_X1 _26780_ (.A1(_04121_),
    .A2(_04117_),
    .ZN(_04434_));
 OAI21_X1 _26781_ (.A(_04434_),
    .B1(_04117_),
    .B2(_04014_),
    .ZN(_04435_));
 AOI21_X1 _26782_ (.A(_04433_),
    .B1(_04435_),
    .B2(_04047_),
    .ZN(_04436_));
 AOI21_X1 _26783_ (.A(_04050_),
    .B1(_04431_),
    .B2(_04436_),
    .ZN(_04437_));
 NOR3_X1 _26784_ (.A1(_04212_),
    .A2(_04125_),
    .A3(_04434_),
    .ZN(_04438_));
 OAI21_X1 _26785_ (.A(_04179_),
    .B1(_04437_),
    .B2(_04438_),
    .ZN(_04439_));
 AOI21_X1 _26786_ (.A(_04166_),
    .B1(_04094_),
    .B2(_04191_),
    .ZN(_04440_));
 BUF_X4 _26787_ (.A(_04160_),
    .Z(_04441_));
 NOR3_X1 _26788_ (.A1(_04086_),
    .A2(_04081_),
    .A3(_04403_),
    .ZN(_04442_));
 NAND3_X1 _26789_ (.A1(_04121_),
    .A2(_04024_),
    .A3(_04154_),
    .ZN(_04443_));
 OAI21_X1 _26790_ (.A(_04443_),
    .B1(_04051_),
    .B2(_04121_),
    .ZN(_04444_));
 NAND2_X1 _26791_ (.A1(_03995_),
    .A2(_04121_),
    .ZN(_04445_));
 OAI22_X1 _26792_ (.A1(_04142_),
    .A2(_04444_),
    .B1(_04445_),
    .B2(_04154_),
    .ZN(_04446_));
 AOI21_X1 _26793_ (.A(_04442_),
    .B1(_04446_),
    .B2(_04053_),
    .ZN(_04447_));
 OAI221_X2 _26794_ (.A(_04439_),
    .B1(_04440_),
    .B2(_04441_),
    .C1(_04447_),
    .C2(_04198_),
    .ZN(_04448_));
 INV_X1 _26795_ (.A(_04448_),
    .ZN(_04449_));
 AOI21_X2 _26796_ (.A(_04375_),
    .B1(_04430_),
    .B2(_04449_),
    .ZN(_04450_));
 BUF_X4 _26797_ (.A(_04047_),
    .Z(_04451_));
 BUF_X4 _26798_ (.A(_04048_),
    .Z(_04452_));
 NOR3_X1 _26799_ (.A1(_04451_),
    .A2(_04452_),
    .A3(_04409_),
    .ZN(_04453_));
 OAI21_X1 _26800_ (.A(_03989_),
    .B1(_04239_),
    .B2(_04453_),
    .ZN(_04454_));
 NOR2_X1 _26801_ (.A1(_04182_),
    .A2(_04188_),
    .ZN(_04455_));
 OAI21_X1 _26802_ (.A(_04166_),
    .B1(_04219_),
    .B2(_04455_),
    .ZN(_04456_));
 NAND2_X4 _26803_ (.A1(_03995_),
    .A2(_04206_),
    .ZN(_04457_));
 NOR2_X1 _26804_ (.A1(_04065_),
    .A2(_04457_),
    .ZN(_04458_));
 NAND2_X4 _26805_ (.A1(_04044_),
    .A2(_04000_),
    .ZN(_04459_));
 NOR2_X2 _26806_ (.A1(_04042_),
    .A2(_04459_),
    .ZN(_04460_));
 NOR2_X4 _26807_ (.A1(_04154_),
    .A2(_04135_),
    .ZN(_04461_));
 NOR2_X4 _26808_ (.A1(_04014_),
    .A2(_04154_),
    .ZN(_04462_));
 NOR2_X2 _26809_ (.A1(_04042_),
    .A2(_04129_),
    .ZN(_04463_));
 AOI221_X2 _26810_ (.A(_04458_),
    .B1(_04460_),
    .B2(_04461_),
    .C1(_04462_),
    .C2(_04463_),
    .ZN(_04464_));
 AND4_X2 _26811_ (.A1(_04450_),
    .A2(_04454_),
    .A3(_04456_),
    .A4(_04464_),
    .ZN(_04465_));
 CLKBUF_X3 _26812_ (.A(_04115_),
    .Z(_04466_));
 CLKBUF_X3 _26813_ (.A(_04143_),
    .Z(_04467_));
 AOI21_X1 _26814_ (.A(_04466_),
    .B1(_04459_),
    .B2(_04467_),
    .ZN(_04468_));
 OAI21_X1 _26815_ (.A(_04169_),
    .B1(_04181_),
    .B2(_04467_),
    .ZN(_04469_));
 BUF_X4 _26816_ (.A(_04132_),
    .Z(_04470_));
 AOI21_X1 _26817_ (.A(_04468_),
    .B1(_04469_),
    .B2(_04470_),
    .ZN(_04471_));
 NOR2_X1 _26818_ (.A1(_04107_),
    .A2(_04471_),
    .ZN(_04472_));
 AOI21_X1 _26819_ (.A(_04183_),
    .B1(_04461_),
    .B2(_04197_),
    .ZN(_04473_));
 AOI21_X1 _26820_ (.A(_04179_),
    .B1(_04219_),
    .B2(_04050_),
    .ZN(_04474_));
 OAI33_X1 _26821_ (.A1(_04181_),
    .A2(_04182_),
    .A3(_04473_),
    .B1(_04474_),
    .B2(_04135_),
    .B3(_04032_),
    .ZN(_04475_));
 NOR2_X1 _26822_ (.A1(_04127_),
    .A2(_04408_),
    .ZN(_04476_));
 OAI33_X1 _26823_ (.A1(_04014_),
    .A2(_04033_),
    .A3(_04222_),
    .B1(_04188_),
    .B2(_04176_),
    .B3(_04182_),
    .ZN(_04477_));
 BUF_X4 _26824_ (.A(_04397_),
    .Z(_04478_));
 NAND2_X4 _26825_ (.A1(_04000_),
    .A2(_04162_),
    .ZN(_04479_));
 AOI21_X1 _26826_ (.A(_04478_),
    .B1(_04457_),
    .B2(_04479_),
    .ZN(_04480_));
 OR4_X1 _26827_ (.A1(_04413_),
    .A2(_04476_),
    .A3(_04477_),
    .A4(_04480_),
    .ZN(_04481_));
 BUF_X4 _26828_ (.A(_04407_),
    .Z(_04482_));
 OAI33_X1 _26829_ (.A1(_04192_),
    .A2(_04112_),
    .A3(_04482_),
    .B1(_04408_),
    .B2(_04104_),
    .B3(_04046_),
    .ZN(_04483_));
 INV_X1 _26830_ (.A(_04483_),
    .ZN(_04484_));
 OAI21_X4 _26831_ (.A(_04484_),
    .B1(_04479_),
    .B2(_04065_),
    .ZN(_04485_));
 NOR4_X2 _26832_ (.A1(_04472_),
    .A2(_04475_),
    .A3(_04481_),
    .A4(_04485_),
    .ZN(_04486_));
 NOR4_X1 _26833_ (.A1(_04058_),
    .A2(_03996_),
    .A3(_04002_),
    .A4(_04174_),
    .ZN(_04487_));
 AOI21_X1 _26834_ (.A(_04487_),
    .B1(_04078_),
    .B2(_04132_),
    .ZN(_04488_));
 NOR2_X1 _26835_ (.A1(_04466_),
    .A2(_04488_),
    .ZN(_04489_));
 NAND2_X2 _26836_ (.A1(_04188_),
    .A2(_04207_),
    .ZN(_04490_));
 OAI22_X1 _26837_ (.A1(_04148_),
    .A2(_04412_),
    .B1(_04490_),
    .B2(_04127_),
    .ZN(_04491_));
 AOI21_X1 _26838_ (.A(_04491_),
    .B1(_04219_),
    .B2(_04110_),
    .ZN(_04492_));
 NOR2_X1 _26839_ (.A1(_04244_),
    .A2(_04461_),
    .ZN(_04493_));
 NAND2_X2 _26840_ (.A1(_03996_),
    .A2(_04091_),
    .ZN(_04494_));
 AOI21_X1 _26841_ (.A(_04139_),
    .B1(_04150_),
    .B2(_04094_),
    .ZN(_04495_));
 OAI221_X2 _26842_ (.A(_04492_),
    .B1(_04493_),
    .B2(_04457_),
    .C1(_04494_),
    .C2(_04495_),
    .ZN(_04496_));
 AOI21_X1 _26843_ (.A(_04139_),
    .B1(_04156_),
    .B2(_04452_),
    .ZN(_04497_));
 NOR2_X1 _26844_ (.A1(_04132_),
    .A2(_04497_),
    .ZN(_04498_));
 OAI21_X1 _26845_ (.A(_04467_),
    .B1(_04133_),
    .B2(_04498_),
    .ZN(_04499_));
 BUF_X4 _26846_ (.A(_04084_),
    .Z(_04500_));
 CLKBUF_X3 _26847_ (.A(_04229_),
    .Z(_04501_));
 NAND4_X1 _26848_ (.A1(_04500_),
    .A2(_04470_),
    .A3(_04501_),
    .A4(_04139_),
    .ZN(_04502_));
 AOI21_X2 _26849_ (.A(_04466_),
    .B1(_04499_),
    .B2(_04502_),
    .ZN(_04503_));
 NOR3_X4 _26850_ (.A1(_04489_),
    .A2(_04496_),
    .A3(_04503_),
    .ZN(_04504_));
 AOI221_X2 _26851_ (.A(_04133_),
    .B1(_04157_),
    .B2(_04229_),
    .C1(_03986_),
    .C2(_18416_),
    .ZN(_04505_));
 AOI21_X1 _26852_ (.A(_04505_),
    .B1(_04165_),
    .B2(_04072_),
    .ZN(_04506_));
 NAND3_X1 _26853_ (.A1(_04467_),
    .A2(_04197_),
    .A3(_04506_),
    .ZN(_04507_));
 AOI21_X2 _26854_ (.A(_04148_),
    .B1(_04414_),
    .B2(_04490_),
    .ZN(_04508_));
 NOR2_X1 _26855_ (.A1(_04193_),
    .A2(_04479_),
    .ZN(_04509_));
 NOR2_X2 _26856_ (.A1(_03994_),
    .A2(_04028_),
    .ZN(_04510_));
 NAND2_X2 _26857_ (.A1(_04206_),
    .A2(_04510_),
    .ZN(_04511_));
 OAI22_X2 _26858_ (.A1(_04055_),
    .A2(_04490_),
    .B1(_04511_),
    .B2(_04077_),
    .ZN(_04512_));
 NOR2_X1 _26859_ (.A1(_04111_),
    .A2(_04459_),
    .ZN(_04513_));
 NAND2_X1 _26860_ (.A1(_04110_),
    .A2(_04513_),
    .ZN(_04514_));
 OAI221_X2 _26861_ (.A(_04514_),
    .B1(_04408_),
    .B2(_04107_),
    .C1(_04397_),
    .C2(_04414_),
    .ZN(_04515_));
 NOR4_X4 _26862_ (.A1(_04508_),
    .A2(_04509_),
    .A3(_04512_),
    .A4(_04515_),
    .ZN(_04516_));
 NAND3_X1 _26863_ (.A1(_04163_),
    .A2(_04507_),
    .A3(_04516_),
    .ZN(_04517_));
 NAND2_X1 _26864_ (.A1(_04001_),
    .A2(_04137_),
    .ZN(_04518_));
 OAI21_X1 _26865_ (.A(_04511_),
    .B1(_04518_),
    .B2(_04441_),
    .ZN(_04519_));
 OAI21_X1 _26866_ (.A(_04519_),
    .B1(_04166_),
    .B2(_04137_),
    .ZN(_04520_));
 AOI21_X1 _26867_ (.A(_04174_),
    .B1(_04457_),
    .B2(_04441_),
    .ZN(_04521_));
 NAND2_X2 _26868_ (.A1(_03989_),
    .A2(_04191_),
    .ZN(_04522_));
 NOR2_X1 _26869_ (.A1(_04522_),
    .A2(_04127_),
    .ZN(_04523_));
 OAI21_X1 _26870_ (.A(_04181_),
    .B1(_04521_),
    .B2(_04523_),
    .ZN(_04524_));
 MUX2_X1 _26871_ (.A(_04068_),
    .B(_04459_),
    .S(_04212_),
    .Z(_04525_));
 OAI22_X1 _26872_ (.A1(_04501_),
    .A2(_04081_),
    .B1(_04525_),
    .B2(_04121_),
    .ZN(_04526_));
 NAND3_X1 _26873_ (.A1(_04098_),
    .A2(_04207_),
    .A3(_04526_),
    .ZN(_04527_));
 AOI21_X1 _26874_ (.A(_04412_),
    .B1(_04095_),
    .B2(_04065_),
    .ZN(_04528_));
 OAI22_X1 _26875_ (.A1(_04192_),
    .A2(_04441_),
    .B1(_04182_),
    .B2(_04193_),
    .ZN(_04529_));
 AOI21_X2 _26876_ (.A(_04528_),
    .B1(_04529_),
    .B2(_04150_),
    .ZN(_04530_));
 NAND4_X2 _26877_ (.A1(_04520_),
    .A2(_04524_),
    .A3(_04527_),
    .A4(_04530_),
    .ZN(_04531_));
 AOI21_X1 _26878_ (.A(_04164_),
    .B1(_04165_),
    .B2(_04061_),
    .ZN(_04532_));
 NOR2_X2 _26879_ (.A1(_04059_),
    .A2(_04229_),
    .ZN(_04533_));
 AOI21_X1 _26880_ (.A(_04532_),
    .B1(_04533_),
    .B2(_04244_),
    .ZN(_04534_));
 OAI21_X1 _26881_ (.A(_04399_),
    .B1(_04534_),
    .B2(_04500_),
    .ZN(_04535_));
 NOR3_X2 _26882_ (.A1(_04517_),
    .A2(_04531_),
    .A3(_04535_),
    .ZN(_04536_));
 NAND4_X2 _26883_ (.A1(_04465_),
    .A2(_04486_),
    .A3(_04504_),
    .A4(_04536_),
    .ZN(_04537_));
 NAND2_X4 _26884_ (.A1(_18416_),
    .A2(_04537_),
    .ZN(_04538_));
 INV_X1 _26885_ (.A(\block_reg[0][25] ),
    .ZN(_04539_));
 NAND2_X1 _26886_ (.A1(_00189_),
    .A2(_16498_),
    .ZN(_04540_));
 AOI22_X1 _26887_ (.A1(\core.keymem.key_mem[12][121] ),
    .A2(_16399_),
    .B1(_17675_),
    .B2(\core.keymem.key_mem[5][121] ),
    .ZN(_04541_));
 AOI22_X1 _26888_ (.A1(\core.keymem.key_mem[14][121] ),
    .A2(_16439_),
    .B1(_16991_),
    .B2(\core.keymem.key_mem[6][121] ),
    .ZN(_04542_));
 AOI22_X1 _26889_ (.A1(\core.keymem.key_mem[1][121] ),
    .A2(_16417_),
    .B1(_16473_),
    .B2(\core.keymem.key_mem[13][121] ),
    .ZN(_04543_));
 AOI22_X1 _26890_ (.A1(\core.keymem.key_mem[7][121] ),
    .A2(_16408_),
    .B1(_17781_),
    .B2(\core.keymem.key_mem[8][121] ),
    .ZN(_04544_));
 AND4_X1 _26891_ (.A1(_04541_),
    .A2(_04542_),
    .A3(_04543_),
    .A4(_04544_),
    .ZN(_04545_));
 AOI22_X2 _26892_ (.A1(\core.keymem.key_mem[2][121] ),
    .A2(_17086_),
    .B1(_17082_),
    .B2(\core.keymem.key_mem[10][121] ),
    .ZN(_04546_));
 AOI22_X2 _26893_ (.A1(\core.keymem.key_mem[3][121] ),
    .A2(_17091_),
    .B1(_17585_),
    .B2(\core.keymem.key_mem[9][121] ),
    .ZN(_04547_));
 AOI22_X2 _26894_ (.A1(\core.keymem.key_mem[4][121] ),
    .A2(_16501_),
    .B1(_17769_),
    .B2(\core.keymem.key_mem[11][121] ),
    .ZN(_04548_));
 NAND4_X2 _26895_ (.A1(_04545_),
    .A2(_04546_),
    .A3(_04547_),
    .A4(_04548_),
    .ZN(_04549_));
 OAI21_X4 _26896_ (.A(_04540_),
    .B1(_04549_),
    .B2(_17578_),
    .ZN(_04550_));
 XNOR2_X1 _26897_ (.A(_04539_),
    .B(_04550_),
    .ZN(_04551_));
 XNOR2_X2 _26898_ (.A(_04372_),
    .B(_04550_),
    .ZN(_04552_));
 OAI221_X1 _26899_ (.A(_16364_),
    .B1(_18078_),
    .B2(_04551_),
    .C1(_04552_),
    .C2(_19180_),
    .ZN(_04553_));
 AOI21_X1 _26900_ (.A(_16544_),
    .B1(_16954_),
    .B2(\core.keymem.key_mem[7][105] ),
    .ZN(_04554_));
 AOI22_X1 _26901_ (.A1(\core.keymem.key_mem[4][105] ),
    .A2(_16455_),
    .B1(_16466_),
    .B2(\core.keymem.key_mem[5][105] ),
    .ZN(_04555_));
 AOI22_X1 _26902_ (.A1(\core.keymem.key_mem[3][105] ),
    .A2(_16864_),
    .B1(_16523_),
    .B2(\core.keymem.key_mem[1][105] ),
    .ZN(_04556_));
 AOI22_X1 _26903_ (.A1(\core.keymem.key_mem[12][105] ),
    .A2(_16396_),
    .B1(_16470_),
    .B2(\core.keymem.key_mem[13][105] ),
    .ZN(_04557_));
 AND4_X1 _26904_ (.A1(_04554_),
    .A2(_04555_),
    .A3(_04556_),
    .A4(_04557_),
    .ZN(_04558_));
 AOI222_X2 _26905_ (.A1(\core.keymem.key_mem[2][105] ),
    .A2(_16858_),
    .B1(_16460_),
    .B2(\core.keymem.key_mem[9][105] ),
    .C1(\core.keymem.key_mem[11][105] ),
    .C2(_16440_),
    .ZN(_04559_));
 AOI22_X1 _26906_ (.A1(\core.keymem.key_mem[14][105] ),
    .A2(_16436_),
    .B1(_16431_),
    .B2(\core.keymem.key_mem[10][105] ),
    .ZN(_04560_));
 AOI22_X1 _26907_ (.A1(\core.keymem.key_mem[6][105] ),
    .A2(_16519_),
    .B1(_16450_),
    .B2(\core.keymem.key_mem[8][105] ),
    .ZN(_04561_));
 AND3_X1 _26908_ (.A1(_04559_),
    .A2(_04560_),
    .A3(_04561_),
    .ZN(_04562_));
 AOI22_X4 _26909_ (.A1(_00193_),
    .A2(_16495_),
    .B1(_04558_),
    .B2(_04562_),
    .ZN(_04563_));
 XOR2_X2 _26910_ (.A(\core.dec_block.block_w0_reg[9] ),
    .B(_04563_),
    .Z(_04564_));
 XOR2_X1 _26911_ (.A(_18410_),
    .B(_04564_),
    .Z(_04565_));
 XNOR2_X1 _26912_ (.A(_18550_),
    .B(_04565_),
    .ZN(_04566_));
 AND2_X1 _26913_ (.A1(_00184_),
    .A2(_16545_),
    .ZN(_04567_));
 NAND3_X1 _26914_ (.A1(\core.keymem.key_mem[2][102] ),
    .A2(_17827_),
    .A3(_17026_),
    .ZN(_04568_));
 NAND3_X1 _26915_ (.A1(\core.keymem.key_mem[3][102] ),
    .A2(_17074_),
    .A3(_17827_),
    .ZN(_04569_));
 OAI211_X2 _26916_ (.A(\core.keymem.key_mem[4][102] ),
    .B(_16893_),
    .C1(_17030_),
    .C2(_16899_),
    .ZN(_04570_));
 OAI211_X2 _26917_ (.A(\core.keymem.key_mem[6][102] ),
    .B(_17163_),
    .C1(_17031_),
    .C2(_16896_),
    .ZN(_04571_));
 NAND4_X2 _26918_ (.A1(_04568_),
    .A2(_04569_),
    .A3(_04570_),
    .A4(_04571_),
    .ZN(_04572_));
 OAI211_X2 _26919_ (.A(\core.keymem.key_mem[11][102] ),
    .B(_16901_),
    .C1(_16927_),
    .C2(_16929_),
    .ZN(_04573_));
 OAI211_X2 _26920_ (.A(\core.keymem.key_mem[7][102] ),
    .B(_16901_),
    .C1(_16896_),
    .C2(_16917_),
    .ZN(_04574_));
 OAI211_X2 _26921_ (.A(\core.keymem.key_mem[13][102] ),
    .B(_16919_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_04575_));
 OAI211_X2 _26922_ (.A(\core.keymem.key_mem[8][102] ),
    .B(_16931_),
    .C1(_16922_),
    .C2(_16923_),
    .ZN(_04576_));
 NAND4_X2 _26923_ (.A1(_04573_),
    .A2(_04574_),
    .A3(_04575_),
    .A4(_04576_),
    .ZN(_04577_));
 OAI221_X2 _26924_ (.A(\core.keymem.key_mem[9][102] ),
    .B1(_16926_),
    .B2(_16928_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_04578_));
 OAI211_X2 _26925_ (.A(\core.keymem.key_mem[1][102] ),
    .B(_16969_),
    .C1(_16935_),
    .C2(_16936_),
    .ZN(_04579_));
 NAND3_X1 _26926_ (.A1(\core.keymem.key_mem[12][102] ),
    .A2(_16881_),
    .A3(_16921_),
    .ZN(_04580_));
 OAI211_X2 _26927_ (.A(\core.keymem.key_mem[10][102] ),
    .B(_17015_),
    .C1(_16885_),
    .C2(_16889_),
    .ZN(_04581_));
 NAND4_X2 _26928_ (.A1(_04578_),
    .A2(_04579_),
    .A3(_04580_),
    .A4(_04581_),
    .ZN(_04582_));
 INV_X1 _26929_ (.A(\core.keymem.key_mem[14][102] ),
    .ZN(_04583_));
 NAND2_X1 _26930_ (.A1(_16919_),
    .A2(_17015_),
    .ZN(_04584_));
 INV_X1 _26931_ (.A(\core.keymem.key_mem[5][102] ),
    .ZN(_04585_));
 OAI22_X4 _26932_ (.A1(_04583_),
    .A2(_04584_),
    .B1(_03591_),
    .B2(_04585_),
    .ZN(_04586_));
 NOR4_X4 _26933_ (.A1(_04572_),
    .A2(_04577_),
    .A3(_04582_),
    .A4(_04586_),
    .ZN(_04587_));
 AOI21_X4 _26934_ (.A(_04567_),
    .B1(_04587_),
    .B2(_16487_),
    .ZN(_04588_));
 XNOR2_X2 _26935_ (.A(\core.dec_block.block_w0_reg[6] ),
    .B(_04588_),
    .ZN(_04589_));
 XNOR2_X2 _26936_ (.A(_04365_),
    .B(_04589_),
    .ZN(_04590_));
 XNOR2_X2 _26937_ (.A(_03510_),
    .B(_04590_),
    .ZN(_04591_));
 XNOR2_X1 _26938_ (.A(_04566_),
    .B(_04591_),
    .ZN(_04592_));
 XNOR2_X2 _26939_ (.A(_19192_),
    .B(_03915_),
    .ZN(_04593_));
 XNOR2_X1 _26940_ (.A(_04263_),
    .B(_04289_),
    .ZN(_04594_));
 XOR2_X1 _26941_ (.A(_04593_),
    .B(_04594_),
    .Z(_04595_));
 XNOR2_X1 _26942_ (.A(_04316_),
    .B(_04595_),
    .ZN(_04596_));
 XNOR2_X1 _26943_ (.A(_04592_),
    .B(_04596_),
    .ZN(_04597_));
 AOI21_X1 _26944_ (.A(_04553_),
    .B1(_04597_),
    .B2(_18332_),
    .ZN(_04598_));
 AOI22_X1 _26945_ (.A1(_04372_),
    .A2(_17744_),
    .B1(_04538_),
    .B2(_04598_),
    .ZN(_00584_));
 OAI221_X2 _26946_ (.A(_04193_),
    .B1(_04459_),
    .B2(_04478_),
    .C1(_04389_),
    .C2(_04451_),
    .ZN(_04599_));
 NAND2_X1 _26947_ (.A1(_04073_),
    .A2(_04083_),
    .ZN(_04600_));
 OAI22_X1 _26948_ (.A1(_04600_),
    .A2(_04060_),
    .B1(_04107_),
    .B2(_04242_),
    .ZN(_04601_));
 AOI22_X2 _26949_ (.A1(_03989_),
    .A2(_04599_),
    .B1(_04601_),
    .B2(_04470_),
    .ZN(_04602_));
 NAND2_X1 _26950_ (.A1(_04445_),
    .A2(_04401_),
    .ZN(_04603_));
 NOR3_X1 _26951_ (.A1(_04048_),
    .A2(_04212_),
    .A3(_04019_),
    .ZN(_04604_));
 OAI21_X1 _26952_ (.A(_04117_),
    .B1(_04400_),
    .B2(_04604_),
    .ZN(_04605_));
 OAI21_X1 _26953_ (.A(_04603_),
    .B1(_04605_),
    .B2(_04445_),
    .ZN(_04606_));
 AOI22_X2 _26954_ (.A1(_04501_),
    .A2(_04103_),
    .B1(_04207_),
    .B2(_04606_),
    .ZN(_04607_));
 NAND3_X2 _26955_ (.A1(_04394_),
    .A2(_04602_),
    .A3(_04607_),
    .ZN(_04608_));
 OAI22_X2 _26956_ (.A1(_04193_),
    .A2(_04414_),
    .B1(_04223_),
    .B2(_04457_),
    .ZN(_04609_));
 NOR3_X1 _26957_ (.A1(_04047_),
    .A2(_04148_),
    .A3(_04408_),
    .ZN(_04610_));
 NOR3_X1 _26958_ (.A1(_04043_),
    .A2(_03995_),
    .A3(_04237_),
    .ZN(_04611_));
 NOR3_X2 _26959_ (.A1(_04609_),
    .A2(_04610_),
    .A3(_04611_),
    .ZN(_04612_));
 NAND2_X1 _26960_ (.A1(_04530_),
    .A2(_04612_),
    .ZN(_04613_));
 BUF_X4 _26961_ (.A(_04229_),
    .Z(_04614_));
 AOI21_X2 _26962_ (.A(_04202_),
    .B1(_04186_),
    .B2(_04614_),
    .ZN(_04615_));
 AOI21_X1 _26963_ (.A(_04002_),
    .B1(_04441_),
    .B2(_04457_),
    .ZN(_04616_));
 AOI21_X2 _26964_ (.A(_04616_),
    .B1(_04101_),
    .B2(_04229_),
    .ZN(_04617_));
 OAI22_X4 _26965_ (.A1(_04412_),
    .A2(_04615_),
    .B1(_04617_),
    .B2(_04127_),
    .ZN(_04618_));
 NOR2_X1 _26966_ (.A1(_04129_),
    .A2(_04482_),
    .ZN(_04619_));
 OAI21_X1 _26967_ (.A(_04619_),
    .B1(_04137_),
    .B2(_04083_),
    .ZN(_04620_));
 OAI221_X1 _26968_ (.A(_04620_),
    .B1(_04222_),
    .B2(_04409_),
    .C1(_04478_),
    .C2(_04494_),
    .ZN(_04621_));
 OAI221_X1 _26969_ (.A(_04415_),
    .B1(_04482_),
    .B2(_04459_),
    .C1(_04151_),
    .C2(_04043_),
    .ZN(_04622_));
 AOI21_X1 _26970_ (.A(_04621_),
    .B1(_04622_),
    .B2(_04157_),
    .ZN(_04623_));
 NOR3_X1 _26971_ (.A1(_04025_),
    .A2(_04139_),
    .A3(_04156_),
    .ZN(_04624_));
 AOI21_X1 _26972_ (.A(_04113_),
    .B1(_04139_),
    .B2(_04460_),
    .ZN(_04625_));
 MUX2_X1 _26973_ (.A(_04192_),
    .B(_04127_),
    .S(_04614_),
    .Z(_04626_));
 OAI221_X2 _26974_ (.A(_04623_),
    .B1(_04624_),
    .B2(_04625_),
    .C1(_04626_),
    .C2(_04522_),
    .ZN(_04627_));
 NOR4_X4 _26975_ (.A1(_04608_),
    .A2(_04613_),
    .A3(_04618_),
    .A4(_04627_),
    .ZN(_04628_));
 NAND2_X1 _26976_ (.A1(_04002_),
    .A2(_04025_),
    .ZN(_04629_));
 NAND2_X1 _26977_ (.A1(_04001_),
    .A2(_04200_),
    .ZN(_04630_));
 NOR2_X1 _26978_ (.A1(_04068_),
    .A2(_04156_),
    .ZN(_04631_));
 AOI221_X2 _26979_ (.A(_04043_),
    .B1(_04068_),
    .B2(_04629_),
    .C1(_04630_),
    .C2(_04631_),
    .ZN(_04632_));
 NAND3_X1 _26980_ (.A1(_04132_),
    .A2(_04501_),
    .A3(_04246_),
    .ZN(_04633_));
 INV_X1 _26981_ (.A(_04133_),
    .ZN(_04634_));
 AOI21_X2 _26982_ (.A(_04482_),
    .B1(_04633_),
    .B2(_04634_),
    .ZN(_04635_));
 OR2_X1 _26983_ (.A1(_04409_),
    .A2(_04412_),
    .ZN(_04636_));
 OAI21_X2 _26984_ (.A(_04636_),
    .B1(_04415_),
    .B2(_04193_),
    .ZN(_04637_));
 NOR4_X4 _26985_ (.A1(_04234_),
    .A2(_04632_),
    .A3(_04635_),
    .A4(_04637_),
    .ZN(_04638_));
 AOI21_X1 _26986_ (.A(_04029_),
    .B1(_04389_),
    .B2(_04107_),
    .ZN(_04639_));
 OAI21_X1 _26987_ (.A(_04047_),
    .B1(_04138_),
    .B2(_04639_),
    .ZN(_04640_));
 NAND2_X1 _26988_ (.A1(_04002_),
    .A2(_04138_),
    .ZN(_04641_));
 AOI21_X2 _26989_ (.A(_04441_),
    .B1(_04640_),
    .B2(_04641_),
    .ZN(_04642_));
 AOI21_X1 _26990_ (.A(_04143_),
    .B1(_04181_),
    .B2(_04246_),
    .ZN(_04643_));
 NOR3_X1 _26991_ (.A1(_04500_),
    .A2(_04110_),
    .A3(_04137_),
    .ZN(_04644_));
 OAI33_X1 _26992_ (.A1(_04181_),
    .A2(_04441_),
    .A3(_04381_),
    .B1(_04643_),
    .B2(_04644_),
    .B3(_04466_),
    .ZN(_04645_));
 AOI21_X2 _26993_ (.A(_04642_),
    .B1(_04645_),
    .B2(_04197_),
    .ZN(_04646_));
 OAI22_X1 _26994_ (.A1(_04222_),
    .A2(_04381_),
    .B1(_04237_),
    .B2(_04479_),
    .ZN(_04647_));
 NAND3_X1 _26995_ (.A1(_04094_),
    .A2(_04179_),
    .A3(_04151_),
    .ZN(_04648_));
 OAI221_X2 _26996_ (.A(_04648_),
    .B1(_04479_),
    .B2(_04173_),
    .C1(_04107_),
    .C2(_04220_),
    .ZN(_04649_));
 OR2_X1 _26997_ (.A1(_04647_),
    .A2(_04649_),
    .ZN(_04650_));
 NOR2_X1 _26998_ (.A1(_04074_),
    .A2(_04107_),
    .ZN(_04651_));
 MUX2_X1 _26999_ (.A(_04417_),
    .B(_04651_),
    .S(_04046_),
    .Z(_04652_));
 AOI22_X2 _27000_ (.A1(_04070_),
    .A2(_04246_),
    .B1(_04169_),
    .B2(_04244_),
    .ZN(_04653_));
 OAI22_X2 _27001_ (.A1(_04061_),
    .A2(_04125_),
    .B1(_04653_),
    .B2(_04047_),
    .ZN(_04654_));
 AOI221_X2 _27002_ (.A(_04650_),
    .B1(_04652_),
    .B2(_04071_),
    .C1(_04143_),
    .C2(_04654_),
    .ZN(_04655_));
 AND3_X1 _27003_ (.A1(_04037_),
    .A2(_04088_),
    .A3(_04655_),
    .ZN(_04656_));
 NAND4_X4 _27004_ (.A1(_04628_),
    .A2(_04638_),
    .A3(_04646_),
    .A4(_04656_),
    .ZN(_04657_));
 AND2_X1 _27005_ (.A1(_00196_),
    .A2(_17013_),
    .ZN(_04658_));
 NAND3_X1 _27006_ (.A1(\core.keymem.key_mem[3][122] ),
    .A2(_17048_),
    .A3(_16970_),
    .ZN(_04659_));
 OAI211_X2 _27007_ (.A(\core.keymem.key_mem[8][122] ),
    .B(_17527_),
    .C1(_17128_),
    .C2(_17129_),
    .ZN(_04660_));
 OAI211_X2 _27008_ (.A(\core.keymem.key_mem[10][122] ),
    .B(_17016_),
    .C1(_17128_),
    .C2(_17129_),
    .ZN(_04661_));
 OAI211_X2 _27009_ (.A(\core.keymem.key_mem[7][122] ),
    .B(_17048_),
    .C1(_17114_),
    .C2(_17115_),
    .ZN(_04662_));
 NAND4_X2 _27010_ (.A1(_04659_),
    .A2(_04660_),
    .A3(_04661_),
    .A4(_04662_),
    .ZN(_04663_));
 NAND3_X1 _27011_ (.A1(\core.keymem.key_mem[14][122] ),
    .A2(_16882_),
    .A3(_17156_),
    .ZN(_04664_));
 NAND3_X1 _27012_ (.A1(\core.keymem.key_mem[2][122] ),
    .A2(_17120_),
    .A3(_17156_),
    .ZN(_04665_));
 OAI211_X2 _27013_ (.A(\core.keymem.key_mem[11][122] ),
    .B(_17111_),
    .C1(_16886_),
    .C2(_16890_),
    .ZN(_04666_));
 OAI211_X2 _27014_ (.A(\core.keymem.key_mem[6][122] ),
    .B(_17156_),
    .C1(_17622_),
    .C2(_17146_),
    .ZN(_04667_));
 NAND4_X2 _27015_ (.A1(_04664_),
    .A2(_04665_),
    .A3(_04666_),
    .A4(_04667_),
    .ZN(_04668_));
 OAI211_X2 _27016_ (.A(\core.keymem.key_mem[13][122] ),
    .B(_17024_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_04669_));
 OAI221_X2 _27017_ (.A(\core.keymem.key_mem[9][122] ),
    .B1(_16927_),
    .B2(_16929_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_04670_));
 OAI211_X2 _27018_ (.A(\core.keymem.key_mem[1][122] ),
    .B(_17827_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_04671_));
 OAI211_X2 _27019_ (.A(\core.keymem.key_mem[4][122] ),
    .B(_17028_),
    .C1(_17030_),
    .C2(_17031_),
    .ZN(_04672_));
 NAND4_X2 _27020_ (.A1(_04669_),
    .A2(_04670_),
    .A3(_04671_),
    .A4(_04672_),
    .ZN(_04673_));
 INV_X1 _27021_ (.A(\core.keymem.key_mem[12][122] ),
    .ZN(_04674_));
 INV_X1 _27022_ (.A(\core.keymem.key_mem[5][122] ),
    .ZN(_04675_));
 OAI22_X2 _27023_ (.A1(_04674_),
    .A2(_17843_),
    .B1(_03591_),
    .B2(_04675_),
    .ZN(_04676_));
 NOR4_X4 _27024_ (.A1(_04663_),
    .A2(_04668_),
    .A3(_04673_),
    .A4(_04676_),
    .ZN(_04677_));
 AOI21_X4 _27025_ (.A(_04658_),
    .B1(_04677_),
    .B2(_17533_),
    .ZN(_04678_));
 XNOR2_X2 _27026_ (.A(\core.dec_block.block_w0_reg[26] ),
    .B(_04678_),
    .ZN(_04679_));
 XNOR2_X1 _27027_ (.A(\block_reg[0][26] ),
    .B(_04678_),
    .ZN(_04680_));
 OAI22_X1 _27028_ (.A1(_16555_),
    .A2(_04679_),
    .B1(_04680_),
    .B2(_18552_),
    .ZN(_04681_));
 NOR2_X1 _27029_ (.A1(_04657_),
    .A2(_04681_),
    .ZN(_04682_));
 XNOR2_X2 _27030_ (.A(_03915_),
    .B(_03976_),
    .ZN(_04683_));
 XNOR2_X2 _27031_ (.A(_19385_),
    .B(_04683_),
    .ZN(_04684_));
 AND2_X1 _27032_ (.A1(_00200_),
    .A2(_16873_),
    .ZN(_04685_));
 AOI22_X1 _27033_ (.A1(\core.keymem.key_mem[11][98] ),
    .A2(_16507_),
    .B1(_17178_),
    .B2(\core.keymem.key_mem[1][98] ),
    .ZN(_04686_));
 AOI22_X2 _27034_ (.A1(\core.keymem.key_mem[8][98] ),
    .A2(_16530_),
    .B1(_16537_),
    .B2(\core.keymem.key_mem[9][98] ),
    .ZN(_04687_));
 AOI22_X2 _27035_ (.A1(\core.keymem.key_mem[4][98] ),
    .A2(_16458_),
    .B1(_16408_),
    .B2(\core.keymem.key_mem[7][98] ),
    .ZN(_04688_));
 AOI21_X1 _27036_ (.A(_16983_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][98] ),
    .ZN(_04689_));
 NAND4_X2 _27037_ (.A1(_04686_),
    .A2(_04687_),
    .A3(_04688_),
    .A4(_04689_),
    .ZN(_04690_));
 MUX2_X1 _27038_ (.A(\core.keymem.key_mem[6][98] ),
    .B(\core.keymem.key_mem[14][98] ),
    .S(_17055_),
    .Z(_04691_));
 AOI22_X2 _27039_ (.A1(\core.keymem.key_mem[2][98] ),
    .A2(_17121_),
    .B1(_17051_),
    .B2(_04691_),
    .ZN(_04692_));
 NOR2_X2 _27040_ (.A1(_16968_),
    .A2(_04692_),
    .ZN(_04693_));
 AOI22_X1 _27041_ (.A1(\core.keymem.key_mem[10][98] ),
    .A2(_16516_),
    .B1(_16469_),
    .B2(\core.keymem.key_mem[5][98] ),
    .ZN(_04694_));
 AOI22_X1 _27042_ (.A1(\core.keymem.key_mem[3][98] ),
    .A2(_16387_),
    .B1(_16540_),
    .B2(\core.keymem.key_mem[12][98] ),
    .ZN(_04695_));
 NAND2_X1 _27043_ (.A1(_04694_),
    .A2(_04695_),
    .ZN(_04696_));
 NOR3_X4 _27044_ (.A1(_04690_),
    .A2(_04693_),
    .A3(_04696_),
    .ZN(_04697_));
 NOR2_X4 _27045_ (.A1(_04685_),
    .A2(_04697_),
    .ZN(_04698_));
 XNOR2_X2 _27046_ (.A(\core.dec_block.block_w0_reg[2] ),
    .B(_04698_),
    .ZN(_04699_));
 XNOR2_X2 _27047_ (.A(_04684_),
    .B(_04699_),
    .ZN(_04700_));
 NAND2_X1 _27048_ (.A1(_00185_),
    .A2(_16983_),
    .ZN(_04701_));
 OAI211_X2 _27049_ (.A(\core.keymem.key_mem[11][103] ),
    .B(_17111_),
    .C1(_16886_),
    .C2(_16890_),
    .ZN(_04702_));
 OAI211_X2 _27050_ (.A(\core.keymem.key_mem[4][103] ),
    .B(_17527_),
    .C1(_17146_),
    .C2(_17622_),
    .ZN(_04703_));
 OAI211_X2 _27051_ (.A(\core.keymem.key_mem[1][103] ),
    .B(_17120_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_04704_));
 OAI221_X1 _27052_ (.A(\core.keymem.key_mem[9][103] ),
    .B1(_16927_),
    .B2(_16929_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_04705_));
 AND4_X1 _27053_ (.A1(_04702_),
    .A2(_04703_),
    .A3(_04704_),
    .A4(_04705_),
    .ZN(_04706_));
 OAI211_X2 _27054_ (.A(\core.keymem.key_mem[13][103] ),
    .B(_17024_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_04707_));
 OAI221_X1 _27055_ (.A(\core.keymem.key_mem[5][103] ),
    .B1(_16896_),
    .B2(_16899_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_04708_));
 NAND3_X1 _27056_ (.A1(\core.keymem.key_mem[14][103] ),
    .A2(_17024_),
    .A3(_17026_),
    .ZN(_04709_));
 AND4_X1 _27057_ (.A1(_16486_),
    .A2(_04707_),
    .A3(_04708_),
    .A4(_04709_),
    .ZN(_04710_));
 INV_X1 _27058_ (.A(\core.keymem.key_mem[6][103] ),
    .ZN(_04711_));
 AOI21_X1 _27059_ (.A(_04711_),
    .B1(_16402_),
    .B2(_16404_),
    .ZN(_04712_));
 MUX2_X1 _27060_ (.A(\core.keymem.key_mem[2][103] ),
    .B(\core.keymem.key_mem[10][103] ),
    .S(_16972_),
    .Z(_04713_));
 AND2_X1 _27061_ (.A1(_17043_),
    .A2(_04713_),
    .ZN(_04714_));
 OAI21_X1 _27062_ (.A(_17101_),
    .B1(_04712_),
    .B2(_04714_),
    .ZN(_04715_));
 OAI211_X2 _27063_ (.A(\core.keymem.key_mem[7][103] ),
    .B(_17074_),
    .C1(_17146_),
    .C2(_17031_),
    .ZN(_04716_));
 NAND3_X1 _27064_ (.A1(\core.keymem.key_mem[3][103] ),
    .A2(_17111_),
    .A3(_17120_),
    .ZN(_04717_));
 OAI211_X2 _27065_ (.A(\core.keymem.key_mem[8][103] ),
    .B(_17028_),
    .C1(_17035_),
    .C2(_17036_),
    .ZN(_04718_));
 NAND3_X1 _27066_ (.A1(\core.keymem.key_mem[12][103] ),
    .A2(_17024_),
    .A3(_17028_),
    .ZN(_04719_));
 AND4_X1 _27067_ (.A1(_04716_),
    .A2(_04717_),
    .A3(_04718_),
    .A4(_04719_),
    .ZN(_04720_));
 NAND4_X2 _27068_ (.A1(_04706_),
    .A2(_04710_),
    .A3(_04715_),
    .A4(_04720_),
    .ZN(_04721_));
 AND2_X2 _27069_ (.A1(_04701_),
    .A2(_04721_),
    .ZN(_04722_));
 XNOR2_X2 _27070_ (.A(_16581_),
    .B(_04722_),
    .ZN(_04723_));
 XNOR2_X2 _27071_ (.A(_04589_),
    .B(_04723_),
    .ZN(_04724_));
 XNOR2_X2 _27072_ (.A(_04700_),
    .B(_04724_),
    .ZN(_04725_));
 XOR2_X1 _27073_ (.A(_04263_),
    .B(_04327_),
    .Z(_04726_));
 XNOR2_X1 _27074_ (.A(_04311_),
    .B(_04726_),
    .ZN(_04727_));
 XNOR2_X2 _27075_ (.A(_04725_),
    .B(_04727_),
    .ZN(_04728_));
 XNOR2_X2 _27076_ (.A(_17740_),
    .B(_18478_),
    .ZN(_04729_));
 XOR2_X1 _27077_ (.A(_19192_),
    .B(_04552_),
    .Z(_04730_));
 XNOR2_X1 _27078_ (.A(_04729_),
    .B(_04730_),
    .ZN(_04731_));
 XNOR2_X2 _27079_ (.A(_04728_),
    .B(_04731_),
    .ZN(_04732_));
 OAI21_X1 _27080_ (.A(_04682_),
    .B1(_04732_),
    .B2(_17204_),
    .ZN(_04733_));
 MUX2_X1 _27081_ (.A(\core.dec_block.block_w0_reg[26] ),
    .B(_04733_),
    .S(_16365_),
    .Z(_00585_));
 NOR2_X2 _27082_ (.A1(_04029_),
    .A2(_04130_),
    .ZN(_04734_));
 NOR2_X1 _27083_ (.A1(_04042_),
    .A2(_04045_),
    .ZN(_04735_));
 OAI21_X1 _27084_ (.A(_04734_),
    .B1(_04162_),
    .B2(_04735_),
    .ZN(_04736_));
 OAI221_X2 _27085_ (.A(_04736_),
    .B1(_04414_),
    .B2(_04409_),
    .C1(_04389_),
    .C2(_04408_),
    .ZN(_04737_));
 OAI21_X1 _27086_ (.A(_04148_),
    .B1(_04112_),
    .B2(_04107_),
    .ZN(_04738_));
 AOI21_X1 _27087_ (.A(_04737_),
    .B1(_04738_),
    .B2(_04179_),
    .ZN(_04739_));
 OAI221_X1 _27088_ (.A(_04068_),
    .B1(_04060_),
    .B2(_04193_),
    .C1(_04381_),
    .C2(_04142_),
    .ZN(_04740_));
 AOI21_X1 _27089_ (.A(_04482_),
    .B1(_04223_),
    .B2(_04095_),
    .ZN(_04741_));
 OAI21_X1 _27090_ (.A(_04740_),
    .B1(_04741_),
    .B2(_04451_),
    .ZN(_04742_));
 NAND2_X1 _27091_ (.A1(_04739_),
    .A2(_04742_),
    .ZN(_04743_));
 MUX2_X1 _27092_ (.A(_04025_),
    .B(_04200_),
    .S(_04059_),
    .Z(_04744_));
 NAND3_X1 _27093_ (.A1(_04500_),
    .A2(_04150_),
    .A3(_04744_),
    .ZN(_04745_));
 OAI221_X2 _27094_ (.A(_04745_),
    .B1(_04223_),
    .B2(_04415_),
    .C1(_04193_),
    .C2(_04511_),
    .ZN(_04746_));
 NAND2_X1 _27095_ (.A1(_04046_),
    .A2(_04200_),
    .ZN(_04747_));
 NOR3_X1 _27096_ (.A1(_04071_),
    .A2(_04452_),
    .A3(_04747_),
    .ZN(_04748_));
 OAI221_X2 _27097_ (.A(_04636_),
    .B1(_04187_),
    .B2(_04169_),
    .C1(_04192_),
    .C2(_04494_),
    .ZN(_04749_));
 NOR4_X2 _27098_ (.A1(_04743_),
    .A2(_04746_),
    .A3(_04748_),
    .A4(_04749_),
    .ZN(_04750_));
 NOR2_X1 _27099_ (.A1(_04094_),
    .A2(_04136_),
    .ZN(_04751_));
 NOR3_X1 _27100_ (.A1(_04001_),
    .A2(_04164_),
    .A3(_04751_),
    .ZN(_04752_));
 NOR2_X1 _27101_ (.A1(_04030_),
    .A2(_04409_),
    .ZN(_04753_));
 AOI21_X1 _27102_ (.A(_04752_),
    .B1(_04753_),
    .B2(_04101_),
    .ZN(_04754_));
 NOR3_X1 _27103_ (.A1(_04074_),
    .A2(_04001_),
    .A3(_04104_),
    .ZN(_04755_));
 AOI21_X1 _27104_ (.A(_04755_),
    .B1(_04137_),
    .B2(_04074_),
    .ZN(_04756_));
 OAI22_X2 _27105_ (.A1(_04142_),
    .A2(_04754_),
    .B1(_04756_),
    .B2(_04059_),
    .ZN(_04757_));
 NOR2_X1 _27106_ (.A1(_04045_),
    .A2(_04111_),
    .ZN(_04758_));
 AOI22_X1 _27107_ (.A1(_04156_),
    .A2(_04172_),
    .B1(_04758_),
    .B2(_04110_),
    .ZN(_04759_));
 OAI21_X1 _27108_ (.A(_04759_),
    .B1(_04412_),
    .B2(_04077_),
    .ZN(_04760_));
 AOI221_X2 _27109_ (.A(_04757_),
    .B1(_04760_),
    .B2(_04229_),
    .C1(_04091_),
    .C2(_04096_),
    .ZN(_04761_));
 NOR3_X1 _27110_ (.A1(_04197_),
    .A2(_04441_),
    .A3(_04237_),
    .ZN(_04762_));
 OAI21_X1 _27111_ (.A(_04600_),
    .B1(_04237_),
    .B2(_04500_),
    .ZN(_04763_));
 AND3_X1 _27112_ (.A1(_04072_),
    .A2(_04451_),
    .A3(_04763_),
    .ZN(_04764_));
 OAI21_X1 _27113_ (.A(_04501_),
    .B1(_04762_),
    .B2(_04764_),
    .ZN(_04765_));
 AND4_X1 _27114_ (.A1(_04232_),
    .A2(_04750_),
    .A3(_04761_),
    .A4(_04765_),
    .ZN(_04766_));
 NAND3_X1 _27115_ (.A1(_04229_),
    .A2(_04462_),
    .A3(_04179_),
    .ZN(_04767_));
 MUX2_X1 _27116_ (.A(_04130_),
    .B(_04174_),
    .S(_04059_),
    .Z(_04768_));
 OAI221_X1 _27117_ (.A(_04767_),
    .B1(_04127_),
    .B2(_04071_),
    .C1(_04143_),
    .C2(_04768_),
    .ZN(_04769_));
 AOI21_X1 _27118_ (.A(_04417_),
    .B1(_04034_),
    .B2(_04142_),
    .ZN(_04770_));
 OAI22_X1 _27119_ (.A1(_04043_),
    .A2(_04061_),
    .B1(_04169_),
    .B2(_04770_),
    .ZN(_04771_));
 NOR3_X1 _27120_ (.A1(_04470_),
    .A2(_04769_),
    .A3(_04771_),
    .ZN(_04772_));
 MUX2_X1 _27121_ (.A(_04478_),
    .B(_04518_),
    .S(_04115_),
    .Z(_04773_));
 OAI21_X1 _27122_ (.A(_04115_),
    .B1(_04048_),
    .B2(_04192_),
    .ZN(_04774_));
 OAI21_X1 _27123_ (.A(_04774_),
    .B1(_04034_),
    .B2(_04115_),
    .ZN(_04775_));
 MUX2_X1 _27124_ (.A(_04773_),
    .B(_04775_),
    .S(_04500_),
    .Z(_04776_));
 AOI21_X2 _27125_ (.A(_04772_),
    .B1(_04776_),
    .B2(_04470_),
    .ZN(_04777_));
 AOI21_X1 _27126_ (.A(_04166_),
    .B1(_04221_),
    .B2(_04246_),
    .ZN(_04778_));
 AOI21_X1 _27127_ (.A(_04157_),
    .B1(_04460_),
    .B2(_04034_),
    .ZN(_04779_));
 NOR2_X1 _27128_ (.A1(_04161_),
    .A2(_04460_),
    .ZN(_04780_));
 NAND2_X2 _27129_ (.A1(_04091_),
    .A2(_04188_),
    .ZN(_04781_));
 OAI222_X2 _27130_ (.A1(_04043_),
    .A2(_04778_),
    .B1(_04779_),
    .B2(_04780_),
    .C1(_04781_),
    .C2(_04478_),
    .ZN(_04782_));
 NAND2_X1 _27131_ (.A1(_03995_),
    .A2(_04083_),
    .ZN(_04783_));
 AOI21_X1 _27132_ (.A(_04452_),
    .B1(_04061_),
    .B2(_04783_),
    .ZN(_04784_));
 AOI21_X1 _27133_ (.A(_04784_),
    .B1(_04188_),
    .B2(_04083_),
    .ZN(_04785_));
 NOR2_X1 _27134_ (.A1(_04043_),
    .A2(_04785_),
    .ZN(_04786_));
 NOR3_X1 _27135_ (.A1(_04043_),
    .A2(_04047_),
    .A3(_04174_),
    .ZN(_04787_));
 NOR3_X1 _27136_ (.A1(_04086_),
    .A2(_04111_),
    .A3(_04381_),
    .ZN(_04788_));
 OAI21_X1 _27137_ (.A(_04614_),
    .B1(_04787_),
    .B2(_04788_),
    .ZN(_04789_));
 OAI221_X2 _27138_ (.A(_04789_),
    .B1(_04511_),
    .B2(_04127_),
    .C1(_04409_),
    .C2(_04781_),
    .ZN(_04790_));
 NOR4_X4 _27139_ (.A1(_04777_),
    .A2(_04782_),
    .A3(_04786_),
    .A4(_04790_),
    .ZN(_04791_));
 NAND4_X4 _27140_ (.A1(_04504_),
    .A2(_04655_),
    .A3(_04766_),
    .A4(_04791_),
    .ZN(_04792_));
 AOI222_X2 _27141_ (.A1(\core.keymem.key_mem[4][123] ),
    .A2(_17713_),
    .B1(_16386_),
    .B2(\core.keymem.key_mem[3][123] ),
    .C1(_16515_),
    .C2(\core.keymem.key_mem[10][123] ),
    .ZN(_04793_));
 AOI22_X1 _27142_ (.A1(\core.keymem.key_mem[14][123] ),
    .A2(_16999_),
    .B1(_17768_),
    .B2(\core.keymem.key_mem[11][123] ),
    .ZN(_04794_));
 AOI22_X1 _27143_ (.A1(\core.keymem.key_mem[1][123] ),
    .A2(_16417_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][123] ),
    .ZN(_04795_));
 NAND3_X1 _27144_ (.A1(_04793_),
    .A2(_04794_),
    .A3(_04795_),
    .ZN(_04796_));
 AOI22_X1 _27145_ (.A1(\core.keymem.key_mem[7][123] ),
    .A2(_17789_),
    .B1(_17786_),
    .B2(\core.keymem.key_mem[2][123] ),
    .ZN(_04797_));
 AOI22_X1 _27146_ (.A1(\core.keymem.key_mem[12][123] ),
    .A2(_17720_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][123] ),
    .ZN(_04798_));
 AOI22_X1 _27147_ (.A1(\core.keymem.key_mem[8][123] ),
    .A2(_17666_),
    .B1(_17668_),
    .B2(\core.keymem.key_mem[9][123] ),
    .ZN(_04799_));
 AOI21_X1 _27148_ (.A(_16495_),
    .B1(_16521_),
    .B2(\core.keymem.key_mem[6][123] ),
    .ZN(_04800_));
 NAND4_X1 _27149_ (.A1(_04797_),
    .A2(_04798_),
    .A3(_04799_),
    .A4(_04800_),
    .ZN(_04801_));
 NOR2_X1 _27150_ (.A1(_04796_),
    .A2(_04801_),
    .ZN(_04802_));
 AOI21_X4 _27151_ (.A(_04802_),
    .B1(_16873_),
    .B2(_00202_),
    .ZN(_04803_));
 XNOR2_X2 _27152_ (.A(\core.dec_block.block_w0_reg[27] ),
    .B(_04803_),
    .ZN(_04804_));
 XNOR2_X1 _27153_ (.A(\block_reg[0][27] ),
    .B(_04803_),
    .ZN(_04805_));
 OAI22_X1 _27154_ (.A1(_19180_),
    .A2(_04804_),
    .B1(_04805_),
    .B2(_18552_),
    .ZN(_04806_));
 XOR2_X2 _27155_ (.A(_03287_),
    .B(_04316_),
    .Z(_04807_));
 XOR2_X1 _27156_ (.A(_16551_),
    .B(_04807_),
    .Z(_04808_));
 XOR2_X2 _27157_ (.A(_18478_),
    .B(_04564_),
    .Z(_04809_));
 XNOR2_X1 _27158_ (.A(_04312_),
    .B(_04809_),
    .ZN(_04810_));
 XNOR2_X2 _27159_ (.A(_04552_),
    .B(_04810_),
    .ZN(_04811_));
 XNOR2_X2 _27160_ (.A(_18410_),
    .B(_04327_),
    .ZN(_04812_));
 XNOR2_X2 _27161_ (.A(_04365_),
    .B(_04723_),
    .ZN(_04813_));
 XNOR2_X1 _27162_ (.A(_04812_),
    .B(_04813_),
    .ZN(_04814_));
 XNOR2_X1 _27163_ (.A(_04263_),
    .B(_04349_),
    .ZN(_04815_));
 XNOR2_X2 _27164_ (.A(_04814_),
    .B(_04815_),
    .ZN(_04816_));
 XNOR2_X1 _27165_ (.A(_04811_),
    .B(_04816_),
    .ZN(_04817_));
 XNOR2_X1 _27166_ (.A(_04808_),
    .B(_04817_),
    .ZN(_04818_));
 XNOR2_X2 _27167_ (.A(_18064_),
    .B(_18550_),
    .ZN(_04819_));
 XNOR2_X2 _27168_ (.A(_04349_),
    .B(_04679_),
    .ZN(_04820_));
 XNOR2_X1 _27169_ (.A(_04819_),
    .B(_04820_),
    .ZN(_04821_));
 AOI222_X2 _27170_ (.A1(\core.keymem.key_mem[14][99] ),
    .A2(_17719_),
    .B1(_16452_),
    .B2(\core.keymem.key_mem[8][99] ),
    .C1(_16472_),
    .C2(\core.keymem.key_mem[13][99] ),
    .ZN(_04822_));
 AOI22_X1 _27171_ (.A1(\core.keymem.key_mem[3][99] ),
    .A2(_16987_),
    .B1(_16989_),
    .B2(\core.keymem.key_mem[10][99] ),
    .ZN(_04823_));
 AOI22_X1 _27172_ (.A1(\core.keymem.key_mem[2][99] ),
    .A2(_17786_),
    .B1(_17720_),
    .B2(\core.keymem.key_mem[12][99] ),
    .ZN(_04824_));
 NAND3_X1 _27173_ (.A1(_04822_),
    .A2(_04823_),
    .A3(_04824_),
    .ZN(_04825_));
 AOI22_X1 _27174_ (.A1(\core.keymem.key_mem[6][99] ),
    .A2(_17695_),
    .B1(_16506_),
    .B2(\core.keymem.key_mem[11][99] ),
    .ZN(_04826_));
 AOI22_X1 _27175_ (.A1(\core.keymem.key_mem[1][99] ),
    .A2(_16855_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][99] ),
    .ZN(_04827_));
 AOI22_X1 _27176_ (.A1(\core.keymem.key_mem[4][99] ),
    .A2(_17713_),
    .B1(_16512_),
    .B2(\core.keymem.key_mem[7][99] ),
    .ZN(_04828_));
 AOI21_X1 _27177_ (.A(_16495_),
    .B1(_17668_),
    .B2(\core.keymem.key_mem[9][99] ),
    .ZN(_04829_));
 NAND4_X1 _27178_ (.A1(_04826_),
    .A2(_04827_),
    .A3(_04828_),
    .A4(_04829_),
    .ZN(_04830_));
 NOR2_X2 _27179_ (.A1(_04825_),
    .A2(_04830_),
    .ZN(_04831_));
 AOI21_X4 _27180_ (.A(_04831_),
    .B1(_17183_),
    .B2(_00205_),
    .ZN(_04832_));
 XNOR2_X2 _27181_ (.A(\core.dec_block.block_w0_reg[3] ),
    .B(_04832_),
    .ZN(_04833_));
 XNOR2_X1 _27182_ (.A(_19385_),
    .B(_04833_),
    .ZN(_04834_));
 XNOR2_X1 _27183_ (.A(_03976_),
    .B(_04834_),
    .ZN(_04835_));
 XNOR2_X1 _27184_ (.A(_04821_),
    .B(_04835_),
    .ZN(_04836_));
 XNOR2_X1 _27185_ (.A(_04818_),
    .B(_04836_),
    .ZN(_04837_));
 NOR2_X1 _27186_ (.A1(_17203_),
    .A2(_04837_),
    .ZN(_04838_));
 NOR4_X1 _27187_ (.A1(_17744_),
    .A2(_04792_),
    .A3(_04806_),
    .A4(_04838_),
    .ZN(_04839_));
 INV_X1 _27188_ (.A(\core.dec_block.block_w0_reg[27] ),
    .ZN(_04840_));
 AOI21_X1 _27189_ (.A(_04839_),
    .B1(_17744_),
    .B2(_04840_),
    .ZN(_00586_));
 OAI21_X1 _27190_ (.A(_04516_),
    .B1(_04488_),
    .B2(_04466_),
    .ZN(_04841_));
 AOI21_X1 _27191_ (.A(_04115_),
    .B1(_04086_),
    .B2(_04084_),
    .ZN(_04842_));
 OAI21_X1 _27192_ (.A(_04083_),
    .B1(_04735_),
    .B2(_04842_),
    .ZN(_04843_));
 NOR3_X1 _27193_ (.A1(_04244_),
    .A2(_04137_),
    .A3(_04156_),
    .ZN(_04844_));
 OAI21_X1 _27194_ (.A(_04843_),
    .B1(_04844_),
    .B2(_04494_),
    .ZN(_04845_));
 NAND4_X1 _27195_ (.A1(_04071_),
    .A2(_04132_),
    .A3(_04614_),
    .A4(_04110_),
    .ZN(_04846_));
 MUX2_X1 _27196_ (.A(_04409_),
    .B(_04237_),
    .S(_04070_),
    .Z(_04847_));
 OAI221_X2 _27197_ (.A(_04846_),
    .B1(_04237_),
    .B2(_04614_),
    .C1(_04132_),
    .C2(_04847_),
    .ZN(_04848_));
 AOI221_X2 _27198_ (.A(_04841_),
    .B1(_04845_),
    .B2(_04501_),
    .C1(_04467_),
    .C2(_04848_),
    .ZN(_04849_));
 MUX2_X1 _27199_ (.A(_04409_),
    .B(_04167_),
    .S(_04614_),
    .Z(_04850_));
 OAI21_X1 _27200_ (.A(_04614_),
    .B1(_04110_),
    .B2(_04461_),
    .ZN(_04851_));
 AOI21_X1 _27201_ (.A(_04197_),
    .B1(_04095_),
    .B2(_04851_),
    .ZN(_04852_));
 AOI21_X1 _27202_ (.A(_04132_),
    .B1(_04389_),
    .B2(_04176_),
    .ZN(_04853_));
 NOR2_X1 _27203_ (.A1(_04852_),
    .A2(_04853_),
    .ZN(_04854_));
 OAI221_X1 _27204_ (.A(_04466_),
    .B1(_04470_),
    .B2(_04850_),
    .C1(_04854_),
    .C2(_04467_),
    .ZN(_04855_));
 NAND2_X1 _27205_ (.A1(_04143_),
    .A2(_04139_),
    .ZN(_04856_));
 OAI21_X1 _27206_ (.A(_04856_),
    .B1(_04409_),
    .B2(_04143_),
    .ZN(_04857_));
 NAND2_X1 _27207_ (.A1(_04197_),
    .A2(_04857_),
    .ZN(_04858_));
 OAI21_X1 _27208_ (.A(_04130_),
    .B1(_04237_),
    .B2(_04181_),
    .ZN(_04859_));
 AOI21_X1 _27209_ (.A(_04734_),
    .B1(_04859_),
    .B2(_04470_),
    .ZN(_04860_));
 OAI221_X1 _27210_ (.A(_04858_),
    .B1(_04860_),
    .B2(_04467_),
    .C1(_04501_),
    .C2(_04856_),
    .ZN(_04861_));
 OAI21_X1 _27211_ (.A(_04855_),
    .B1(_04861_),
    .B2(_04466_),
    .ZN(_04862_));
 OAI22_X1 _27212_ (.A1(_04111_),
    .A2(_04129_),
    .B1(_04479_),
    .B2(_04061_),
    .ZN(_04863_));
 NAND3_X1 _27213_ (.A1(_04212_),
    .A2(_04051_),
    .A3(_04863_),
    .ZN(_04864_));
 OAI21_X1 _27214_ (.A(_04381_),
    .B1(_04192_),
    .B2(_04048_),
    .ZN(_04865_));
 NAND3_X1 _27215_ (.A1(_04207_),
    .A2(_04459_),
    .A3(_04865_),
    .ZN(_04866_));
 OAI21_X1 _27216_ (.A(_04083_),
    .B1(_04162_),
    .B2(_04219_),
    .ZN(_04867_));
 NAND3_X1 _27217_ (.A1(_04451_),
    .A2(_04246_),
    .A3(_04091_),
    .ZN(_04868_));
 NAND4_X1 _27218_ (.A1(_04864_),
    .A2(_04866_),
    .A3(_04867_),
    .A4(_04868_),
    .ZN(_04869_));
 AOI21_X1 _27219_ (.A(_04164_),
    .B1(_04165_),
    .B2(_04167_),
    .ZN(_04870_));
 AOI21_X1 _27220_ (.A(_04182_),
    .B1(_04223_),
    .B2(_04747_),
    .ZN(_04871_));
 NOR4_X1 _27221_ (.A1(_04194_),
    .A2(_04869_),
    .A3(_04870_),
    .A4(_04871_),
    .ZN(_04872_));
 AOI22_X1 _27222_ (.A1(_04461_),
    .A2(_04161_),
    .B1(_04758_),
    .B2(_04025_),
    .ZN(_04873_));
 NAND3_X1 _27223_ (.A1(_03989_),
    .A2(_04244_),
    .A3(_04188_),
    .ZN(_04874_));
 OAI21_X1 _27224_ (.A(_04156_),
    .B1(_04463_),
    .B2(_04513_),
    .ZN(_04875_));
 NAND3_X2 _27225_ (.A1(_04873_),
    .A2(_04874_),
    .A3(_04875_),
    .ZN(_04876_));
 NOR3_X1 _27226_ (.A1(_04649_),
    .A2(_04746_),
    .A3(_04876_),
    .ZN(_04877_));
 AOI21_X1 _27227_ (.A(_04482_),
    .B1(_04783_),
    .B2(_04747_),
    .ZN(_04878_));
 AOI21_X1 _27228_ (.A(_04878_),
    .B1(_04651_),
    .B2(_04150_),
    .ZN(_04879_));
 MUX2_X1 _27229_ (.A(_04107_),
    .B(_04126_),
    .S(_04041_),
    .Z(_04880_));
 MUX2_X1 _27230_ (.A(_04381_),
    .B(_04880_),
    .S(_04084_),
    .Z(_04881_));
 AOI21_X1 _27231_ (.A(_04025_),
    .B1(_04376_),
    .B2(_04452_),
    .ZN(_04882_));
 OAI221_X2 _27232_ (.A(_04879_),
    .B1(_04881_),
    .B2(_04125_),
    .C1(_04522_),
    .C2(_04882_),
    .ZN(_04883_));
 NOR3_X1 _27233_ (.A1(_04070_),
    .A2(_04002_),
    .A3(_04077_),
    .ZN(_04884_));
 AOI21_X1 _27234_ (.A(_04884_),
    .B1(_04376_),
    .B2(_04070_),
    .ZN(_04885_));
 OAI33_X1 _27235_ (.A1(_04389_),
    .A2(_04146_),
    .A3(_04482_),
    .B1(_04885_),
    .B2(_04500_),
    .B3(_04191_),
    .ZN(_04886_));
 NOR2_X1 _27236_ (.A1(_04057_),
    .A2(_04389_),
    .ZN(_04887_));
 OAI21_X1 _27237_ (.A(_04198_),
    .B1(_04078_),
    .B2(_04887_),
    .ZN(_04888_));
 NAND3_X1 _27238_ (.A1(_04500_),
    .A2(_04071_),
    .A3(_04376_),
    .ZN(_04889_));
 AOI21_X1 _27239_ (.A(_04129_),
    .B1(_04888_),
    .B2(_04889_),
    .ZN(_04890_));
 NOR3_X1 _27240_ (.A1(_04883_),
    .A2(_04886_),
    .A3(_04890_),
    .ZN(_04891_));
 OAI21_X1 _27241_ (.A(_04029_),
    .B1(_04094_),
    .B2(_04137_),
    .ZN(_04892_));
 AOI21_X1 _27242_ (.A(_04160_),
    .B1(_04630_),
    .B2(_04892_),
    .ZN(_04893_));
 AOI21_X1 _27243_ (.A(_04169_),
    .B1(_04201_),
    .B2(_04223_),
    .ZN(_04894_));
 OR2_X1 _27244_ (.A1(_04893_),
    .A2(_04894_),
    .ZN(_04895_));
 AOI21_X1 _27245_ (.A(_04030_),
    .B1(_04381_),
    .B2(_04174_),
    .ZN(_04896_));
 OAI21_X1 _27246_ (.A(_04047_),
    .B1(_04133_),
    .B2(_04896_),
    .ZN(_04897_));
 OAI21_X1 _27247_ (.A(_04897_),
    .B1(_04641_),
    .B2(_04068_),
    .ZN(_04898_));
 AOI221_X2 _27248_ (.A(_04642_),
    .B1(_04895_),
    .B2(_04191_),
    .C1(_04898_),
    .C2(_03989_),
    .ZN(_04899_));
 AND4_X1 _27249_ (.A1(_04872_),
    .A2(_04877_),
    .A3(_04891_),
    .A4(_04899_),
    .ZN(_04900_));
 NAND4_X2 _27250_ (.A1(_04450_),
    .A2(_04849_),
    .A3(_04862_),
    .A4(_04900_),
    .ZN(_04901_));
 NAND2_X4 _27251_ (.A1(_18416_),
    .A2(_04901_),
    .ZN(_04902_));
 NAND2_X1 _27252_ (.A1(_00207_),
    .A2(_17578_),
    .ZN(_04903_));
 AOI222_X2 _27253_ (.A1(\core.keymem.key_mem[3][124] ),
    .A2(_17091_),
    .B1(_16537_),
    .B2(\core.keymem.key_mem[9][124] ),
    .C1(\core.keymem.key_mem[12][124] ),
    .C2(_16540_),
    .ZN(_04904_));
 AOI22_X2 _27254_ (.A1(\core.keymem.key_mem[11][124] ),
    .A2(_17769_),
    .B1(_16510_),
    .B2(\core.keymem.key_mem[5][124] ),
    .ZN(_04905_));
 AOI22_X2 _27255_ (.A1(\core.keymem.key_mem[2][124] ),
    .A2(_17086_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][124] ),
    .ZN(_04906_));
 NAND3_X2 _27256_ (.A1(_04904_),
    .A2(_04905_),
    .A3(_04906_),
    .ZN(_04907_));
 AOI22_X2 _27257_ (.A1(\core.keymem.key_mem[4][124] ),
    .A2(_16501_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][124] ),
    .ZN(_04908_));
 AOI21_X1 _27258_ (.A(_16547_),
    .B1(_17085_),
    .B2(\core.keymem.key_mem[7][124] ),
    .ZN(_04909_));
 AOI22_X2 _27259_ (.A1(\core.keymem.key_mem[14][124] ),
    .A2(_17581_),
    .B1(_16522_),
    .B2(\core.keymem.key_mem[6][124] ),
    .ZN(_04910_));
 AOI22_X2 _27260_ (.A1(\core.keymem.key_mem[8][124] ),
    .A2(_17765_),
    .B1(_17082_),
    .B2(\core.keymem.key_mem[10][124] ),
    .ZN(_04911_));
 NAND4_X2 _27261_ (.A1(_04908_),
    .A2(_04909_),
    .A3(_04910_),
    .A4(_04911_),
    .ZN(_04912_));
 OAI21_X4 _27262_ (.A(_04903_),
    .B1(_04907_),
    .B2(_04912_),
    .ZN(_04913_));
 XOR2_X2 _27263_ (.A(\core.dec_block.block_w0_reg[28] ),
    .B(_04913_),
    .Z(_04914_));
 XOR2_X1 _27264_ (.A(\block_reg[0][28] ),
    .B(_04913_),
    .Z(_04915_));
 OAI22_X1 _27265_ (.A1(_19180_),
    .A2(_04914_),
    .B1(_04915_),
    .B2(_18552_),
    .ZN(_04916_));
 INV_X1 _27266_ (.A(_04916_),
    .ZN(_04917_));
 XOR2_X2 _27267_ (.A(_04593_),
    .B(_04811_),
    .Z(_04918_));
 XNOR2_X2 _27268_ (.A(_18326_),
    .B(_18410_),
    .ZN(_04919_));
 XNOR2_X1 _27269_ (.A(_03857_),
    .B(_04919_),
    .ZN(_04920_));
 XNOR2_X1 _27270_ (.A(_04918_),
    .B(_04920_),
    .ZN(_04921_));
 XNOR2_X1 _27271_ (.A(_17740_),
    .B(_18550_),
    .ZN(_04922_));
 XNOR2_X2 _27272_ (.A(_04820_),
    .B(_04922_),
    .ZN(_04923_));
 XOR2_X2 _27273_ (.A(_04311_),
    .B(_04923_),
    .Z(_04924_));
 INV_X1 _27274_ (.A(\core.dec_block.block_w0_reg[4] ),
    .ZN(_04925_));
 AOI22_X1 _27275_ (.A1(\core.keymem.key_mem[2][100] ),
    .A2(_16860_),
    .B1(_16855_),
    .B2(\core.keymem.key_mem[1][100] ),
    .ZN(_04926_));
 AOI22_X1 _27276_ (.A1(\core.keymem.key_mem[3][100] ),
    .A2(_16866_),
    .B1(_16515_),
    .B2(\core.keymem.key_mem[10][100] ),
    .ZN(_04927_));
 AOI22_X1 _27277_ (.A1(\core.keymem.key_mem[9][100] ),
    .A2(_16536_),
    .B1(_16539_),
    .B2(\core.keymem.key_mem[12][100] ),
    .ZN(_04928_));
 AOI22_X1 _27278_ (.A1(\core.keymem.key_mem[4][100] ),
    .A2(_16457_),
    .B1(_16468_),
    .B2(\core.keymem.key_mem[5][100] ),
    .ZN(_04929_));
 NAND4_X1 _27279_ (.A1(_04926_),
    .A2(_04927_),
    .A3(_04928_),
    .A4(_04929_),
    .ZN(_04930_));
 AOI22_X1 _27280_ (.A1(\core.keymem.key_mem[6][100] ),
    .A2(_17695_),
    .B1(_16532_),
    .B2(\core.keymem.key_mem[13][100] ),
    .ZN(_04931_));
 AOI22_X1 _27281_ (.A1(\core.keymem.key_mem[14][100] ),
    .A2(_17719_),
    .B1(_16512_),
    .B2(\core.keymem.key_mem[7][100] ),
    .ZN(_04932_));
 AOI22_X1 _27282_ (.A1(\core.keymem.key_mem[8][100] ),
    .A2(_16529_),
    .B1(_16506_),
    .B2(\core.keymem.key_mem[11][100] ),
    .ZN(_04933_));
 NAND3_X1 _27283_ (.A1(_04931_),
    .A2(_04932_),
    .A3(_04933_),
    .ZN(_04934_));
 NOR2_X1 _27284_ (.A1(_04930_),
    .A2(_04934_),
    .ZN(_04935_));
 MUX2_X2 _27285_ (.A(_00210_),
    .B(_04935_),
    .S(_17533_),
    .Z(_04936_));
 XNOR2_X2 _27286_ (.A(_04925_),
    .B(_04936_),
    .ZN(_04937_));
 XOR2_X1 _27287_ (.A(_18478_),
    .B(_04937_),
    .Z(_04938_));
 XNOR2_X1 _27288_ (.A(_04591_),
    .B(_04938_),
    .ZN(_04939_));
 XNOR2_X2 _27289_ (.A(_04924_),
    .B(_04939_),
    .ZN(_04940_));
 XNOR2_X2 _27290_ (.A(_04349_),
    .B(_04804_),
    .ZN(_04941_));
 XNOR2_X2 _27291_ (.A(_03287_),
    .B(_03976_),
    .ZN(_04942_));
 XNOR2_X2 _27292_ (.A(_03724_),
    .B(_04942_),
    .ZN(_04943_));
 XNOR2_X1 _27293_ (.A(_04941_),
    .B(_04943_),
    .ZN(_04944_));
 XNOR2_X1 _27294_ (.A(_04940_),
    .B(_04944_),
    .ZN(_04945_));
 XNOR2_X1 _27295_ (.A(_04921_),
    .B(_04945_),
    .ZN(_04946_));
 NAND2_X1 _27296_ (.A1(_17748_),
    .A2(_04946_),
    .ZN(_04947_));
 NAND3_X1 _27297_ (.A1(_04902_),
    .A2(_04917_),
    .A3(_04947_),
    .ZN(_04948_));
 MUX2_X1 _27298_ (.A(\core.dec_block.block_w0_reg[28] ),
    .B(_04948_),
    .S(_16365_),
    .Z(_00587_));
 OAI22_X1 _27299_ (.A1(_04130_),
    .A2(_04494_),
    .B1(_04482_),
    .B2(_04223_),
    .ZN(_04949_));
 NAND2_X1 _27300_ (.A1(_04501_),
    .A2(_04949_),
    .ZN(_04950_));
 NAND2_X1 _27301_ (.A1(_04466_),
    .A2(_04887_),
    .ZN(_04951_));
 OAI21_X1 _27302_ (.A(_04951_),
    .B1(_04130_),
    .B2(_04182_),
    .ZN(_04952_));
 AOI21_X1 _27303_ (.A(_04637_),
    .B1(_04952_),
    .B2(_04470_),
    .ZN(_04953_));
 OAI21_X1 _27304_ (.A(_04950_),
    .B1(_04953_),
    .B2(_04501_),
    .ZN(_04954_));
 NOR3_X1 _27305_ (.A1(_04072_),
    .A2(_04501_),
    .A3(_04201_),
    .ZN(_04955_));
 NOR3_X1 _27306_ (.A1(_04142_),
    .A2(_04129_),
    .A3(_04174_),
    .ZN(_04956_));
 NAND2_X1 _27307_ (.A1(_04013_),
    .A2(_04117_),
    .ZN(_04957_));
 NOR4_X1 _27308_ (.A1(_04074_),
    .A2(_03994_),
    .A3(_04050_),
    .A4(_04957_),
    .ZN(_04958_));
 OAI21_X1 _27309_ (.A(_04008_),
    .B1(_04401_),
    .B2(_04958_),
    .ZN(_04959_));
 NOR3_X1 _27310_ (.A1(_04058_),
    .A2(_04212_),
    .A3(_04019_),
    .ZN(_04960_));
 OAI21_X1 _27311_ (.A(_04423_),
    .B1(_04212_),
    .B2(_04058_),
    .ZN(_04961_));
 AOI21_X1 _27312_ (.A(_04960_),
    .B1(_04961_),
    .B2(_04047_),
    .ZN(_04962_));
 OAI21_X1 _27313_ (.A(_04959_),
    .B1(_04962_),
    .B2(_04434_),
    .ZN(_04963_));
 AOI221_X2 _27314_ (.A(_04956_),
    .B1(_04963_),
    .B2(_04452_),
    .C1(_04143_),
    .C2(_04461_),
    .ZN(_04964_));
 NOR2_X1 _27315_ (.A1(_04466_),
    .A2(_04964_),
    .ZN(_04965_));
 NOR3_X2 _27316_ (.A1(_04954_),
    .A2(_04955_),
    .A3(_04965_),
    .ZN(_04966_));
 NOR3_X1 _27317_ (.A1(_04084_),
    .A2(_04127_),
    .A3(_04129_),
    .ZN(_04967_));
 OAI21_X1 _27318_ (.A(_04513_),
    .B1(_04157_),
    .B2(_04186_),
    .ZN(_04968_));
 AOI22_X1 _27319_ (.A1(_04025_),
    .A2(_04091_),
    .B1(_04109_),
    .B2(_04069_),
    .ZN(_04969_));
 OAI221_X1 _27320_ (.A(_04968_),
    .B1(_04518_),
    .B2(_04482_),
    .C1(_03996_),
    .C2(_04969_),
    .ZN(_04970_));
 OR2_X1 _27321_ (.A1(_04967_),
    .A2(_04970_),
    .ZN(_04971_));
 NAND2_X1 _27322_ (.A1(_04244_),
    .A2(_04146_),
    .ZN(_04972_));
 OAI221_X1 _27323_ (.A(_04467_),
    .B1(_04060_),
    .B2(_04381_),
    .C1(_04972_),
    .C2(_04466_),
    .ZN(_04973_));
 OAI221_X1 _27324_ (.A(_04500_),
    .B1(_04198_),
    .B2(_04065_),
    .C1(_04107_),
    .C2(_04164_),
    .ZN(_04974_));
 AOI21_X1 _27325_ (.A(_04971_),
    .B1(_04973_),
    .B2(_04974_),
    .ZN(_04975_));
 AOI21_X1 _27326_ (.A(_04414_),
    .B1(_04223_),
    .B2(_04421_),
    .ZN(_04976_));
 NAND3_X1 _27327_ (.A1(_04115_),
    .A2(_04137_),
    .A3(_04188_),
    .ZN(_04977_));
 NAND3_X1 _27328_ (.A1(_04142_),
    .A2(_04068_),
    .A3(_04462_),
    .ZN(_04978_));
 OAI21_X1 _27329_ (.A(_04977_),
    .B1(_04978_),
    .B2(_04198_),
    .ZN(_04979_));
 NOR4_X2 _27330_ (.A1(_04618_),
    .A2(_04737_),
    .A3(_04976_),
    .A4(_04979_),
    .ZN(_04980_));
 OAI22_X2 _27331_ (.A1(_04415_),
    .A2(_04237_),
    .B1(_04781_),
    .B2(_04061_),
    .ZN(_04981_));
 NOR4_X4 _27332_ (.A1(_04422_),
    .A2(_04485_),
    .A3(_04876_),
    .A4(_04981_),
    .ZN(_04982_));
 NAND4_X2 _27333_ (.A1(_04180_),
    .A2(_04975_),
    .A3(_04980_),
    .A4(_04982_),
    .ZN(_04983_));
 AOI22_X1 _27334_ (.A1(_04198_),
    .A2(_04461_),
    .B1(_04139_),
    .B2(_04101_),
    .ZN(_04984_));
 NOR2_X1 _27335_ (.A1(_04181_),
    .A2(_04984_),
    .ZN(_04985_));
 AOI21_X1 _27336_ (.A(_04213_),
    .B1(_04121_),
    .B2(_04115_),
    .ZN(_04986_));
 AOI22_X1 _27337_ (.A1(_04229_),
    .A2(_04208_),
    .B1(_04213_),
    .B2(_04019_),
    .ZN(_04987_));
 OAI33_X1 _27338_ (.A1(_04212_),
    .A2(_04033_),
    .A3(_04986_),
    .B1(_04987_),
    .B2(_04957_),
    .B3(_04198_),
    .ZN(_04988_));
 AOI21_X1 _27339_ (.A(_04985_),
    .B1(_04988_),
    .B2(_04470_),
    .ZN(_04989_));
 AOI21_X1 _27340_ (.A(_04086_),
    .B1(_04389_),
    .B2(_04193_),
    .ZN(_04990_));
 AOI21_X1 _27341_ (.A(_04990_),
    .B1(_04376_),
    .B2(_04614_),
    .ZN(_04991_));
 MUX2_X1 _27342_ (.A(_04035_),
    .B(_04991_),
    .S(_04198_),
    .Z(_04992_));
 AOI21_X1 _27343_ (.A(_04467_),
    .B1(_04989_),
    .B2(_04992_),
    .ZN(_04993_));
 OAI33_X1 _27344_ (.A1(_04070_),
    .A2(_04478_),
    .A3(_04125_),
    .B1(_04482_),
    .B2(_04055_),
    .B3(_04112_),
    .ZN(_04994_));
 OAI21_X1 _27345_ (.A(_04479_),
    .B1(_04129_),
    .B2(_04182_),
    .ZN(_04995_));
 AOI221_X2 _27346_ (.A(_04994_),
    .B1(_04156_),
    .B2(_04162_),
    .C1(_04462_),
    .C2(_04995_),
    .ZN(_04996_));
 NOR2_X1 _27347_ (.A1(_04072_),
    .A2(_04478_),
    .ZN(_04997_));
 NAND3_X1 _27348_ (.A1(_04451_),
    .A2(_04452_),
    .A3(_04246_),
    .ZN(_04998_));
 OAI21_X1 _27349_ (.A(_04998_),
    .B1(_04518_),
    .B2(_04197_),
    .ZN(_04999_));
 AOI21_X1 _27350_ (.A(_04997_),
    .B1(_04999_),
    .B2(_04072_),
    .ZN(_05000_));
 OAI21_X2 _27351_ (.A(_04996_),
    .B1(_05000_),
    .B2(_04500_),
    .ZN(_05001_));
 NOR3_X2 _27352_ (.A1(_04983_),
    .A2(_04993_),
    .A3(_05001_),
    .ZN(_05002_));
 NAND2_X4 _27353_ (.A1(_04966_),
    .A2(_05002_),
    .ZN(_05003_));
 XNOR2_X1 _27354_ (.A(\block_reg[0][29] ),
    .B(_04288_),
    .ZN(_05004_));
 OAI22_X1 _27355_ (.A1(_16555_),
    .A2(_04289_),
    .B1(_05004_),
    .B2(_18552_),
    .ZN(_05005_));
 NOR2_X1 _27356_ (.A1(_05003_),
    .A2(_05005_),
    .ZN(_05006_));
 XNOR2_X2 _27357_ (.A(_04311_),
    .B(_04590_),
    .ZN(_05007_));
 XNOR2_X2 _27358_ (.A(_04699_),
    .B(_04723_),
    .ZN(_05008_));
 XNOR2_X2 _27359_ (.A(_04820_),
    .B(_05008_),
    .ZN(_05009_));
 XNOR2_X1 _27360_ (.A(_05007_),
    .B(_05009_),
    .ZN(_05010_));
 XNOR2_X1 _27361_ (.A(_18064_),
    .B(_04941_),
    .ZN(_05011_));
 XNOR2_X1 _27362_ (.A(_04729_),
    .B(_05011_),
    .ZN(_05012_));
 XNOR2_X1 _27363_ (.A(_04684_),
    .B(_05012_),
    .ZN(_05013_));
 XNOR2_X2 _27364_ (.A(_05010_),
    .B(_05013_),
    .ZN(_05014_));
 XNOR2_X2 _27365_ (.A(_18410_),
    .B(_03857_),
    .ZN(_05015_));
 XNOR2_X2 _27366_ (.A(_03724_),
    .B(_04914_),
    .ZN(_05016_));
 XNOR2_X1 _27367_ (.A(_05015_),
    .B(_05016_),
    .ZN(_05017_));
 XNOR2_X2 _27368_ (.A(_05014_),
    .B(_05017_),
    .ZN(_05018_));
 OAI21_X1 _27369_ (.A(_05006_),
    .B1(_05018_),
    .B2(_17204_),
    .ZN(_05019_));
 MUX2_X1 _27370_ (.A(\core.dec_block.block_w0_reg[29] ),
    .B(_05019_),
    .S(_16365_),
    .Z(_00588_));
 NOR2_X1 _27371_ (.A1(\core.dec_block.block_w0_reg[2] ),
    .A2(_18330_),
    .ZN(_05020_));
 BUF_X4 _27372_ (.A(_16555_),
    .Z(_05021_));
 OAI21_X1 _27373_ (.A(_18329_),
    .B1(_05021_),
    .B2(_04699_),
    .ZN(_05022_));
 NAND2_X2 _27374_ (.A1(_00239_),
    .A2(_16548_),
    .ZN(_05023_));
 AOI222_X2 _27375_ (.A1(\core.keymem.key_mem[12][66] ),
    .A2(_17093_),
    .B1(_16507_),
    .B2(\core.keymem.key_mem[11][66] ),
    .C1(_16469_),
    .C2(\core.keymem.key_mem[5][66] ),
    .ZN(_05024_));
 AOI22_X2 _27376_ (.A1(\core.keymem.key_mem[14][66] ),
    .A2(_17581_),
    .B1(_16522_),
    .B2(\core.keymem.key_mem[6][66] ),
    .ZN(_05025_));
 AOI22_X2 _27377_ (.A1(\core.keymem.key_mem[8][66] ),
    .A2(_17765_),
    .B1(_17585_),
    .B2(\core.keymem.key_mem[9][66] ),
    .ZN(_05026_));
 NAND3_X2 _27378_ (.A1(_05024_),
    .A2(_05025_),
    .A3(_05026_),
    .ZN(_05027_));
 AOI22_X1 _27379_ (.A1(\core.keymem.key_mem[10][66] ),
    .A2(_16516_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][66] ),
    .ZN(_05028_));
 AOI21_X1 _27380_ (.A(_16872_),
    .B1(_17085_),
    .B2(\core.keymem.key_mem[7][66] ),
    .ZN(_05029_));
 AOI22_X2 _27381_ (.A1(\core.keymem.key_mem[2][66] ),
    .A2(_16425_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][66] ),
    .ZN(_05030_));
 AOI22_X2 _27382_ (.A1(\core.keymem.key_mem[4][66] ),
    .A2(_16501_),
    .B1(_16387_),
    .B2(\core.keymem.key_mem[3][66] ),
    .ZN(_05031_));
 NAND4_X2 _27383_ (.A1(_05028_),
    .A2(_05029_),
    .A3(_05030_),
    .A4(_05031_),
    .ZN(_05032_));
 OAI21_X4 _27384_ (.A(_05023_),
    .B1(_05027_),
    .B2(_05032_),
    .ZN(_05033_));
 XNOR2_X1 _27385_ (.A(\block_reg[1][2] ),
    .B(_05033_),
    .ZN(_05034_));
 AOI21_X1 _27386_ (.A(_05022_),
    .B1(_05034_),
    .B2(_16372_),
    .ZN(_05035_));
 NAND2_X1 _27387_ (.A1(_16794_),
    .A2(_16847_),
    .ZN(_05036_));
 AOI21_X1 _27388_ (.A(_05036_),
    .B1(_03382_),
    .B2(_16793_),
    .ZN(_05037_));
 AOI21_X1 _27389_ (.A(_05037_),
    .B1(_16723_),
    .B2(_16717_),
    .ZN(_05038_));
 NOR2_X1 _27390_ (.A1(_16828_),
    .A2(_16712_),
    .ZN(_05039_));
 MUX2_X1 _27391_ (.A(_05039_),
    .B(_03382_),
    .S(_05036_),
    .Z(_05040_));
 MUX2_X1 _27392_ (.A(_05038_),
    .B(_05040_),
    .S(_16714_),
    .Z(_05041_));
 NOR2_X1 _27393_ (.A1(_16678_),
    .A2(_05041_),
    .ZN(_05042_));
 NOR3_X1 _27394_ (.A1(_16689_),
    .A2(_16694_),
    .A3(_16800_),
    .ZN(_05043_));
 OAI22_X2 _27395_ (.A1(_16738_),
    .A2(_03470_),
    .B1(_16800_),
    .B2(_16724_),
    .ZN(_05044_));
 NAND2_X1 _27396_ (.A1(_16644_),
    .A2(_16828_),
    .ZN(_05045_));
 OAI22_X2 _27397_ (.A1(_16681_),
    .A2(_05045_),
    .B1(_03397_),
    .B2(_16844_),
    .ZN(_05046_));
 AOI221_X2 _27398_ (.A(_05043_),
    .B1(_05044_),
    .B2(_16722_),
    .C1(_16705_),
    .C2(_05046_),
    .ZN(_05047_));
 NOR2_X1 _27399_ (.A1(_16737_),
    .A2(_16639_),
    .ZN(_05048_));
 AOI21_X1 _27400_ (.A(_05048_),
    .B1(_03449_),
    .B2(_16760_),
    .ZN(_05049_));
 OAI21_X2 _27401_ (.A(_05047_),
    .B1(_05049_),
    .B2(_16726_),
    .ZN(_05050_));
 NOR3_X2 _27402_ (.A1(_16807_),
    .A2(_05042_),
    .A3(_05050_),
    .ZN(_05051_));
 NOR2_X1 _27403_ (.A1(_16796_),
    .A2(_16699_),
    .ZN(_05052_));
 AOI21_X1 _27404_ (.A(_03366_),
    .B1(_16845_),
    .B2(_16685_),
    .ZN(_05053_));
 OAI21_X1 _27405_ (.A(_16666_),
    .B1(_05052_),
    .B2(_05053_),
    .ZN(_05054_));
 NAND3_X1 _27406_ (.A1(_03399_),
    .A2(_03454_),
    .A3(_05054_),
    .ZN(_05055_));
 OAI22_X1 _27407_ (.A1(_16655_),
    .A2(_16738_),
    .B1(_16713_),
    .B2(_16803_),
    .ZN(_05056_));
 NAND3_X1 _27408_ (.A1(_16714_),
    .A2(_16799_),
    .A3(_05056_),
    .ZN(_05057_));
 OAI21_X2 _27409_ (.A(_16845_),
    .B1(_16631_),
    .B2(_16667_),
    .ZN(_05058_));
 AOI21_X1 _27410_ (.A(_16836_),
    .B1(_05058_),
    .B2(_16706_),
    .ZN(_05059_));
 AOI21_X1 _27411_ (.A(_03386_),
    .B1(_16685_),
    .B2(_16793_),
    .ZN(_05060_));
 AOI21_X1 _27412_ (.A(_16800_),
    .B1(_03382_),
    .B2(_16845_),
    .ZN(_05061_));
 OAI21_X1 _27413_ (.A(_16811_),
    .B1(_05060_),
    .B2(_05061_),
    .ZN(_05062_));
 CLKBUF_X3 _27414_ (.A(_16834_),
    .Z(_05063_));
 XNOR2_X1 _27415_ (.A(_16715_),
    .B(_16775_),
    .ZN(_05064_));
 OAI22_X1 _27416_ (.A1(_16691_),
    .A2(_16713_),
    .B1(_05064_),
    .B2(_16604_),
    .ZN(_05065_));
 NAND2_X1 _27417_ (.A1(_05063_),
    .A2(_05065_),
    .ZN(_05066_));
 NAND4_X1 _27418_ (.A1(_05057_),
    .A2(_05059_),
    .A3(_05062_),
    .A4(_05066_),
    .ZN(_05067_));
 NOR3_X1 _27419_ (.A1(_16663_),
    .A2(_16703_),
    .A3(_16710_),
    .ZN(_05068_));
 NOR2_X1 _27420_ (.A1(_03366_),
    .A2(_16785_),
    .ZN(_05069_));
 AOI21_X2 _27421_ (.A(_05068_),
    .B1(_05069_),
    .B2(_16603_),
    .ZN(_05070_));
 OAI21_X1 _27422_ (.A(_03381_),
    .B1(_03386_),
    .B2(_16821_),
    .ZN(_05071_));
 NAND4_X1 _27423_ (.A1(_16808_),
    .A2(_16810_),
    .A3(_16636_),
    .A4(_05071_),
    .ZN(_05072_));
 NAND2_X1 _27424_ (.A1(_05070_),
    .A2(_05072_),
    .ZN(_05073_));
 OAI33_X1 _27425_ (.A1(_16834_),
    .A2(_16680_),
    .A3(_16825_),
    .B1(_16727_),
    .B2(_16811_),
    .B3(_16793_),
    .ZN(_05074_));
 AOI21_X2 _27426_ (.A(_05073_),
    .B1(_05074_),
    .B2(_03466_),
    .ZN(_05075_));
 OAI22_X2 _27427_ (.A1(_03386_),
    .A2(_16841_),
    .B1(_16800_),
    .B2(_16699_),
    .ZN(_05076_));
 OAI21_X1 _27428_ (.A(_03461_),
    .B1(_16798_),
    .B2(_16793_),
    .ZN(_05077_));
 OAI21_X1 _27429_ (.A(_03479_),
    .B1(_03470_),
    .B2(_05064_),
    .ZN(_05078_));
 AOI221_X2 _27430_ (.A(_05076_),
    .B1(_05077_),
    .B2(_16782_),
    .C1(_16822_),
    .C2(_05078_),
    .ZN(_05079_));
 AOI21_X1 _27431_ (.A(_16770_),
    .B1(_16796_),
    .B2(_16587_),
    .ZN(_05080_));
 NOR2_X1 _27432_ (.A1(_16808_),
    .A2(_16821_),
    .ZN(_05081_));
 AOI21_X1 _27433_ (.A(_05080_),
    .B1(_05081_),
    .B2(_16741_),
    .ZN(_05082_));
 NOR3_X1 _27434_ (.A1(_16810_),
    .A2(_16670_),
    .A3(_05082_),
    .ZN(_05083_));
 NAND2_X1 _27435_ (.A1(_16808_),
    .A2(_16821_),
    .ZN(_05084_));
 OAI22_X1 _27436_ (.A1(_16691_),
    .A2(_05084_),
    .B1(_16816_),
    .B2(_16676_),
    .ZN(_05085_));
 AND3_X1 _27437_ (.A1(_16810_),
    .A2(_16670_),
    .A3(_05085_),
    .ZN(_05086_));
 OAI21_X1 _27438_ (.A(_16733_),
    .B1(_05083_),
    .B2(_05086_),
    .ZN(_05087_));
 OAI22_X1 _27439_ (.A1(_16759_),
    .A2(_16841_),
    .B1(_16800_),
    .B2(_16732_),
    .ZN(_05088_));
 NAND3_X1 _27440_ (.A1(_16656_),
    .A2(_16667_),
    .A3(_16717_),
    .ZN(_05089_));
 OAI21_X1 _27441_ (.A(_05089_),
    .B1(_16672_),
    .B2(_16656_),
    .ZN(_05090_));
 AOI21_X2 _27442_ (.A(_05088_),
    .B1(_05090_),
    .B2(_03447_),
    .ZN(_05091_));
 NAND4_X2 _27443_ (.A1(_05075_),
    .A2(_05079_),
    .A3(_05087_),
    .A4(_05091_),
    .ZN(_05092_));
 NAND3_X1 _27444_ (.A1(_16767_),
    .A2(_16613_),
    .A3(_16710_),
    .ZN(_05093_));
 AOI22_X1 _27445_ (.A1(_16673_),
    .A2(_16745_),
    .B1(_16747_),
    .B2(_16798_),
    .ZN(_05094_));
 OAI21_X1 _27446_ (.A(_05093_),
    .B1(_05094_),
    .B2(_16767_),
    .ZN(_05095_));
 NAND2_X2 _27447_ (.A1(_16632_),
    .A2(_16638_),
    .ZN(_05096_));
 NAND3_X1 _27448_ (.A1(_16811_),
    .A2(_16677_),
    .A3(_16717_),
    .ZN(_05097_));
 AOI21_X1 _27449_ (.A(_16767_),
    .B1(_05096_),
    .B2(_05097_),
    .ZN(_05098_));
 MUX2_X2 _27450_ (.A(_05095_),
    .B(_05098_),
    .S(_16714_),
    .Z(_05099_));
 NOR4_X2 _27451_ (.A1(_05055_),
    .A2(_05067_),
    .A3(_05092_),
    .A4(_05099_),
    .ZN(_05100_));
 NAND2_X4 _27452_ (.A1(_05051_),
    .A2(_05100_),
    .ZN(_05101_));
 AND2_X1 _27453_ (.A1(\core.keymem.key_mem[14][79] ),
    .A2(_17025_),
    .ZN(_05102_));
 INV_X1 _27454_ (.A(\core.keymem.key_mem[13][79] ),
    .ZN(_05103_));
 AOI21_X1 _27455_ (.A(_05103_),
    .B1(_16411_),
    .B2(_16413_),
    .ZN(_05104_));
 OAI21_X1 _27456_ (.A(_17099_),
    .B1(_05102_),
    .B2(_05104_),
    .ZN(_05105_));
 AOI21_X1 _27457_ (.A(_16544_),
    .B1(_16858_),
    .B2(\core.keymem.key_mem[2][79] ),
    .ZN(_05106_));
 AOI22_X1 _27458_ (.A1(\core.keymem.key_mem[4][79] ),
    .A2(_16455_),
    .B1(_16396_),
    .B2(\core.keymem.key_mem[12][79] ),
    .ZN(_05107_));
 AOI22_X1 _27459_ (.A1(\core.keymem.key_mem[9][79] ),
    .A2(_16460_),
    .B1(_16431_),
    .B2(\core.keymem.key_mem[10][79] ),
    .ZN(_05108_));
 AND4_X1 _27460_ (.A1(_05105_),
    .A2(_05106_),
    .A3(_05107_),
    .A4(_05108_),
    .ZN(_05109_));
 AOI22_X1 _27461_ (.A1(\core.keymem.key_mem[7][79] ),
    .A2(_16954_),
    .B1(_16519_),
    .B2(\core.keymem.key_mem[6][79] ),
    .ZN(_05110_));
 AOI222_X2 _27462_ (.A1(\core.keymem.key_mem[11][79] ),
    .A2(_16504_),
    .B1(_16523_),
    .B2(\core.keymem.key_mem[1][79] ),
    .C1(_16466_),
    .C2(\core.keymem.key_mem[5][79] ),
    .ZN(_05111_));
 AOI22_X1 _27463_ (.A1(\core.keymem.key_mem[8][79] ),
    .A2(_16451_),
    .B1(_16864_),
    .B2(\core.keymem.key_mem[3][79] ),
    .ZN(_05112_));
 AND3_X1 _27464_ (.A1(_05110_),
    .A2(_05111_),
    .A3(_05112_),
    .ZN(_05113_));
 AOI22_X4 _27465_ (.A1(_00222_),
    .A2(_17013_),
    .B1(_05109_),
    .B2(_05113_),
    .ZN(_05114_));
 XNOR2_X2 _27466_ (.A(\core.dec_block.block_w1_reg[15] ),
    .B(_05114_),
    .ZN(_05115_));
 XNOR2_X2 _27467_ (.A(_03596_),
    .B(_05115_),
    .ZN(_05116_));
 AND2_X1 _27468_ (.A1(_00236_),
    .A2(_16983_),
    .ZN(_05117_));
 OAI211_X2 _27469_ (.A(\core.keymem.key_mem[11][90] ),
    .B(_17112_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_05118_));
 NAND3_X1 _27470_ (.A1(\core.keymem.key_mem[2][90] ),
    .A2(_17121_),
    .A3(_17101_),
    .ZN(_05119_));
 OAI211_X2 _27471_ (.A(\core.keymem.key_mem[7][90] ),
    .B(_17112_),
    .C1(_17107_),
    .C2(_17106_),
    .ZN(_05120_));
 OAI211_X2 _27472_ (.A(\core.keymem.key_mem[6][90] ),
    .B(_17050_),
    .C1(_17106_),
    .C2(_17107_),
    .ZN(_05121_));
 NAND4_X2 _27473_ (.A1(_05118_),
    .A2(_05119_),
    .A3(_05120_),
    .A4(_05121_),
    .ZN(_05122_));
 OAI211_X2 _27474_ (.A(\core.keymem.key_mem[4][90] ),
    .B(_17057_),
    .C1(_17114_),
    .C2(_17115_),
    .ZN(_05123_));
 OAI211_X2 _27475_ (.A(\core.keymem.key_mem[13][90] ),
    .B(_17100_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_05124_));
 NAND3_X1 _27476_ (.A1(\core.keymem.key_mem[3][90] ),
    .A2(_17048_),
    .A3(_16970_),
    .ZN(_05125_));
 OAI211_X2 _27477_ (.A(\core.keymem.key_mem[1][90] ),
    .B(_16970_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_05126_));
 NAND4_X2 _27478_ (.A1(_05123_),
    .A2(_05124_),
    .A3(_05125_),
    .A4(_05126_),
    .ZN(_05127_));
 OAI211_X2 _27479_ (.A(\core.keymem.key_mem[10][90] ),
    .B(_17050_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_05128_));
 NAND3_X1 _27480_ (.A1(\core.keymem.key_mem[14][90] ),
    .A2(_17100_),
    .A3(_17016_),
    .ZN(_05129_));
 OAI211_X2 _27481_ (.A(\core.keymem.key_mem[8][90] ),
    .B(_17527_),
    .C1(_17128_),
    .C2(_17129_),
    .ZN(_05130_));
 OAI221_X2 _27482_ (.A(\core.keymem.key_mem[9][90] ),
    .B1(_16886_),
    .B2(_16890_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_05131_));
 NAND4_X2 _27483_ (.A1(_05128_),
    .A2(_05129_),
    .A3(_05130_),
    .A4(_05131_),
    .ZN(_05132_));
 INV_X1 _27484_ (.A(\core.keymem.key_mem[12][90] ),
    .ZN(_05133_));
 INV_X1 _27485_ (.A(\core.keymem.key_mem[5][90] ),
    .ZN(_05134_));
 OAI22_X2 _27486_ (.A1(_05133_),
    .A2(_17843_),
    .B1(_03591_),
    .B2(_05134_),
    .ZN(_05135_));
 NOR4_X4 _27487_ (.A1(_05122_),
    .A2(_05127_),
    .A3(_05132_),
    .A4(_05135_),
    .ZN(_05136_));
 AOI21_X4 _27488_ (.A(_05117_),
    .B1(_05136_),
    .B2(_17533_),
    .ZN(_05137_));
 XNOR2_X2 _27489_ (.A(\core.dec_block.block_w1_reg[26] ),
    .B(_05137_),
    .ZN(_05138_));
 INV_X1 _27490_ (.A(_00240_),
    .ZN(_05139_));
 NAND3_X1 _27491_ (.A1(\core.keymem.key_mem[3][74] ),
    .A2(_17111_),
    .A3(_17120_),
    .ZN(_05140_));
 OAI221_X1 _27492_ (.A(\core.keymem.key_mem[9][74] ),
    .B1(_16927_),
    .B2(_16929_),
    .C1(_17143_),
    .C2(_17144_),
    .ZN(_05141_));
 OAI211_X2 _27493_ (.A(\core.keymem.key_mem[10][74] ),
    .B(_17026_),
    .C1(_16886_),
    .C2(_16890_),
    .ZN(_05142_));
 NAND3_X1 _27494_ (.A1(\core.keymem.key_mem[2][74] ),
    .A2(_17120_),
    .A3(_17026_),
    .ZN(_05143_));
 AND4_X1 _27495_ (.A1(_05140_),
    .A2(_05141_),
    .A3(_05142_),
    .A4(_05143_),
    .ZN(_05144_));
 OAI211_X2 _27496_ (.A(\core.keymem.key_mem[4][74] ),
    .B(_17028_),
    .C1(_17146_),
    .C2(_17031_),
    .ZN(_05145_));
 NAND3_X1 _27497_ (.A1(\core.keymem.key_mem[12][74] ),
    .A2(_17024_),
    .A3(_17527_),
    .ZN(_05146_));
 OAI211_X2 _27498_ (.A(\core.keymem.key_mem[13][74] ),
    .B(_17099_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_05147_));
 OAI221_X1 _27499_ (.A(\core.keymem.key_mem[5][74] ),
    .B1(_16908_),
    .B2(_16917_),
    .C1(_17149_),
    .C2(_16915_),
    .ZN(_05148_));
 AND4_X1 _27500_ (.A1(_05145_),
    .A2(_05146_),
    .A3(_05147_),
    .A4(_05148_),
    .ZN(_05149_));
 OAI211_X2 _27501_ (.A(\core.keymem.key_mem[6][74] ),
    .B(_17026_),
    .C1(_17622_),
    .C2(_17030_),
    .ZN(_05150_));
 OAI211_X2 _27502_ (.A(\core.keymem.key_mem[11][74] ),
    .B(_17074_),
    .C1(_17035_),
    .C2(_17036_),
    .ZN(_05151_));
 OAI211_X2 _27503_ (.A(\core.keymem.key_mem[1][74] ),
    .B(_17827_),
    .C1(_17149_),
    .C2(_17117_),
    .ZN(_05152_));
 OAI211_X2 _27504_ (.A(\core.keymem.key_mem[8][74] ),
    .B(_16893_),
    .C1(_17035_),
    .C2(_17036_),
    .ZN(_05153_));
 AND4_X1 _27505_ (.A1(_05150_),
    .A2(_05151_),
    .A3(_05152_),
    .A4(_05153_),
    .ZN(_05154_));
 AOI22_X4 _27506_ (.A1(\core.keymem.key_mem[14][74] ),
    .A2(_16998_),
    .B1(_16407_),
    .B2(\core.keymem.key_mem[7][74] ),
    .ZN(_05155_));
 NAND4_X4 _27507_ (.A1(_05144_),
    .A2(_05149_),
    .A3(_05154_),
    .A4(_05155_),
    .ZN(_05156_));
 MUX2_X2 _27508_ (.A(_05139_),
    .B(_05156_),
    .S(_16488_),
    .Z(_05157_));
 XNOR2_X2 _27509_ (.A(\core.dec_block.block_w1_reg[10] ),
    .B(_05157_),
    .ZN(_05158_));
 XNOR2_X1 _27510_ (.A(_05138_),
    .B(_05158_),
    .ZN(_05159_));
 XNOR2_X1 _27511_ (.A(_05116_),
    .B(_05159_),
    .ZN(_05160_));
 XNOR2_X2 _27512_ (.A(_03542_),
    .B(_05160_),
    .ZN(_05161_));
 XNOR2_X2 _27513_ (.A(_17139_),
    .B(_03525_),
    .ZN(_05162_));
 XNOR2_X1 _27514_ (.A(_16978_),
    .B(_05162_),
    .ZN(_05163_));
 XNOR2_X1 _27515_ (.A(_05161_),
    .B(_05163_),
    .ZN(_05164_));
 AOI222_X2 _27516_ (.A1(\core.keymem.key_mem[4][82] ),
    .A2(_16457_),
    .B1(_16512_),
    .B2(\core.keymem.key_mem[7][82] ),
    .C1(\core.keymem.key_mem[8][82] ),
    .C2(_16452_),
    .ZN(_05165_));
 AOI22_X1 _27517_ (.A1(\core.keymem.key_mem[10][82] ),
    .A2(_16989_),
    .B1(_17720_),
    .B2(\core.keymem.key_mem[12][82] ),
    .ZN(_05166_));
 AOI22_X1 _27518_ (.A1(\core.keymem.key_mem[9][82] ),
    .A2(_17668_),
    .B1(_17722_),
    .B2(\core.keymem.key_mem[13][82] ),
    .ZN(_05167_));
 NAND3_X1 _27519_ (.A1(_05165_),
    .A2(_05166_),
    .A3(_05167_),
    .ZN(_05168_));
 AOI22_X1 _27520_ (.A1(\core.keymem.key_mem[2][82] ),
    .A2(_17786_),
    .B1(_16509_),
    .B2(\core.keymem.key_mem[5][82] ),
    .ZN(_05169_));
 AOI22_X1 _27521_ (.A1(\core.keymem.key_mem[3][82] ),
    .A2(_16866_),
    .B1(_16506_),
    .B2(\core.keymem.key_mem[11][82] ),
    .ZN(_05170_));
 AOI22_X1 _27522_ (.A1(\core.keymem.key_mem[14][82] ),
    .A2(_17719_),
    .B1(_16855_),
    .B2(\core.keymem.key_mem[1][82] ),
    .ZN(_05171_));
 AOI21_X1 _27523_ (.A(_16495_),
    .B1(_17695_),
    .B2(\core.keymem.key_mem[6][82] ),
    .ZN(_05172_));
 NAND4_X1 _27524_ (.A1(_05169_),
    .A2(_05170_),
    .A3(_05171_),
    .A4(_05172_),
    .ZN(_05173_));
 NOR2_X2 _27525_ (.A1(_05168_),
    .A2(_05173_),
    .ZN(_05174_));
 AOI21_X4 _27526_ (.A(_05174_),
    .B1(_17183_),
    .B2(_00238_),
    .ZN(_05175_));
 XNOR2_X2 _27527_ (.A(\core.dec_block.block_w1_reg[18] ),
    .B(_05175_),
    .ZN(_05176_));
 XNOR2_X2 _27528_ (.A(\core.dec_block.block_w1_reg[1] ),
    .B(_03520_),
    .ZN(_05177_));
 XNOR2_X2 _27529_ (.A(_05176_),
    .B(_05177_),
    .ZN(_05178_));
 XNOR2_X1 _27530_ (.A(_16875_),
    .B(_03556_),
    .ZN(_05179_));
 XOR2_X1 _27531_ (.A(_05178_),
    .B(_05179_),
    .Z(_05180_));
 XNOR2_X1 _27532_ (.A(_05164_),
    .B(_05180_),
    .ZN(_05181_));
 AOI21_X1 _27533_ (.A(_05101_),
    .B1(_05181_),
    .B2(_19031_),
    .ZN(_05182_));
 AOI21_X1 _27534_ (.A(_05020_),
    .B1(_05035_),
    .B2(_05182_),
    .ZN(_00589_));
 XNOR2_X2 _27535_ (.A(_04914_),
    .B(_04942_),
    .ZN(_05183_));
 XNOR2_X2 _27536_ (.A(_04804_),
    .B(_04833_),
    .ZN(_05184_));
 XOR2_X1 _27537_ (.A(_04349_),
    .B(_05184_),
    .Z(_05185_));
 XNOR2_X1 _27538_ (.A(_04819_),
    .B(_05185_),
    .ZN(_05186_));
 XNOR2_X1 _27539_ (.A(_05183_),
    .B(_05186_),
    .ZN(_05187_));
 XNOR2_X2 _27540_ (.A(_03857_),
    .B(_04289_),
    .ZN(_05188_));
 XNOR2_X1 _27541_ (.A(_04724_),
    .B(_05188_),
    .ZN(_05189_));
 XNOR2_X2 _27542_ (.A(_18478_),
    .B(_03915_),
    .ZN(_05190_));
 XOR2_X1 _27543_ (.A(_18326_),
    .B(_05190_),
    .Z(_05191_));
 XNOR2_X1 _27544_ (.A(_05189_),
    .B(_05191_),
    .ZN(_05192_));
 XNOR2_X1 _27545_ (.A(_05187_),
    .B(_05192_),
    .ZN(_05193_));
 INV_X1 _27546_ (.A(\block_reg[0][30] ),
    .ZN(_05194_));
 XNOR2_X2 _27547_ (.A(_05194_),
    .B(_04310_),
    .ZN(_05195_));
 OAI222_X2 _27548_ (.A1(_16556_),
    .A2(_04311_),
    .B1(_05193_),
    .B2(_17203_),
    .C1(_05195_),
    .C2(_18412_),
    .ZN(_05196_));
 AOI22_X2 _27549_ (.A1(_04198_),
    .A2(_04246_),
    .B1(_04533_),
    .B2(_04025_),
    .ZN(_05197_));
 OAI22_X2 _27550_ (.A1(_04222_),
    .A2(_04223_),
    .B1(_05197_),
    .B2(_04143_),
    .ZN(_05198_));
 NAND3_X1 _27551_ (.A1(_04132_),
    .A2(_04452_),
    .A3(_04246_),
    .ZN(_05199_));
 OAI21_X1 _27552_ (.A(_04451_),
    .B1(_04186_),
    .B2(_04139_),
    .ZN(_05200_));
 AOI21_X2 _27553_ (.A(_04441_),
    .B1(_05199_),
    .B2(_05200_),
    .ZN(_05201_));
 AOI21_X1 _27554_ (.A(_04111_),
    .B1(_04065_),
    .B2(_04478_),
    .ZN(_05202_));
 OAI21_X1 _27555_ (.A(_04191_),
    .B1(_04476_),
    .B2(_05202_),
    .ZN(_05203_));
 NOR3_X1 _27556_ (.A1(_04084_),
    .A2(_04061_),
    .A3(_04459_),
    .ZN(_05204_));
 NOR3_X1 _27557_ (.A1(_04058_),
    .A2(_04104_),
    .A3(_04510_),
    .ZN(_05205_));
 OAI21_X1 _27558_ (.A(_04071_),
    .B1(_05204_),
    .B2(_05205_),
    .ZN(_05206_));
 NAND4_X1 _27559_ (.A1(_04037_),
    .A2(_04612_),
    .A3(_05203_),
    .A4(_05206_),
    .ZN(_05207_));
 NOR4_X2 _27560_ (.A1(_04790_),
    .A2(_05198_),
    .A3(_05201_),
    .A4(_05207_),
    .ZN(_05208_));
 NOR4_X1 _27561_ (.A1(_04084_),
    .A2(_04059_),
    .A3(_04047_),
    .A4(_04130_),
    .ZN(_05209_));
 AND2_X1 _27562_ (.A1(_04244_),
    .A2(_04168_),
    .ZN(_05210_));
 AOI21_X1 _27563_ (.A(_05209_),
    .B1(_05210_),
    .B2(_04068_),
    .ZN(_05211_));
 AOI21_X1 _27564_ (.A(_04463_),
    .B1(_04188_),
    .B2(_04091_),
    .ZN(_05212_));
 AOI21_X1 _27565_ (.A(_03996_),
    .B1(_04148_),
    .B2(_04193_),
    .ZN(_05213_));
 AOI21_X1 _27566_ (.A(_05213_),
    .B1(_04461_),
    .B2(_04452_),
    .ZN(_05214_));
 OAI221_X2 _27567_ (.A(_05211_),
    .B1(_05212_),
    .B2(_04223_),
    .C1(_04182_),
    .C2(_05214_),
    .ZN(_05215_));
 NOR3_X1 _27568_ (.A1(_04886_),
    .A2(_04890_),
    .A3(_05215_),
    .ZN(_05216_));
 NAND2_X2 _27569_ (.A1(_05208_),
    .A2(_05216_),
    .ZN(_05217_));
 OAI21_X1 _27570_ (.A(_04201_),
    .B1(_04478_),
    .B2(_04084_),
    .ZN(_05218_));
 AOI21_X1 _27571_ (.A(_04100_),
    .B1(_04110_),
    .B2(_04070_),
    .ZN(_05219_));
 NOR2_X1 _27572_ (.A1(_04142_),
    .A2(_05219_),
    .ZN(_05220_));
 AOI221_X2 _27573_ (.A(_04452_),
    .B1(_04101_),
    .B2(_05218_),
    .C1(_05220_),
    .C2(_04132_),
    .ZN(_05221_));
 AOI21_X1 _27574_ (.A(_04115_),
    .B1(_04086_),
    .B2(_04142_),
    .ZN(_05222_));
 OAI22_X1 _27575_ (.A1(_04148_),
    .A2(_04441_),
    .B1(_04187_),
    .B2(_04071_),
    .ZN(_05223_));
 AOI221_X2 _27576_ (.A(_04614_),
    .B1(_04462_),
    .B2(_05222_),
    .C1(_05223_),
    .C2(_04451_),
    .ZN(_05224_));
 OAI21_X2 _27577_ (.A(_04144_),
    .B1(_05221_),
    .B2(_05224_),
    .ZN(_05225_));
 NOR4_X4 _27578_ (.A1(_04448_),
    .A2(_05001_),
    .A3(_05217_),
    .A4(_05225_),
    .ZN(_05226_));
 AOI21_X4 _27579_ (.A(_17379_),
    .B1(_04465_),
    .B2(_05226_),
    .ZN(_05227_));
 OAI21_X1 _27580_ (.A(_16366_),
    .B1(_05196_),
    .B2(_05227_),
    .ZN(_05228_));
 OAI21_X1 _27581_ (.A(_05228_),
    .B1(_16366_),
    .B2(_04290_),
    .ZN(_00590_));
 NOR2_X1 _27582_ (.A1(_04003_),
    .A2(_16365_),
    .ZN(_05229_));
 NOR2_X1 _27583_ (.A1(_04883_),
    .A2(_05215_),
    .ZN(_05230_));
 NOR2_X1 _27584_ (.A1(_04376_),
    .A2(_04157_),
    .ZN(_05231_));
 NOR2_X1 _27585_ (.A1(_04069_),
    .A2(_04510_),
    .ZN(_05232_));
 OAI33_X1 _27586_ (.A1(_04151_),
    .A2(_04407_),
    .A3(_05231_),
    .B1(_05232_),
    .B2(_04057_),
    .B3(_04173_),
    .ZN(_05233_));
 OR2_X1 _27587_ (.A1(_04190_),
    .A2(_05233_),
    .ZN(_05234_));
 NAND2_X1 _27588_ (.A1(_04046_),
    .A2(_04461_),
    .ZN(_05235_));
 MUX2_X1 _27589_ (.A(_04077_),
    .B(_04104_),
    .S(_03994_),
    .Z(_05236_));
 OAI221_X2 _27590_ (.A(_05235_),
    .B1(_05236_),
    .B2(_04002_),
    .C1(_04381_),
    .C2(_04046_),
    .ZN(_05237_));
 OAI21_X1 _27591_ (.A(_04081_),
    .B1(_04135_),
    .B2(_04019_),
    .ZN(_05238_));
 AOI22_X1 _27592_ (.A1(_04050_),
    .A2(_04054_),
    .B1(_04150_),
    .B2(_05238_),
    .ZN(_05239_));
 OAI21_X1 _27593_ (.A(_04629_),
    .B1(_05239_),
    .B2(_04117_),
    .ZN(_05240_));
 AOI221_X2 _27594_ (.A(_05234_),
    .B1(_05237_),
    .B2(_03989_),
    .C1(_04207_),
    .C2(_05240_),
    .ZN(_05241_));
 AOI22_X1 _27595_ (.A1(_04083_),
    .A2(_04221_),
    .B1(_04510_),
    .B2(_04034_),
    .ZN(_05242_));
 AOI21_X1 _27596_ (.A(_04246_),
    .B1(_04188_),
    .B2(_04156_),
    .ZN(_05243_));
 AOI21_X1 _27597_ (.A(_04182_),
    .B1(_05242_),
    .B2(_05243_),
    .ZN(_05244_));
 OAI21_X1 _27598_ (.A(_03994_),
    .B1(_04083_),
    .B2(_04887_),
    .ZN(_05245_));
 AOI221_X1 _27599_ (.A(_04030_),
    .B1(_04600_),
    .B2(_05245_),
    .C1(_03986_),
    .C2(_18416_),
    .ZN(_05246_));
 NOR4_X1 _27600_ (.A1(_04782_),
    .A2(_04971_),
    .A3(_05244_),
    .A4(_05246_),
    .ZN(_05247_));
 AND4_X1 _27601_ (.A1(_04420_),
    .A2(_04454_),
    .A3(_05241_),
    .A4(_05247_),
    .ZN(_05248_));
 AOI221_X2 _27602_ (.A(_04059_),
    .B1(_03994_),
    .B2(_04029_),
    .C1(_04148_),
    .C2(_04055_),
    .ZN(_05249_));
 NAND2_X1 _27603_ (.A1(_04478_),
    .A2(_04130_),
    .ZN(_05250_));
 AOI221_X2 _27604_ (.A(_05249_),
    .B1(_04462_),
    .B2(_04048_),
    .C1(_04451_),
    .C2(_05250_),
    .ZN(_05251_));
 NOR2_X1 _27605_ (.A1(_04083_),
    .A2(_04139_),
    .ZN(_05252_));
 OAI221_X1 _27606_ (.A(_04061_),
    .B1(_05252_),
    .B2(_04191_),
    .C1(_04614_),
    .C2(_04192_),
    .ZN(_05253_));
 AOI21_X1 _27607_ (.A(_04470_),
    .B1(_05253_),
    .B2(_04072_),
    .ZN(_05254_));
 OAI21_X1 _27608_ (.A(_04174_),
    .B1(_04061_),
    .B2(_04451_),
    .ZN(_05255_));
 AOI22_X1 _27609_ (.A1(_04197_),
    .A2(_04734_),
    .B1(_05255_),
    .B2(_04181_),
    .ZN(_05256_));
 OAI22_X1 _27610_ (.A1(_05251_),
    .A2(_05254_),
    .B1(_05256_),
    .B2(_04072_),
    .ZN(_05257_));
 NAND2_X1 _27611_ (.A1(_04467_),
    .A2(_05257_),
    .ZN(_05258_));
 AND4_X4 _27612_ (.A1(_04638_),
    .A2(_05230_),
    .A3(_05248_),
    .A4(_05258_),
    .ZN(_05259_));
 XNOR2_X1 _27613_ (.A(\block_reg[0][31] ),
    .B(_04348_),
    .ZN(_05260_));
 OAI221_X1 _27614_ (.A(_05259_),
    .B1(_05260_),
    .B2(_18466_),
    .C1(_04349_),
    .C2(_18399_),
    .ZN(_05261_));
 XNOR2_X2 _27615_ (.A(_18326_),
    .B(_04937_),
    .ZN(_05262_));
 XOR2_X1 _27616_ (.A(_05016_),
    .B(_05262_),
    .Z(_05263_));
 XNOR2_X1 _27617_ (.A(_04723_),
    .B(_05263_),
    .ZN(_05264_));
 XNOR2_X2 _27618_ (.A(_18550_),
    .B(_04683_),
    .ZN(_05265_));
 XNOR2_X1 _27619_ (.A(_04313_),
    .B(_05265_),
    .ZN(_05266_));
 XNOR2_X2 _27620_ (.A(_05264_),
    .B(_05266_),
    .ZN(_05267_));
 AOI21_X1 _27621_ (.A(_05261_),
    .B1(_05267_),
    .B2(_04370_),
    .ZN(_05268_));
 AOI21_X1 _27622_ (.A(_05229_),
    .B1(_05268_),
    .B2(_16366_),
    .ZN(_00591_));
 AND2_X2 _27623_ (.A1(_00244_),
    .A2(_16984_),
    .ZN(_05269_));
 AOI22_X1 _27624_ (.A1(\core.keymem.key_mem[11][67] ),
    .A2(_16443_),
    .B1(_17003_),
    .B2(\core.keymem.key_mem[1][67] ),
    .ZN(_05270_));
 AOI22_X2 _27625_ (.A1(\core.keymem.key_mem[8][67] ),
    .A2(_17781_),
    .B1(_17914_),
    .B2(\core.keymem.key_mem[9][67] ),
    .ZN(_05271_));
 AOI22_X2 _27626_ (.A1(\core.keymem.key_mem[7][67] ),
    .A2(_17789_),
    .B1(_16989_),
    .B2(\core.keymem.key_mem[10][67] ),
    .ZN(_05272_));
 AOI21_X1 _27627_ (.A(_17013_),
    .B1(_16399_),
    .B2(\core.keymem.key_mem[12][67] ),
    .ZN(_05273_));
 NAND4_X2 _27628_ (.A1(_05270_),
    .A2(_05271_),
    .A3(_05272_),
    .A4(_05273_),
    .ZN(_05274_));
 MUX2_X1 _27629_ (.A(\core.keymem.key_mem[6][67] ),
    .B(\core.keymem.key_mem[14][67] ),
    .S(_17054_),
    .Z(_05275_));
 AOI22_X1 _27630_ (.A1(\core.keymem.key_mem[2][67] ),
    .A2(_17121_),
    .B1(_17051_),
    .B2(_05275_),
    .ZN(_05276_));
 NOR2_X1 _27631_ (.A1(_16968_),
    .A2(_05276_),
    .ZN(_05277_));
 AOI22_X1 _27632_ (.A1(\core.keymem.key_mem[4][67] ),
    .A2(_16500_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][67] ),
    .ZN(_05278_));
 AOI22_X1 _27633_ (.A1(\core.keymem.key_mem[3][67] ),
    .A2(_16987_),
    .B1(_17005_),
    .B2(\core.keymem.key_mem[5][67] ),
    .ZN(_05279_));
 NAND2_X1 _27634_ (.A1(_05278_),
    .A2(_05279_),
    .ZN(_05280_));
 NOR3_X4 _27635_ (.A1(_05274_),
    .A2(_05277_),
    .A3(_05280_),
    .ZN(_05281_));
 NOR2_X4 _27636_ (.A1(_05269_),
    .A2(_05281_),
    .ZN(_05282_));
 XNOR2_X1 _27637_ (.A(\block_reg[1][3] ),
    .B(_05282_),
    .ZN(_05283_));
 OAI221_X1 _27638_ (.A(_16365_),
    .B1(_03858_),
    .B2(_04833_),
    .C1(_05283_),
    .C2(_04266_),
    .ZN(_05284_));
 MUX2_X1 _27639_ (.A(_16638_),
    .B(_16790_),
    .S(_16714_),
    .Z(_05285_));
 NAND3_X1 _27640_ (.A1(_03466_),
    .A2(_16740_),
    .A3(_05285_),
    .ZN(_05286_));
 NOR4_X1 _27641_ (.A1(_16587_),
    .A2(_16628_),
    .A3(_16667_),
    .A4(_16683_),
    .ZN(_05287_));
 AOI21_X1 _27642_ (.A(_05287_),
    .B1(_05081_),
    .B2(_16670_),
    .ZN(_05288_));
 OAI22_X1 _27643_ (.A1(_16808_),
    .A2(_16637_),
    .B1(_05288_),
    .B2(_16803_),
    .ZN(_05289_));
 AOI22_X2 _27644_ (.A1(_16803_),
    .A2(_03402_),
    .B1(_05289_),
    .B2(_16810_),
    .ZN(_05290_));
 OAI221_X2 _27645_ (.A(_05286_),
    .B1(_05290_),
    .B2(_16785_),
    .C1(_16728_),
    .C2(_16759_),
    .ZN(_05291_));
 OAI33_X1 _27646_ (.A1(_16681_),
    .A2(_16690_),
    .A3(_16738_),
    .B1(_16699_),
    .B2(_16647_),
    .B3(_16692_),
    .ZN(_05292_));
 MUX2_X1 _27647_ (.A(_16603_),
    .B(_16789_),
    .S(_16632_),
    .Z(_05293_));
 OAI22_X2 _27648_ (.A1(_16792_),
    .A2(_16781_),
    .B1(_05096_),
    .B2(_16785_),
    .ZN(_05294_));
 AOI221_X2 _27649_ (.A(_05292_),
    .B1(_05293_),
    .B2(_16666_),
    .C1(_05294_),
    .C2(_16737_),
    .ZN(_05295_));
 NAND2_X1 _27650_ (.A1(_05075_),
    .A2(_05295_),
    .ZN(_05296_));
 NOR2_X1 _27651_ (.A1(_16735_),
    .A2(_05296_),
    .ZN(_05297_));
 OAI22_X1 _27652_ (.A1(_16737_),
    .A2(_05084_),
    .B1(_16816_),
    .B2(_16701_),
    .ZN(_05298_));
 AOI22_X1 _27653_ (.A1(_16683_),
    .A2(_03422_),
    .B1(_05298_),
    .B2(_16670_),
    .ZN(_05299_));
 NOR2_X1 _27654_ (.A1(_16657_),
    .A2(_05299_),
    .ZN(_05300_));
 NOR4_X1 _27655_ (.A1(_16810_),
    .A2(_16636_),
    .A3(_16691_),
    .A4(_05084_),
    .ZN(_05301_));
 OAI21_X1 _27656_ (.A(_16686_),
    .B1(_05300_),
    .B2(_05301_),
    .ZN(_05302_));
 NAND2_X1 _27657_ (.A1(_16613_),
    .A2(_16710_),
    .ZN(_05303_));
 OAI221_X2 _27658_ (.A(_05302_),
    .B1(_03479_),
    .B2(_16845_),
    .C1(_16736_),
    .C2(_05303_),
    .ZN(_05304_));
 AOI22_X1 _27659_ (.A1(_16803_),
    .A2(_16603_),
    .B1(_16828_),
    .B2(_16767_),
    .ZN(_05305_));
 AOI221_X1 _27660_ (.A(_16659_),
    .B1(_16745_),
    .B2(_16708_),
    .C1(_16603_),
    .C2(_16798_),
    .ZN(_05306_));
 OAI221_X1 _27661_ (.A(_05063_),
    .B1(_16811_),
    .B2(_05305_),
    .C1(_05306_),
    .C2(_03466_),
    .ZN(_05307_));
 OAI221_X1 _27662_ (.A(_16714_),
    .B1(_16799_),
    .B2(_16823_),
    .C1(_16791_),
    .C2(_16742_),
    .ZN(_05308_));
 AOI21_X1 _27663_ (.A(_05304_),
    .B1(_05307_),
    .B2(_05308_),
    .ZN(_05309_));
 NAND4_X1 _27664_ (.A1(_16770_),
    .A2(_16677_),
    .A3(_16679_),
    .A4(_16733_),
    .ZN(_05310_));
 OAI221_X2 _27665_ (.A(_05310_),
    .B1(_16732_),
    .B2(_03386_),
    .C1(_16694_),
    .C2(_16800_),
    .ZN(_05311_));
 OAI21_X1 _27666_ (.A(_03470_),
    .B1(_03446_),
    .B2(_16808_),
    .ZN(_05312_));
 NAND4_X1 _27667_ (.A1(_16810_),
    .A2(_16847_),
    .A3(_16683_),
    .A4(_05312_),
    .ZN(_05313_));
 OAI21_X1 _27668_ (.A(_05313_),
    .B1(_16727_),
    .B2(_16672_),
    .ZN(_05314_));
 AOI22_X2 _27669_ (.A1(_16811_),
    .A2(_05311_),
    .B1(_05314_),
    .B2(_03466_),
    .ZN(_05315_));
 NOR2_X1 _27670_ (.A1(_16659_),
    .A2(_16746_),
    .ZN(_05316_));
 AOI21_X1 _27671_ (.A(_16783_),
    .B1(_05316_),
    .B2(_16663_),
    .ZN(_05317_));
 OAI33_X1 _27672_ (.A1(_16663_),
    .A2(_16811_),
    .A3(_03386_),
    .B1(_03440_),
    .B2(_16680_),
    .B3(_16754_),
    .ZN(_05318_));
 AOI22_X1 _27673_ (.A1(_16666_),
    .A2(_16717_),
    .B1(_03430_),
    .B2(_16746_),
    .ZN(_05319_));
 NAND2_X1 _27674_ (.A1(_16723_),
    .A2(_16797_),
    .ZN(_05320_));
 OAI21_X1 _27675_ (.A(_05319_),
    .B1(_05320_),
    .B2(_16631_),
    .ZN(_05321_));
 NOR3_X1 _27676_ (.A1(_05317_),
    .A2(_05318_),
    .A3(_05321_),
    .ZN(_05322_));
 NAND3_X1 _27677_ (.A1(_03494_),
    .A2(_05315_),
    .A3(_05322_),
    .ZN(_05323_));
 NOR2_X2 _27678_ (.A1(_16847_),
    .A2(_16841_),
    .ZN(_05324_));
 NAND3_X1 _27679_ (.A1(_03466_),
    .A2(_16834_),
    .A3(_05324_),
    .ZN(_05325_));
 AOI22_X1 _27680_ (.A1(_16618_),
    .A2(_16676_),
    .B1(_16629_),
    .B2(_16741_),
    .ZN(_05326_));
 NOR3_X1 _27681_ (.A1(_16767_),
    .A2(_16637_),
    .A3(_05326_),
    .ZN(_05327_));
 NOR3_X1 _27682_ (.A1(_16847_),
    .A2(_16796_),
    .A3(_16841_),
    .ZN(_05328_));
 NOR2_X1 _27683_ (.A1(_05327_),
    .A2(_05328_),
    .ZN(_05329_));
 OAI21_X1 _27684_ (.A(_16660_),
    .B1(_16845_),
    .B2(_16656_),
    .ZN(_05330_));
 AOI221_X1 _27685_ (.A(_16745_),
    .B1(_16828_),
    .B2(_16656_),
    .C1(_05330_),
    .C2(_16794_),
    .ZN(_05331_));
 NOR2_X2 _27686_ (.A1(_16792_),
    .A2(_16775_),
    .ZN(_05332_));
 OAI21_X1 _27687_ (.A(_16841_),
    .B1(_16737_),
    .B2(_16663_),
    .ZN(_05333_));
 AOI221_X2 _27688_ (.A(_16676_),
    .B1(_16686_),
    .B2(_05332_),
    .C1(_05333_),
    .C2(_16733_),
    .ZN(_05334_));
 OAI221_X1 _27689_ (.A(_05325_),
    .B1(_05329_),
    .B2(_05063_),
    .C1(_05331_),
    .C2(_05334_),
    .ZN(_05335_));
 NAND3_X1 _27690_ (.A1(_16733_),
    .A2(_16638_),
    .A3(_16740_),
    .ZN(_05336_));
 AOI21_X1 _27691_ (.A(_16796_),
    .B1(_16831_),
    .B2(_16794_),
    .ZN(_05337_));
 MUX2_X1 _27692_ (.A(_16630_),
    .B(_16699_),
    .S(_16715_),
    .Z(_05338_));
 AOI21_X1 _27693_ (.A(_05337_),
    .B1(_05338_),
    .B2(_16803_),
    .ZN(_05339_));
 AOI21_X1 _27694_ (.A(_03460_),
    .B1(_05339_),
    .B2(_16834_),
    .ZN(_05340_));
 OAI21_X1 _27695_ (.A(_05336_),
    .B1(_05340_),
    .B2(_16799_),
    .ZN(_05341_));
 NOR3_X1 _27696_ (.A1(_05323_),
    .A2(_05335_),
    .A3(_05341_),
    .ZN(_05342_));
 NAND3_X2 _27697_ (.A1(_05297_),
    .A2(_05309_),
    .A3(_05342_),
    .ZN(_05343_));
 NOR2_X4 _27698_ (.A1(_05291_),
    .A2(_05343_),
    .ZN(_05344_));
 XNOR2_X2 _27699_ (.A(_16978_),
    .B(_03616_),
    .ZN(_05345_));
 XOR2_X1 _27700_ (.A(_17198_),
    .B(_05177_),
    .Z(_05346_));
 XNOR2_X1 _27701_ (.A(_16875_),
    .B(_05346_),
    .ZN(_05347_));
 XNOR2_X2 _27702_ (.A(_05345_),
    .B(_05347_),
    .ZN(_05348_));
 XNOR2_X1 _27703_ (.A(_17185_),
    .B(_03525_),
    .ZN(_05349_));
 XNOR2_X2 _27704_ (.A(_05348_),
    .B(_05349_),
    .ZN(_05350_));
 XNOR2_X1 _27705_ (.A(_17063_),
    .B(_03628_),
    .ZN(_05351_));
 AOI22_X1 _27706_ (.A1(\core.keymem.key_mem[4][91] ),
    .A2(_16457_),
    .B1(_16398_),
    .B2(\core.keymem.key_mem[12][91] ),
    .ZN(_05352_));
 AOI21_X1 _27707_ (.A(_16982_),
    .B1(_16536_),
    .B2(\core.keymem.key_mem[9][91] ),
    .ZN(_05353_));
 AOI22_X1 _27708_ (.A1(\core.keymem.key_mem[6][91] ),
    .A2(_16448_),
    .B1(_16993_),
    .B2(\core.keymem.key_mem[2][91] ),
    .ZN(_05354_));
 AOI22_X1 _27709_ (.A1(\core.keymem.key_mem[10][91] ),
    .A2(_16432_),
    .B1(_16416_),
    .B2(\core.keymem.key_mem[1][91] ),
    .ZN(_05355_));
 AND4_X2 _27710_ (.A1(_05352_),
    .A2(_05353_),
    .A3(_05354_),
    .A4(_05355_),
    .ZN(_05356_));
 AOI222_X2 _27711_ (.A1(\core.keymem.key_mem[7][91] ),
    .A2(_16407_),
    .B1(_17175_),
    .B2(\core.keymem.key_mem[3][91] ),
    .C1(_17007_),
    .C2(\core.keymem.key_mem[11][91] ),
    .ZN(_05357_));
 AOI22_X1 _27712_ (.A1(\core.keymem.key_mem[14][91] ),
    .A2(_16438_),
    .B1(_16472_),
    .B2(\core.keymem.key_mem[13][91] ),
    .ZN(_05358_));
 AOI22_X1 _27713_ (.A1(\core.keymem.key_mem[8][91] ),
    .A2(_16529_),
    .B1(_16949_),
    .B2(\core.keymem.key_mem[5][91] ),
    .ZN(_05359_));
 AND3_X2 _27714_ (.A1(_05357_),
    .A2(_05358_),
    .A3(_05359_),
    .ZN(_05360_));
 AOI22_X4 _27715_ (.A1(_00242_),
    .A2(_16984_),
    .B1(_05356_),
    .B2(_05360_),
    .ZN(_05361_));
 XNOR2_X2 _27716_ (.A(\core.dec_block.block_w1_reg[27] ),
    .B(_05361_),
    .ZN(_05362_));
 XNOR2_X2 _27717_ (.A(_17169_),
    .B(_05362_),
    .ZN(_05363_));
 AND2_X1 _27718_ (.A1(_00245_),
    .A2(_16983_),
    .ZN(_05364_));
 OAI211_X2 _27719_ (.A(\core.keymem.key_mem[7][75] ),
    .B(_17112_),
    .C1(_17107_),
    .C2(_17106_),
    .ZN(_05365_));
 OAI211_X2 _27720_ (.A(\core.keymem.key_mem[10][75] ),
    .B(_17101_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_05366_));
 NAND3_X1 _27721_ (.A1(\core.keymem.key_mem[3][75] ),
    .A2(_17112_),
    .A3(_17121_),
    .ZN(_05367_));
 OAI221_X2 _27722_ (.A(\core.keymem.key_mem[9][75] ),
    .B1(_17103_),
    .B2(_17104_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_05368_));
 NAND4_X2 _27723_ (.A1(_05365_),
    .A2(_05366_),
    .A3(_05367_),
    .A4(_05368_),
    .ZN(_05369_));
 OAI211_X2 _27724_ (.A(\core.keymem.key_mem[13][75] ),
    .B(_17100_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_05370_));
 OAI211_X2 _27725_ (.A(\core.keymem.key_mem[4][75] ),
    .B(_17057_),
    .C1(_17107_),
    .C2(_17106_),
    .ZN(_05371_));
 NAND3_X1 _27726_ (.A1(\core.keymem.key_mem[14][75] ),
    .A2(_17100_),
    .A3(_17050_),
    .ZN(_05372_));
 OAI211_X2 _27727_ (.A(\core.keymem.key_mem[1][75] ),
    .B(_16970_),
    .C1(_17116_),
    .C2(_17118_),
    .ZN(_05373_));
 NAND4_X2 _27728_ (.A1(_05370_),
    .A2(_05371_),
    .A3(_05372_),
    .A4(_05373_),
    .ZN(_05374_));
 OAI211_X2 _27729_ (.A(\core.keymem.key_mem[6][75] ),
    .B(_17050_),
    .C1(_17106_),
    .C2(_17114_),
    .ZN(_05375_));
 OAI211_X2 _27730_ (.A(\core.keymem.key_mem[11][75] ),
    .B(_17048_),
    .C1(_17103_),
    .C2(_17104_),
    .ZN(_05376_));
 OAI221_X2 _27731_ (.A(\core.keymem.key_mem[5][75] ),
    .B1(_17146_),
    .B2(_17622_),
    .C1(_17019_),
    .C2(_17021_),
    .ZN(_05377_));
 NAND3_X1 _27732_ (.A1(\core.keymem.key_mem[2][75] ),
    .A2(_16970_),
    .A3(_17050_),
    .ZN(_05378_));
 NAND4_X2 _27733_ (.A1(_05375_),
    .A2(_05376_),
    .A3(_05377_),
    .A4(_05378_),
    .ZN(_05379_));
 INV_X1 _27734_ (.A(\core.keymem.key_mem[8][75] ),
    .ZN(_05380_));
 INV_X1 _27735_ (.A(\core.keymem.key_mem[12][75] ),
    .ZN(_05381_));
 OAI22_X4 _27736_ (.A1(_05380_),
    .A2(_17134_),
    .B1(_17843_),
    .B2(_05381_),
    .ZN(_05382_));
 NOR4_X4 _27737_ (.A1(_05369_),
    .A2(_05374_),
    .A3(_05379_),
    .A4(_05382_),
    .ZN(_05383_));
 AOI21_X4 _27738_ (.A(_05364_),
    .B1(_05383_),
    .B2(_17533_),
    .ZN(_05384_));
 XNOR2_X2 _27739_ (.A(\core.dec_block.block_w1_reg[11] ),
    .B(_05384_),
    .ZN(_05385_));
 XNOR2_X2 _27740_ (.A(_05115_),
    .B(_05385_),
    .ZN(_05386_));
 XNOR2_X1 _27741_ (.A(_05363_),
    .B(_05386_),
    .ZN(_05387_));
 XNOR2_X1 _27742_ (.A(_05351_),
    .B(_05387_),
    .ZN(_05388_));
 XNOR2_X1 _27743_ (.A(_17141_),
    .B(_05388_),
    .ZN(_05389_));
 XNOR2_X2 _27744_ (.A(_05350_),
    .B(_05389_),
    .ZN(_05390_));
 INV_X1 _27745_ (.A(\core.dec_block.block_w1_reg[2] ),
    .ZN(_05391_));
 XNOR2_X2 _27746_ (.A(_05391_),
    .B(_05033_),
    .ZN(_05392_));
 XNOR2_X2 _27747_ (.A(_17185_),
    .B(_05392_),
    .ZN(_05393_));
 INV_X1 _27748_ (.A(\core.dec_block.block_w1_reg[19] ),
    .ZN(_05394_));
 NAND2_X1 _27749_ (.A1(_00243_),
    .A2(_17183_),
    .ZN(_05395_));
 AOI22_X1 _27750_ (.A1(\core.keymem.key_mem[2][83] ),
    .A2(_16860_),
    .B1(_16515_),
    .B2(\core.keymem.key_mem[10][83] ),
    .ZN(_05396_));
 AOI22_X1 _27751_ (.A1(\core.keymem.key_mem[14][83] ),
    .A2(_16438_),
    .B1(_16448_),
    .B2(\core.keymem.key_mem[6][83] ),
    .ZN(_05397_));
 AOI22_X1 _27752_ (.A1(\core.keymem.key_mem[3][83] ),
    .A2(_16386_),
    .B1(_16416_),
    .B2(\core.keymem.key_mem[1][83] ),
    .ZN(_05398_));
 AOI22_X1 _27753_ (.A1(\core.keymem.key_mem[9][83] ),
    .A2(_16462_),
    .B1(_16472_),
    .B2(\core.keymem.key_mem[13][83] ),
    .ZN(_05399_));
 AND4_X1 _27754_ (.A1(_05396_),
    .A2(_05397_),
    .A3(_05398_),
    .A4(_05399_),
    .ZN(_05400_));
 AOI22_X2 _27755_ (.A1(\core.keymem.key_mem[4][83] ),
    .A2(_16458_),
    .B1(_16507_),
    .B2(\core.keymem.key_mem[11][83] ),
    .ZN(_05401_));
 AOI22_X2 _27756_ (.A1(\core.keymem.key_mem[7][83] ),
    .A2(_16513_),
    .B1(_16469_),
    .B2(\core.keymem.key_mem[5][83] ),
    .ZN(_05402_));
 AOI22_X4 _27757_ (.A1(\core.keymem.key_mem[8][83] ),
    .A2(_16530_),
    .B1(_16540_),
    .B2(\core.keymem.key_mem[12][83] ),
    .ZN(_05403_));
 NAND4_X4 _27758_ (.A1(_05400_),
    .A2(_05401_),
    .A3(_05402_),
    .A4(_05403_),
    .ZN(_05404_));
 OAI21_X4 _27759_ (.A(_05395_),
    .B1(_05404_),
    .B2(_16873_),
    .ZN(_05405_));
 XNOR2_X2 _27760_ (.A(_05394_),
    .B(_05405_),
    .ZN(_05406_));
 XNOR2_X2 _27761_ (.A(_17169_),
    .B(_05138_),
    .ZN(_05407_));
 XOR2_X1 _27762_ (.A(_05406_),
    .B(_05407_),
    .Z(_05408_));
 XNOR2_X1 _27763_ (.A(_05393_),
    .B(_05408_),
    .ZN(_05409_));
 XNOR2_X2 _27764_ (.A(_05390_),
    .B(_05409_),
    .ZN(_05410_));
 OAI21_X1 _27765_ (.A(_05344_),
    .B1(_05410_),
    .B2(_17204_),
    .ZN(_05411_));
 OAI22_X1 _27766_ (.A1(\core.dec_block.block_w0_reg[3] ),
    .A2(_16366_),
    .B1(_05284_),
    .B2(_05411_),
    .ZN(_05412_));
 INV_X1 _27767_ (.A(_05412_),
    .ZN(_00592_));
 NOR3_X1 _27768_ (.A1(_16692_),
    .A2(_16694_),
    .A3(_16742_),
    .ZN(_05413_));
 NOR3_X1 _27769_ (.A1(_16682_),
    .A2(_16631_),
    .A3(_16710_),
    .ZN(_05414_));
 OR3_X2 _27770_ (.A1(_03427_),
    .A2(_05413_),
    .A3(_05414_),
    .ZN(_05415_));
 NAND2_X1 _27771_ (.A1(_16722_),
    .A2(_16789_),
    .ZN(_05416_));
 AOI22_X1 _27772_ (.A1(_16678_),
    .A2(_16760_),
    .B1(_16790_),
    .B2(_16811_),
    .ZN(_05417_));
 OAI221_X1 _27773_ (.A(_05063_),
    .B1(_16803_),
    .B2(_05416_),
    .C1(_05417_),
    .C2(_16655_),
    .ZN(_05418_));
 NOR2_X2 _27774_ (.A1(_16648_),
    .A2(_16675_),
    .ZN(_05419_));
 OAI21_X1 _27775_ (.A(_05419_),
    .B1(_03483_),
    .B2(_16760_),
    .ZN(_05420_));
 NAND2_X1 _27776_ (.A1(_16650_),
    .A2(_16701_),
    .ZN(_05421_));
 NAND2_X1 _27777_ (.A1(_03466_),
    .A2(_16678_),
    .ZN(_05422_));
 NOR3_X1 _27778_ (.A1(_16743_),
    .A2(_16790_),
    .A3(_05058_),
    .ZN(_05423_));
 OAI221_X1 _27779_ (.A(_05420_),
    .B1(_05421_),
    .B2(_03466_),
    .C1(_05422_),
    .C2(_05423_),
    .ZN(_05424_));
 OAI21_X1 _27780_ (.A(_05418_),
    .B1(_05424_),
    .B2(_05063_),
    .ZN(_05425_));
 OAI22_X1 _27781_ (.A1(_16847_),
    .A2(_16732_),
    .B1(_16841_),
    .B2(_16701_),
    .ZN(_05426_));
 AOI22_X1 _27782_ (.A1(_16760_),
    .A2(_16761_),
    .B1(_05426_),
    .B2(_16664_),
    .ZN(_05427_));
 NOR2_X1 _27783_ (.A1(_16655_),
    .A2(_05427_),
    .ZN(_05428_));
 OAI21_X1 _27784_ (.A(_16758_),
    .B1(_16805_),
    .B2(_16659_),
    .ZN(_05429_));
 AOI21_X1 _27785_ (.A(_16701_),
    .B1(_16841_),
    .B2(_16738_),
    .ZN(_05430_));
 OAI21_X1 _27786_ (.A(_16733_),
    .B1(_05328_),
    .B2(_05430_),
    .ZN(_05431_));
 NAND4_X1 _27787_ (.A1(_03487_),
    .A2(_05070_),
    .A3(_05429_),
    .A4(_05431_),
    .ZN(_05432_));
 NOR2_X1 _27788_ (.A1(_16708_),
    .A2(_16763_),
    .ZN(_05433_));
 OAI221_X2 _27789_ (.A(_16794_),
    .B1(_16667_),
    .B2(_05096_),
    .C1(_05433_),
    .C2(_16745_),
    .ZN(_05434_));
 OAI21_X1 _27790_ (.A(_16753_),
    .B1(_16847_),
    .B2(_16725_),
    .ZN(_05435_));
 NAND3_X1 _27791_ (.A1(_16664_),
    .A2(_05434_),
    .A3(_05435_),
    .ZN(_05436_));
 OAI21_X2 _27792_ (.A(_05436_),
    .B1(_16826_),
    .B2(_16685_),
    .ZN(_05437_));
 NOR4_X1 _27793_ (.A1(_03434_),
    .A2(_05428_),
    .A3(_05432_),
    .A4(_05437_),
    .ZN(_05438_));
 AOI22_X1 _27794_ (.A1(_16708_),
    .A2(_16704_),
    .B1(_16761_),
    .B2(_16686_),
    .ZN(_05439_));
 AOI21_X1 _27795_ (.A(_05439_),
    .B1(_16631_),
    .B2(_16663_),
    .ZN(_05440_));
 AOI22_X1 _27796_ (.A1(_16790_),
    .A2(_05069_),
    .B1(_03476_),
    .B2(_16746_),
    .ZN(_05441_));
 NAND3_X1 _27797_ (.A1(_16737_),
    .A2(_03446_),
    .A3(_03470_),
    .ZN(_05442_));
 MUX2_X1 _27798_ (.A(_16680_),
    .B(_16732_),
    .S(_16654_),
    .Z(_05443_));
 OAI221_X1 _27799_ (.A(_05441_),
    .B1(_05442_),
    .B2(_05443_),
    .C1(_16725_),
    .C2(_03397_),
    .ZN(_05444_));
 NOR2_X1 _27800_ (.A1(_16664_),
    .A2(_05052_),
    .ZN(_05445_));
 NOR2_X1 _27801_ (.A1(_16715_),
    .A2(_16761_),
    .ZN(_05446_));
 OAI221_X1 _27802_ (.A(_05446_),
    .B1(_16747_),
    .B2(_16743_),
    .C1(_16754_),
    .C2(_16691_),
    .ZN(_05447_));
 NOR2_X1 _27803_ (.A1(_05445_),
    .A2(_05447_),
    .ZN(_05448_));
 NOR3_X1 _27804_ (.A1(_05440_),
    .A2(_05444_),
    .A3(_05448_),
    .ZN(_05449_));
 OAI21_X1 _27805_ (.A(_16603_),
    .B1(_16704_),
    .B2(_03430_),
    .ZN(_05450_));
 OAI21_X2 _27806_ (.A(_05450_),
    .B1(_16823_),
    .B2(_16682_),
    .ZN(_05451_));
 NOR3_X2 _27807_ (.A1(_16753_),
    .A2(_16727_),
    .A3(_03382_),
    .ZN(_05452_));
 NOR3_X2 _27808_ (.A1(_16794_),
    .A2(_16793_),
    .A3(_16647_),
    .ZN(_05453_));
 OAI21_X1 _27809_ (.A(_16764_),
    .B1(_16685_),
    .B2(_16775_),
    .ZN(_05454_));
 OAI21_X1 _27810_ (.A(_05454_),
    .B1(_16716_),
    .B2(_16764_),
    .ZN(_05455_));
 AOI21_X2 _27811_ (.A(_16785_),
    .B1(_05045_),
    .B2(_05455_),
    .ZN(_05456_));
 NOR4_X4 _27812_ (.A1(_05451_),
    .A2(_05452_),
    .A3(_05453_),
    .A4(_05456_),
    .ZN(_05457_));
 NAND2_X1 _27813_ (.A1(_16698_),
    .A2(_16689_),
    .ZN(_05458_));
 NAND2_X1 _27814_ (.A1(_16675_),
    .A2(_05458_),
    .ZN(_05459_));
 OAI21_X1 _27815_ (.A(_16635_),
    .B1(_16659_),
    .B2(_05459_),
    .ZN(_05460_));
 NAND2_X1 _27816_ (.A1(_16659_),
    .A2(_16691_),
    .ZN(_05461_));
 NOR2_X1 _27817_ (.A1(_16625_),
    .A2(_16747_),
    .ZN(_05462_));
 OAI21_X1 _27818_ (.A(_16722_),
    .B1(_16675_),
    .B2(_16790_),
    .ZN(_05463_));
 AOI221_X2 _27819_ (.A(_05460_),
    .B1(_05461_),
    .B2(_05462_),
    .C1(_05463_),
    .C2(_16634_),
    .ZN(_05464_));
 NOR3_X1 _27820_ (.A1(_16656_),
    .A2(_16728_),
    .A3(_05446_),
    .ZN(_05465_));
 OAI222_X2 _27821_ (.A1(_16631_),
    .A2(_03479_),
    .B1(_16781_),
    .B2(_16738_),
    .C1(_16845_),
    .C2(_16759_),
    .ZN(_05466_));
 NOR4_X1 _27822_ (.A1(_16778_),
    .A2(_05464_),
    .A3(_05465_),
    .A4(_05466_),
    .ZN(_05467_));
 NAND3_X1 _27823_ (.A1(_05449_),
    .A2(_05457_),
    .A3(_05467_),
    .ZN(_05468_));
 NAND3_X1 _27824_ (.A1(_03466_),
    .A2(_16822_),
    .A3(_16678_),
    .ZN(_05469_));
 AOI21_X1 _27825_ (.A(_16750_),
    .B1(_16746_),
    .B2(_16847_),
    .ZN(_05470_));
 OAI21_X1 _27826_ (.A(_16718_),
    .B1(_05470_),
    .B2(_16753_),
    .ZN(_05471_));
 AOI22_X1 _27827_ (.A1(_16673_),
    .A2(_16782_),
    .B1(_05471_),
    .B2(_16834_),
    .ZN(_05472_));
 OAI21_X1 _27828_ (.A(_05469_),
    .B1(_05472_),
    .B2(_16678_),
    .ZN(_05473_));
 NOR3_X1 _27829_ (.A1(_05341_),
    .A2(_05468_),
    .A3(_05473_),
    .ZN(_05474_));
 NAND3_X1 _27830_ (.A1(_05425_),
    .A2(_05438_),
    .A3(_05474_),
    .ZN(_05475_));
 NOR2_X2 _27831_ (.A1(_05415_),
    .A2(_05475_),
    .ZN(_05476_));
 NOR2_X2 _27832_ (.A1(_17379_),
    .A2(_05476_),
    .ZN(_05477_));
 NAND2_X1 _27833_ (.A1(_00249_),
    .A2(_17578_),
    .ZN(_05478_));
 AOI222_X2 _27834_ (.A1(\core.keymem.key_mem[4][68] ),
    .A2(_16501_),
    .B1(_17585_),
    .B2(\core.keymem.key_mem[9][68] ),
    .C1(\core.keymem.key_mem[11][68] ),
    .C2(_17769_),
    .ZN(_05479_));
 AOI22_X2 _27835_ (.A1(\core.keymem.key_mem[8][68] ),
    .A2(_17765_),
    .B1(_17082_),
    .B2(\core.keymem.key_mem[10][68] ),
    .ZN(_05480_));
 AOI22_X2 _27836_ (.A1(\core.keymem.key_mem[7][68] ),
    .A2(_17085_),
    .B1(_17086_),
    .B2(\core.keymem.key_mem[2][68] ),
    .ZN(_05481_));
 NAND3_X2 _27837_ (.A1(_05479_),
    .A2(_05480_),
    .A3(_05481_),
    .ZN(_05482_));
 AOI21_X1 _27838_ (.A(_16984_),
    .B1(_16526_),
    .B2(\core.keymem.key_mem[1][68] ),
    .ZN(_05483_));
 AOI22_X2 _27839_ (.A1(\core.keymem.key_mem[6][68] ),
    .A2(_16522_),
    .B1(_17091_),
    .B2(\core.keymem.key_mem[3][68] ),
    .ZN(_05484_));
 AOI22_X2 _27840_ (.A1(\core.keymem.key_mem[14][68] ),
    .A2(_17581_),
    .B1(_16510_),
    .B2(\core.keymem.key_mem[5][68] ),
    .ZN(_05485_));
 AOI22_X2 _27841_ (.A1(\core.keymem.key_mem[12][68] ),
    .A2(_17093_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][68] ),
    .ZN(_05486_));
 NAND4_X2 _27842_ (.A1(_05483_),
    .A2(_05484_),
    .A3(_05485_),
    .A4(_05486_),
    .ZN(_05487_));
 OAI21_X4 _27843_ (.A(_05478_),
    .B1(_05482_),
    .B2(_05487_),
    .ZN(_05488_));
 XNOR2_X1 _27844_ (.A(\block_reg[1][4] ),
    .B(_05488_),
    .ZN(_05489_));
 AOI21_X1 _27845_ (.A(_16367_),
    .B1(_16371_),
    .B2(_05489_),
    .ZN(_05490_));
 XNOR2_X2 _27846_ (.A(_17079_),
    .B(_03541_),
    .ZN(_05491_));
 XNOR2_X2 _27847_ (.A(_16943_),
    .B(_03556_),
    .ZN(_05492_));
 XNOR2_X2 _27848_ (.A(_05491_),
    .B(_05492_),
    .ZN(_05493_));
 XOR2_X2 _27849_ (.A(_03597_),
    .B(_05493_),
    .Z(_05494_));
 XNOR2_X1 _27850_ (.A(_03627_),
    .B(_05392_),
    .ZN(_05495_));
 XNOR2_X1 _27851_ (.A(_03616_),
    .B(_05178_),
    .ZN(_05496_));
 XNOR2_X1 _27852_ (.A(_05495_),
    .B(_05496_),
    .ZN(_05497_));
 XNOR2_X2 _27853_ (.A(_05494_),
    .B(_05497_),
    .ZN(_05498_));
 AOI222_X2 _27854_ (.A1(\core.keymem.key_mem[14][92] ),
    .A2(_16502_),
    .B1(_16425_),
    .B2(\core.keymem.key_mem[2][92] ),
    .C1(_16417_),
    .C2(\core.keymem.key_mem[1][92] ),
    .ZN(_05499_));
 AOI22_X1 _27855_ (.A1(\core.keymem.key_mem[10][92] ),
    .A2(_16516_),
    .B1(_16533_),
    .B2(\core.keymem.key_mem[13][92] ),
    .ZN(_05500_));
 AOI22_X1 _27856_ (.A1(\core.keymem.key_mem[3][92] ),
    .A2(_17091_),
    .B1(_17093_),
    .B2(\core.keymem.key_mem[12][92] ),
    .ZN(_05501_));
 NAND3_X1 _27857_ (.A1(_05499_),
    .A2(_05500_),
    .A3(_05501_),
    .ZN(_05502_));
 AOI22_X1 _27858_ (.A1(\core.keymem.key_mem[6][92] ),
    .A2(_16449_),
    .B1(_16507_),
    .B2(\core.keymem.key_mem[11][92] ),
    .ZN(_05503_));
 AOI22_X1 _27859_ (.A1(\core.keymem.key_mem[7][92] ),
    .A2(_17085_),
    .B1(_16530_),
    .B2(\core.keymem.key_mem[8][92] ),
    .ZN(_05504_));
 AOI22_X1 _27860_ (.A1(\core.keymem.key_mem[9][92] ),
    .A2(_16537_),
    .B1(_16469_),
    .B2(\core.keymem.key_mem[5][92] ),
    .ZN(_05505_));
 AOI21_X1 _27861_ (.A(_16496_),
    .B1(_16458_),
    .B2(\core.keymem.key_mem[4][92] ),
    .ZN(_05506_));
 NAND4_X1 _27862_ (.A1(_05503_),
    .A2(_05504_),
    .A3(_05505_),
    .A4(_05506_),
    .ZN(_05507_));
 NOR2_X2 _27863_ (.A1(_05502_),
    .A2(_05507_),
    .ZN(_05508_));
 AOI21_X4 _27864_ (.A(_05508_),
    .B1(_17578_),
    .B2(_00247_),
    .ZN(_05509_));
 XNOR2_X2 _27865_ (.A(\core.dec_block.block_w1_reg[28] ),
    .B(_05509_),
    .ZN(_05510_));
 XNOR2_X1 _27866_ (.A(_05363_),
    .B(_05510_),
    .ZN(_05511_));
 XNOR2_X2 _27867_ (.A(_17199_),
    .B(_05511_),
    .ZN(_05512_));
 AOI222_X2 _27868_ (.A1(\core.keymem.key_mem[8][84] ),
    .A2(_17666_),
    .B1(_16509_),
    .B2(\core.keymem.key_mem[5][84] ),
    .C1(_16442_),
    .C2(\core.keymem.key_mem[11][84] ),
    .ZN(_05513_));
 AOI22_X1 _27869_ (.A1(\core.keymem.key_mem[4][84] ),
    .A2(_18232_),
    .B1(_16999_),
    .B2(\core.keymem.key_mem[14][84] ),
    .ZN(_05514_));
 AOI22_X1 _27870_ (.A1(\core.keymem.key_mem[3][84] ),
    .A2(_17683_),
    .B1(_17001_),
    .B2(\core.keymem.key_mem[12][84] ),
    .ZN(_05515_));
 NAND3_X1 _27871_ (.A1(_05513_),
    .A2(_05514_),
    .A3(_05515_),
    .ZN(_05516_));
 AOI22_X1 _27872_ (.A1(\core.keymem.key_mem[7][84] ),
    .A2(_17789_),
    .B1(_16521_),
    .B2(\core.keymem.key_mem[6][84] ),
    .ZN(_05517_));
 AOI22_X1 _27873_ (.A1(\core.keymem.key_mem[10][84] ),
    .A2(_16989_),
    .B1(_17784_),
    .B2(\core.keymem.key_mem[13][84] ),
    .ZN(_05518_));
 AOI22_X1 _27874_ (.A1(\core.keymem.key_mem[2][84] ),
    .A2(_17786_),
    .B1(_16525_),
    .B2(\core.keymem.key_mem[1][84] ),
    .ZN(_05519_));
 AOI21_X1 _27875_ (.A(_17013_),
    .B1(_17914_),
    .B2(\core.keymem.key_mem[9][84] ),
    .ZN(_05520_));
 NAND4_X1 _27876_ (.A1(_05517_),
    .A2(_05518_),
    .A3(_05519_),
    .A4(_05520_),
    .ZN(_05521_));
 NOR2_X2 _27877_ (.A1(_05516_),
    .A2(_05521_),
    .ZN(_05522_));
 AOI21_X4 _27878_ (.A(_05522_),
    .B1(_16548_),
    .B2(_00248_),
    .ZN(_05523_));
 XNOR2_X2 _27879_ (.A(\core.dec_block.block_w1_reg[20] ),
    .B(_05523_),
    .ZN(_05524_));
 INV_X1 _27880_ (.A(\core.dec_block.block_w1_reg[12] ),
    .ZN(_05525_));
 NAND2_X1 _27881_ (.A1(_00250_),
    .A2(_16549_),
    .ZN(_05526_));
 AOI22_X1 _27882_ (.A1(\core.keymem.key_mem[10][76] ),
    .A2(_16516_),
    .B1(_16469_),
    .B2(\core.keymem.key_mem[5][76] ),
    .ZN(_05527_));
 AOI22_X1 _27883_ (.A1(\core.keymem.key_mem[7][76] ),
    .A2(_16513_),
    .B1(_17178_),
    .B2(\core.keymem.key_mem[1][76] ),
    .ZN(_05528_));
 AOI22_X1 _27884_ (.A1(\core.keymem.key_mem[14][76] ),
    .A2(_16502_),
    .B1(_16449_),
    .B2(\core.keymem.key_mem[6][76] ),
    .ZN(_05529_));
 AOI22_X1 _27885_ (.A1(\core.keymem.key_mem[2][76] ),
    .A2(_16425_),
    .B1(_16540_),
    .B2(\core.keymem.key_mem[12][76] ),
    .ZN(_05530_));
 AND4_X1 _27886_ (.A1(_05527_),
    .A2(_05528_),
    .A3(_05529_),
    .A4(_05530_),
    .ZN(_05531_));
 AOI22_X2 _27887_ (.A1(\core.keymem.key_mem[4][76] ),
    .A2(_16501_),
    .B1(_17765_),
    .B2(\core.keymem.key_mem[8][76] ),
    .ZN(_05532_));
 AOI22_X2 _27888_ (.A1(\core.keymem.key_mem[9][76] ),
    .A2(_17585_),
    .B1(_17771_),
    .B2(\core.keymem.key_mem[13][76] ),
    .ZN(_05533_));
 AOI22_X2 _27889_ (.A1(\core.keymem.key_mem[3][76] ),
    .A2(_17091_),
    .B1(_17769_),
    .B2(\core.keymem.key_mem[11][76] ),
    .ZN(_05534_));
 NAND4_X2 _27890_ (.A1(_05531_),
    .A2(_05532_),
    .A3(_05533_),
    .A4(_05534_),
    .ZN(_05535_));
 OAI21_X4 _27891_ (.A(_05526_),
    .B1(_05535_),
    .B2(_16549_),
    .ZN(_05536_));
 XNOR2_X2 _27892_ (.A(_05525_),
    .B(_05536_),
    .ZN(_05537_));
 XNOR2_X2 _27893_ (.A(_05524_),
    .B(_05537_),
    .ZN(_05538_));
 XNOR2_X2 _27894_ (.A(\core.dec_block.block_w1_reg[3] ),
    .B(_05282_),
    .ZN(_05539_));
 XNOR2_X2 _27895_ (.A(_17185_),
    .B(_05539_),
    .ZN(_05540_));
 XOR2_X1 _27896_ (.A(_05538_),
    .B(_05540_),
    .Z(_05541_));
 XNOR2_X1 _27897_ (.A(_05512_),
    .B(_05541_),
    .ZN(_05542_));
 XNOR2_X1 _27898_ (.A(_05498_),
    .B(_05542_),
    .ZN(_05543_));
 OAI221_X1 _27899_ (.A(_05490_),
    .B1(_05543_),
    .B2(_17203_),
    .C1(_05021_),
    .C2(_04937_),
    .ZN(_05544_));
 NOR2_X1 _27900_ (.A1(_05477_),
    .A2(_05544_),
    .ZN(_05545_));
 AOI21_X1 _27901_ (.A(_05545_),
    .B1(_17744_),
    .B2(_04925_),
    .ZN(_00593_));
 XNOR2_X1 _27902_ (.A(\block_reg[1][5] ),
    .B(_17197_),
    .ZN(_05546_));
 OAI221_X1 _27903_ (.A(_16365_),
    .B1(_03858_),
    .B2(_04365_),
    .C1(_05546_),
    .C2(_04266_),
    .ZN(_05547_));
 OAI22_X1 _27904_ (.A1(_16676_),
    .A2(_16728_),
    .B1(_16846_),
    .B2(_16793_),
    .ZN(_05548_));
 NOR2_X1 _27905_ (.A1(_16648_),
    .A2(_16740_),
    .ZN(_05549_));
 AOI22_X1 _27906_ (.A1(_16799_),
    .A2(_05548_),
    .B1(_05549_),
    .B2(_16828_),
    .ZN(_05550_));
 OR2_X1 _27907_ (.A1(_05063_),
    .A2(_05550_),
    .ZN(_05551_));
 NOR2_X1 _27908_ (.A1(_16717_),
    .A2(_16747_),
    .ZN(_05552_));
 OAI221_X1 _27909_ (.A(_16672_),
    .B1(_16691_),
    .B2(_16845_),
    .C1(_03366_),
    .C2(_05552_),
    .ZN(_05553_));
 NAND3_X1 _27910_ (.A1(_16655_),
    .A2(_05063_),
    .A3(_05553_),
    .ZN(_05554_));
 NAND2_X1 _27911_ (.A1(_16698_),
    .A2(_16669_),
    .ZN(_05555_));
 AOI21_X1 _27912_ (.A(_16609_),
    .B1(_03446_),
    .B2(_05555_),
    .ZN(_05556_));
 NOR3_X1 _27913_ (.A1(_16698_),
    .A2(_16669_),
    .A3(_16649_),
    .ZN(_05557_));
 OR2_X1 _27914_ (.A1(_05556_),
    .A2(_05557_),
    .ZN(_05558_));
 AOI221_X2 _27915_ (.A(_16715_),
    .B1(_16698_),
    .B2(_16650_),
    .C1(_05558_),
    .C2(_16808_),
    .ZN(_05559_));
 AOI22_X1 _27916_ (.A1(_16664_),
    .A2(_16659_),
    .B1(_16765_),
    .B2(_16747_),
    .ZN(_05560_));
 AOI21_X1 _27917_ (.A(_05559_),
    .B1(_05560_),
    .B2(_16767_),
    .ZN(_05561_));
 OAI21_X1 _27918_ (.A(_16799_),
    .B1(_05076_),
    .B2(_05561_),
    .ZN(_05562_));
 OAI33_X1 _27919_ (.A1(_16654_),
    .A2(_16705_),
    .A3(_16684_),
    .B1(_05549_),
    .B2(_16612_),
    .B3(_16649_),
    .ZN(_05563_));
 AOI22_X2 _27920_ (.A1(_16825_),
    .A2(_16695_),
    .B1(_05563_),
    .B2(_16656_),
    .ZN(_05564_));
 NOR3_X1 _27921_ (.A1(_16775_),
    .A2(_16764_),
    .A3(_05316_),
    .ZN(_05565_));
 AOI21_X1 _27922_ (.A(_05565_),
    .B1(_16750_),
    .B2(_16676_),
    .ZN(_05566_));
 OAI21_X1 _27923_ (.A(_05564_),
    .B1(_05566_),
    .B2(_16736_),
    .ZN(_05567_));
 OAI22_X2 _27924_ (.A1(_16647_),
    .A2(_16725_),
    .B1(_05416_),
    .B2(_16764_),
    .ZN(_05568_));
 OAI22_X1 _27925_ (.A1(_16698_),
    .A2(_16725_),
    .B1(_05458_),
    .B2(_16685_),
    .ZN(_05569_));
 AOI22_X2 _27926_ (.A1(_16733_),
    .A2(_05568_),
    .B1(_05569_),
    .B2(_05419_),
    .ZN(_05570_));
 NAND2_X1 _27927_ (.A1(_16662_),
    .A2(_16630_),
    .ZN(_05571_));
 AOI21_X1 _27928_ (.A(_05571_),
    .B1(_16831_),
    .B2(_03366_),
    .ZN(_05572_));
 MUX2_X1 _27929_ (.A(_16630_),
    .B(_05316_),
    .S(_16764_),
    .Z(_05573_));
 OAI221_X2 _27930_ (.A(_05570_),
    .B1(_05572_),
    .B2(_16785_),
    .C1(_05573_),
    .C2(_16736_),
    .ZN(_05574_));
 NOR4_X2 _27931_ (.A1(_16768_),
    .A2(_05050_),
    .A3(_05567_),
    .A4(_05574_),
    .ZN(_05575_));
 NAND4_X2 _27932_ (.A1(_05551_),
    .A2(_05554_),
    .A3(_05562_),
    .A4(_05575_),
    .ZN(_05576_));
 AOI22_X1 _27933_ (.A1(_16726_),
    .A2(_16831_),
    .B1(_03488_),
    .B2(_05458_),
    .ZN(_05577_));
 OAI21_X1 _27934_ (.A(_03457_),
    .B1(_05577_),
    .B2(_16655_),
    .ZN(_05578_));
 AOI22_X4 _27935_ (.A1(_16828_),
    .A2(_16704_),
    .B1(_05332_),
    .B2(_16733_),
    .ZN(_05579_));
 AOI21_X2 _27936_ (.A(_16743_),
    .B1(_03449_),
    .B2(_16603_),
    .ZN(_05580_));
 OR2_X1 _27937_ (.A1(_16733_),
    .A2(_16758_),
    .ZN(_05581_));
 AOI22_X1 _27938_ (.A1(_16758_),
    .A2(_05571_),
    .B1(_05581_),
    .B2(_16712_),
    .ZN(_05582_));
 OAI221_X2 _27939_ (.A(_05579_),
    .B1(_05580_),
    .B2(_03470_),
    .C1(_05582_),
    .C2(_16799_),
    .ZN(_05583_));
 NOR2_X1 _27940_ (.A1(_05578_),
    .A2(_05583_),
    .ZN(_05584_));
 AOI22_X1 _27941_ (.A1(_16834_),
    .A2(_16661_),
    .B1(_16686_),
    .B2(_16821_),
    .ZN(_05585_));
 NOR3_X1 _27942_ (.A1(_16612_),
    .A2(_16647_),
    .A3(_05585_),
    .ZN(_05586_));
 AOI21_X1 _27943_ (.A(_05586_),
    .B1(_05324_),
    .B2(_05063_),
    .ZN(_05587_));
 NAND3_X1 _27944_ (.A1(_16829_),
    .A2(_05584_),
    .A3(_05587_),
    .ZN(_05588_));
 NOR4_X4 _27945_ (.A1(_05304_),
    .A2(_05437_),
    .A3(_05576_),
    .A4(_05588_),
    .ZN(_05589_));
 XOR2_X2 _27946_ (.A(\core.dec_block.block_w1_reg[4] ),
    .B(_05488_),
    .Z(_05590_));
 XNOR2_X2 _27947_ (.A(_16875_),
    .B(_05590_),
    .ZN(_05591_));
 XNOR2_X2 _27948_ (.A(_03627_),
    .B(_05176_),
    .ZN(_05592_));
 XOR2_X2 _27949_ (.A(_16979_),
    .B(_05592_),
    .Z(_05593_));
 XNOR2_X2 _27950_ (.A(_05161_),
    .B(_05593_),
    .ZN(_05594_));
 XNOR2_X2 _27951_ (.A(_05591_),
    .B(_05594_),
    .ZN(_05595_));
 XNOR2_X2 _27952_ (.A(_03627_),
    .B(_05406_),
    .ZN(_05596_));
 XNOR2_X2 _27953_ (.A(_05510_),
    .B(_05596_),
    .ZN(_05597_));
 XNOR2_X2 _27954_ (.A(_17062_),
    .B(_17079_),
    .ZN(_05598_));
 XOR2_X1 _27955_ (.A(_05392_),
    .B(_05539_),
    .Z(_05599_));
 XNOR2_X1 _27956_ (.A(_05598_),
    .B(_05599_),
    .ZN(_05600_));
 XNOR2_X1 _27957_ (.A(_05597_),
    .B(_05600_),
    .ZN(_05601_));
 XNOR2_X2 _27958_ (.A(_05595_),
    .B(_05601_),
    .ZN(_05602_));
 OAI21_X1 _27959_ (.A(_05589_),
    .B1(_05602_),
    .B2(_17204_),
    .ZN(_05603_));
 OAI22_X1 _27960_ (.A1(\core.dec_block.block_w0_reg[5] ),
    .A2(_16366_),
    .B1(_05547_),
    .B2(_05603_),
    .ZN(_05604_));
 INV_X1 _27961_ (.A(_05604_),
    .ZN(_00594_));
 NOR2_X1 _27962_ (.A1(\core.dec_block.block_w0_reg[6] ),
    .A2(_16365_),
    .ZN(_05605_));
 XNOR2_X2 _27963_ (.A(\block_reg[1][6] ),
    .B(_16874_),
    .ZN(_05606_));
 OAI221_X1 _27964_ (.A(_18329_),
    .B1(_18052_),
    .B2(_04589_),
    .C1(_05606_),
    .C2(_04266_),
    .ZN(_05607_));
 XNOR2_X2 _27965_ (.A(_05524_),
    .B(_05590_),
    .ZN(_05608_));
 XNOR2_X1 _27966_ (.A(_05491_),
    .B(_05608_),
    .ZN(_05609_));
 XOR2_X1 _27967_ (.A(_05385_),
    .B(_05539_),
    .Z(_05610_));
 XNOR2_X1 _27968_ (.A(_16978_),
    .B(_05610_),
    .ZN(_05611_));
 XNOR2_X1 _27969_ (.A(_05609_),
    .B(_05611_),
    .ZN(_05612_));
 XNOR2_X2 _27970_ (.A(_17199_),
    .B(_05116_),
    .ZN(_05613_));
 XNOR2_X2 _27971_ (.A(_05363_),
    .B(_05596_),
    .ZN(_05614_));
 XNOR2_X1 _27972_ (.A(_05613_),
    .B(_05614_),
    .ZN(_05615_));
 XNOR2_X2 _27973_ (.A(_05612_),
    .B(_05615_),
    .ZN(_05616_));
 AOI21_X1 _27974_ (.A(_05607_),
    .B1(_05616_),
    .B2(_04370_),
    .ZN(_05617_));
 NAND3_X1 _27975_ (.A1(_16839_),
    .A2(_16843_),
    .A3(_16849_),
    .ZN(_05618_));
 INV_X1 _27976_ (.A(_05567_),
    .ZN(_05619_));
 OAI22_X1 _27977_ (.A1(_16634_),
    .A2(_16694_),
    .B1(_16725_),
    .B2(_16726_),
    .ZN(_05620_));
 AOI221_X2 _27978_ (.A(_16737_),
    .B1(_16686_),
    .B2(_03488_),
    .C1(_05620_),
    .C2(_16794_),
    .ZN(_05621_));
 NAND3_X1 _27979_ (.A1(_16654_),
    .A2(_16705_),
    .A3(_16743_),
    .ZN(_05622_));
 NAND3_X1 _27980_ (.A1(_16715_),
    .A2(_16764_),
    .A3(_16790_),
    .ZN(_05623_));
 NAND2_X1 _27981_ (.A1(_05622_),
    .A2(_05623_),
    .ZN(_05624_));
 AOI221_X1 _27982_ (.A(_16667_),
    .B1(_16603_),
    .B2(_16706_),
    .C1(_05624_),
    .C2(_16754_),
    .ZN(_05625_));
 OAI21_X1 _27983_ (.A(_05619_),
    .B1(_05621_),
    .B2(_05625_),
    .ZN(_05626_));
 OAI21_X1 _27984_ (.A(_05419_),
    .B1(_16763_),
    .B2(_16712_),
    .ZN(_05627_));
 NOR2_X1 _27985_ (.A1(_16654_),
    .A2(_16705_),
    .ZN(_05628_));
 AOI21_X1 _27986_ (.A(_05628_),
    .B1(_16741_),
    .B2(_16794_),
    .ZN(_05629_));
 OAI21_X1 _27987_ (.A(_05627_),
    .B1(_05629_),
    .B2(_16738_),
    .ZN(_05630_));
 NAND2_X1 _27988_ (.A1(_16834_),
    .A2(_05630_),
    .ZN(_05631_));
 AOI22_X1 _27989_ (.A1(_16626_),
    .A2(_16716_),
    .B1(_16828_),
    .B2(_16758_),
    .ZN(_05632_));
 OAI21_X1 _27990_ (.A(_16730_),
    .B1(_05632_),
    .B2(_16847_),
    .ZN(_05633_));
 OAI21_X1 _27991_ (.A(_16822_),
    .B1(_16782_),
    .B2(_03476_),
    .ZN(_05634_));
 OAI221_X1 _27992_ (.A(_05634_),
    .B1(_16845_),
    .B2(_03386_),
    .C1(_16793_),
    .C2(_03479_),
    .ZN(_05635_));
 NOR3_X1 _27993_ (.A1(_16787_),
    .A2(_05633_),
    .A3(_05635_),
    .ZN(_05636_));
 NAND4_X1 _27994_ (.A1(_05091_),
    .A2(_05295_),
    .A3(_05631_),
    .A4(_05636_),
    .ZN(_05637_));
 OR4_X2 _27995_ (.A1(_05618_),
    .A2(_03485_),
    .A3(_05626_),
    .A4(_05637_),
    .ZN(_05638_));
 AOI221_X1 _27996_ (.A(_16805_),
    .B1(_16723_),
    .B2(_16712_),
    .C1(_16794_),
    .C2(_16747_),
    .ZN(_05639_));
 OAI221_X1 _27997_ (.A(_16678_),
    .B1(_16841_),
    .B2(_16736_),
    .C1(_05639_),
    .C2(_05063_),
    .ZN(_05640_));
 NAND4_X1 _27998_ (.A1(_16655_),
    .A2(_16664_),
    .A3(_16811_),
    .A4(_16712_),
    .ZN(_05641_));
 OAI21_X1 _27999_ (.A(_05641_),
    .B1(_16840_),
    .B2(_16714_),
    .ZN(_05642_));
 OAI21_X1 _28000_ (.A(_05640_),
    .B1(_05642_),
    .B2(_16678_),
    .ZN(_05643_));
 NOR2_X1 _28001_ (.A1(_16708_),
    .A2(_16743_),
    .ZN(_05644_));
 NAND2_X1 _28002_ (.A1(_16775_),
    .A2(_16746_),
    .ZN(_05645_));
 OAI221_X1 _28003_ (.A(_05645_),
    .B1(_16680_),
    .B2(_16799_),
    .C1(_16602_),
    .C2(_16707_),
    .ZN(_05646_));
 AOI21_X1 _28004_ (.A(_05324_),
    .B1(_05646_),
    .B2(_16678_),
    .ZN(_05647_));
 OAI221_X2 _28005_ (.A(_05643_),
    .B1(_05644_),
    .B2(_03479_),
    .C1(_05647_),
    .C2(_16736_),
    .ZN(_05648_));
 NOR4_X4 _28006_ (.A1(_03379_),
    .A2(_05415_),
    .A3(_05638_),
    .A4(_05648_),
    .ZN(_05649_));
 OR2_X2 _28007_ (.A1(_17379_),
    .A2(_05649_),
    .ZN(_05650_));
 AOI21_X1 _28008_ (.A(_05605_),
    .B1(_05617_),
    .B2(_05650_),
    .ZN(_00595_));
 NOR2_X1 _28009_ (.A1(_16581_),
    .A2(_16365_),
    .ZN(_05651_));
 NOR3_X1 _28010_ (.A1(_16798_),
    .A2(_16745_),
    .A3(_16845_),
    .ZN(_05652_));
 OAI21_X1 _28011_ (.A(_16767_),
    .B1(_16847_),
    .B2(_16685_),
    .ZN(_05653_));
 OAI22_X1 _28012_ (.A1(_03466_),
    .A2(_05324_),
    .B1(_05652_),
    .B2(_05653_),
    .ZN(_05654_));
 NOR3_X1 _28013_ (.A1(_16753_),
    .A2(_16808_),
    .A3(_16770_),
    .ZN(_05655_));
 OAI21_X1 _28014_ (.A(_16670_),
    .B1(_16701_),
    .B2(_16657_),
    .ZN(_05656_));
 AOI22_X1 _28015_ (.A1(_16767_),
    .A2(_03402_),
    .B1(_05655_),
    .B2(_05656_),
    .ZN(_05657_));
 MUX2_X1 _28016_ (.A(_05654_),
    .B(_05657_),
    .S(_05063_),
    .Z(_05658_));
 AOI22_X2 _28017_ (.A1(_16677_),
    .A2(_16831_),
    .B1(_05419_),
    .B2(_16659_),
    .ZN(_05659_));
 OAI221_X2 _28018_ (.A(_05579_),
    .B1(_05580_),
    .B2(_03470_),
    .C1(_05659_),
    .C2(_16834_),
    .ZN(_05660_));
 NOR2_X1 _28019_ (.A1(_16648_),
    .A2(_16705_),
    .ZN(_05661_));
 OAI21_X1 _28020_ (.A(_16634_),
    .B1(_05661_),
    .B2(_03447_),
    .ZN(_05662_));
 OAI22_X1 _28021_ (.A1(_16731_),
    .A2(_05039_),
    .B1(_05645_),
    .B2(_05662_),
    .ZN(_05663_));
 AOI21_X1 _28022_ (.A(_05663_),
    .B1(_16704_),
    .B2(_16717_),
    .ZN(_05664_));
 NOR3_X1 _28023_ (.A1(_16754_),
    .A2(_16667_),
    .A3(_05628_),
    .ZN(_05665_));
 AOI21_X1 _28024_ (.A(_05665_),
    .B1(_16701_),
    .B2(_16666_),
    .ZN(_05666_));
 AOI22_X2 _28025_ (.A1(_16733_),
    .A2(_16717_),
    .B1(_16603_),
    .B2(_16758_),
    .ZN(_05667_));
 OAI221_X2 _28026_ (.A(_05664_),
    .B1(_05666_),
    .B2(_03382_),
    .C1(_16799_),
    .C2(_05667_),
    .ZN(_05668_));
 NOR2_X1 _28027_ (.A1(_16676_),
    .A2(_05645_),
    .ZN(_05669_));
 AOI21_X1 _28028_ (.A(_05669_),
    .B1(_05058_),
    .B2(_16677_),
    .ZN(_05670_));
 NOR2_X1 _28029_ (.A1(_16736_),
    .A2(_05670_),
    .ZN(_05671_));
 NOR4_X2 _28030_ (.A1(_03391_),
    .A2(_05660_),
    .A3(_05668_),
    .A4(_05671_),
    .ZN(_05672_));
 NAND4_X2 _28031_ (.A1(_16837_),
    .A2(_05457_),
    .A3(_05658_),
    .A4(_05672_),
    .ZN(_05673_));
 NOR4_X4 _28032_ (.A1(_05099_),
    .A2(_05291_),
    .A3(_05648_),
    .A4(_05673_),
    .ZN(_05674_));
 INV_X1 _28033_ (.A(\block_reg[1][7] ),
    .ZN(_05675_));
 XNOR2_X1 _28034_ (.A(_05675_),
    .B(_17184_),
    .ZN(_05676_));
 OAI221_X1 _28035_ (.A(_16364_),
    .B1(_17741_),
    .B2(_04723_),
    .C1(_05676_),
    .C2(_18553_),
    .ZN(_05677_));
 XNOR2_X1 _28036_ (.A(_05115_),
    .B(_05510_),
    .ZN(_05678_));
 XNOR2_X1 _28037_ (.A(_05538_),
    .B(_05678_),
    .ZN(_05679_));
 XOR2_X1 _28038_ (.A(_17198_),
    .B(_05591_),
    .Z(_05680_));
 XNOR2_X1 _28039_ (.A(_03542_),
    .B(_03628_),
    .ZN(_05681_));
 XNOR2_X1 _28040_ (.A(_05680_),
    .B(_05681_),
    .ZN(_05682_));
 XNOR2_X1 _28041_ (.A(_05679_),
    .B(_05682_),
    .ZN(_05683_));
 AOI21_X1 _28042_ (.A(_05677_),
    .B1(_05683_),
    .B2(_19031_),
    .ZN(_05684_));
 AOI21_X1 _28043_ (.A(_05651_),
    .B1(_05674_),
    .B2(_05684_),
    .ZN(_00596_));
 NOR2_X1 _28044_ (.A1(\core.dec_block.block_w0_reg[8] ),
    .A2(_16365_),
    .ZN(_05685_));
 AOI21_X1 _28045_ (.A(_17300_),
    .B1(_17475_),
    .B2(_17214_),
    .ZN(_05686_));
 NOR2_X1 _28046_ (.A1(_17364_),
    .A2(_05686_),
    .ZN(_05687_));
 AOI21_X1 _28047_ (.A(_05687_),
    .B1(_17475_),
    .B2(_17434_),
    .ZN(_05688_));
 NOR2_X1 _28048_ (.A1(_17459_),
    .A2(_05688_),
    .ZN(_05689_));
 OAI21_X1 _28049_ (.A(_18044_),
    .B1(_17461_),
    .B2(_18164_),
    .ZN(_05690_));
 OAI21_X1 _28050_ (.A(_18164_),
    .B1(_17364_),
    .B2(_17368_),
    .ZN(_05691_));
 OAI21_X1 _28051_ (.A(_17273_),
    .B1(_17441_),
    .B2(_17214_),
    .ZN(_05692_));
 AOI22_X1 _28052_ (.A1(_17294_),
    .A2(_05690_),
    .B1(_05691_),
    .B2(_05692_),
    .ZN(_05693_));
 OAI21_X1 _28053_ (.A(_17431_),
    .B1(_05693_),
    .B2(_17221_),
    .ZN(_05694_));
 NOR3_X2 _28054_ (.A1(_18351_),
    .A2(_05689_),
    .A3(_05694_),
    .ZN(_05695_));
 OAI21_X1 _28055_ (.A(_17963_),
    .B1(_17325_),
    .B2(_17228_),
    .ZN(_05696_));
 AOI22_X2 _28056_ (.A1(_17464_),
    .A2(_17987_),
    .B1(_17304_),
    .B2(_17371_),
    .ZN(_05697_));
 OAI221_X2 _28057_ (.A(_05696_),
    .B1(_05697_),
    .B2(_17468_),
    .C1(_17338_),
    .C2(_17461_),
    .ZN(_05698_));
 OAI22_X1 _28058_ (.A1(_17310_),
    .A2(_17989_),
    .B1(_17461_),
    .B2(_17987_),
    .ZN(_05699_));
 NAND2_X1 _28059_ (.A1(_17391_),
    .A2(_17486_),
    .ZN(_05700_));
 AOI221_X2 _28060_ (.A(_05698_),
    .B1(_05699_),
    .B2(_17325_),
    .C1(_05700_),
    .C2(_18186_),
    .ZN(_05701_));
 OAI21_X1 _28061_ (.A(_18214_),
    .B1(_17461_),
    .B2(_17987_),
    .ZN(_05702_));
 NAND2_X1 _28062_ (.A1(_17294_),
    .A2(_05702_),
    .ZN(_05703_));
 NAND4_X2 _28063_ (.A1(_17994_),
    .A2(_18193_),
    .A3(_05701_),
    .A4(_05703_),
    .ZN(_05704_));
 NAND2_X1 _28064_ (.A1(_17434_),
    .A2(_18120_),
    .ZN(_05705_));
 AOI22_X1 _28065_ (.A1(_17220_),
    .A2(_17360_),
    .B1(_18120_),
    .B2(_17213_),
    .ZN(_05706_));
 OAI21_X1 _28066_ (.A(_05705_),
    .B1(_05706_),
    .B2(_17319_),
    .ZN(_05707_));
 NAND2_X1 _28067_ (.A1(_17229_),
    .A2(_05707_),
    .ZN(_05708_));
 NAND3_X1 _28068_ (.A1(_17321_),
    .A2(_17434_),
    .A3(_17491_),
    .ZN(_05709_));
 OAI21_X1 _28069_ (.A(_18393_),
    .B1(_17437_),
    .B2(_17268_),
    .ZN(_05710_));
 NAND2_X1 _28070_ (.A1(_18364_),
    .A2(_05710_),
    .ZN(_05711_));
 NAND4_X1 _28071_ (.A1(_18362_),
    .A2(_05708_),
    .A3(_05709_),
    .A4(_05711_),
    .ZN(_05712_));
 NOR2_X1 _28072_ (.A1(_05704_),
    .A2(_05712_),
    .ZN(_05713_));
 NAND4_X4 _28073_ (.A1(_18424_),
    .A2(_18523_),
    .A3(_05695_),
    .A4(_05713_),
    .ZN(_05714_));
 NOR2_X4 _28074_ (.A1(_18105_),
    .A2(_05714_),
    .ZN(_05715_));
 INV_X1 _28075_ (.A(\block_reg[2][8] ),
    .ZN(_05716_));
 XNOR2_X1 _28076_ (.A(_05716_),
    .B(_17617_),
    .ZN(_05717_));
 OAI221_X1 _28077_ (.A(_16364_),
    .B1(_17741_),
    .B2(_04327_),
    .C1(_05717_),
    .C2(_18553_),
    .ZN(_05718_));
 XNOR2_X2 _28078_ (.A(_17891_),
    .B(_18560_),
    .ZN(_05719_));
 XOR2_X1 _28079_ (.A(_17780_),
    .B(_05719_),
    .Z(_05720_));
 XNOR2_X2 _28080_ (.A(_17604_),
    .B(_17848_),
    .ZN(_05721_));
 XNOR2_X1 _28081_ (.A(_17947_),
    .B(_05721_),
    .ZN(_05722_));
 XNOR2_X1 _28082_ (.A(_17906_),
    .B(_05722_),
    .ZN(_05723_));
 XNOR2_X1 _28083_ (.A(_05720_),
    .B(_05723_),
    .ZN(_05724_));
 AOI21_X1 _28084_ (.A(_05718_),
    .B1(_05724_),
    .B2(_19031_),
    .ZN(_05725_));
 AOI21_X1 _28085_ (.A(_05685_),
    .B1(_05715_),
    .B2(_05725_),
    .ZN(_00597_));
 AND4_X1 _28086_ (.A1(_18362_),
    .A2(_05708_),
    .A3(_05709_),
    .A4(_05711_),
    .ZN(_05726_));
 NAND2_X1 _28087_ (.A1(_17372_),
    .A2(_17491_),
    .ZN(_05727_));
 MUX2_X1 _28088_ (.A(_17318_),
    .B(_05727_),
    .S(_17272_),
    .Z(_05728_));
 OAI21_X1 _28089_ (.A(_18392_),
    .B1(_05728_),
    .B2(_17427_),
    .ZN(_05729_));
 NOR2_X1 _28090_ (.A1(_18009_),
    .A2(_05729_),
    .ZN(_05730_));
 NAND4_X2 _28091_ (.A1(_17341_),
    .A2(_18462_),
    .A3(_05726_),
    .A4(_05730_),
    .ZN(_05731_));
 OAI21_X1 _28092_ (.A(_17434_),
    .B1(_17384_),
    .B2(_17350_),
    .ZN(_05732_));
 AOI21_X1 _28093_ (.A(_17989_),
    .B1(_17397_),
    .B2(_05732_),
    .ZN(_05733_));
 AOI22_X2 _28094_ (.A1(_17366_),
    .A2(_17398_),
    .B1(_17456_),
    .B2(_17445_),
    .ZN(_05734_));
 AOI21_X1 _28095_ (.A(_17355_),
    .B1(_17366_),
    .B2(_18014_),
    .ZN(_05735_));
 AOI21_X1 _28096_ (.A(_18014_),
    .B1(_17434_),
    .B2(_17321_),
    .ZN(_05736_));
 OAI22_X1 _28097_ (.A1(_17374_),
    .A2(_05734_),
    .B1(_05735_),
    .B2(_05736_),
    .ZN(_05737_));
 NAND2_X1 _28098_ (.A1(_17313_),
    .A2(_17433_),
    .ZN(_05738_));
 AOI21_X1 _28099_ (.A(_05738_),
    .B1(_17474_),
    .B2(_17391_),
    .ZN(_05739_));
 OAI222_X2 _28100_ (.A1(_17305_),
    .A2(_17448_),
    .B1(_17418_),
    .B2(_17955_),
    .C1(_17439_),
    .C2(_17307_),
    .ZN(_05740_));
 NAND3_X1 _28101_ (.A1(_17276_),
    .A2(_17288_),
    .A3(_17433_),
    .ZN(_05741_));
 OAI21_X1 _28102_ (.A(_05741_),
    .B1(_17450_),
    .B2(_17276_),
    .ZN(_05742_));
 NAND4_X1 _28103_ (.A1(_17239_),
    .A2(_17281_),
    .A3(_17304_),
    .A4(_05742_),
    .ZN(_05743_));
 OAI221_X1 _28104_ (.A(_05743_),
    .B1(_17399_),
    .B2(_17317_),
    .C1(_17459_),
    .C2(_17391_),
    .ZN(_05744_));
 NOR3_X1 _28105_ (.A1(_05739_),
    .A2(_05740_),
    .A3(_05744_),
    .ZN(_05745_));
 AOI21_X1 _28106_ (.A(_18006_),
    .B1(_17485_),
    .B2(_17464_),
    .ZN(_05746_));
 MUX2_X1 _28107_ (.A(_17463_),
    .B(_18495_),
    .S(_17271_),
    .Z(_05747_));
 OAI221_X1 _28108_ (.A(_05745_),
    .B1(_05746_),
    .B2(_18214_),
    .C1(_17482_),
    .C2(_05747_),
    .ZN(_05748_));
 OR4_X1 _28109_ (.A1(_18508_),
    .A2(_05733_),
    .A3(_05737_),
    .A4(_05748_),
    .ZN(_05749_));
 AOI21_X1 _28110_ (.A(_18017_),
    .B1(_17463_),
    .B2(_18044_),
    .ZN(_05750_));
 AOI21_X1 _28111_ (.A(_05750_),
    .B1(_17369_),
    .B2(_17377_),
    .ZN(_05751_));
 OAI21_X1 _28112_ (.A(_18110_),
    .B1(_05751_),
    .B2(_17364_),
    .ZN(_05752_));
 NOR3_X2 _28113_ (.A1(_05731_),
    .A2(_05749_),
    .A3(_05752_),
    .ZN(_05753_));
 AOI21_X4 _28114_ (.A(_17379_),
    .B1(_18158_),
    .B2(_05753_),
    .ZN(_05754_));
 INV_X1 _28115_ (.A(_16553_),
    .ZN(_05755_));
 XOR2_X2 _28116_ (.A(\block_reg[2][9] ),
    .B(_17688_),
    .Z(_05756_));
 AOI221_X1 _28117_ (.A(_16367_),
    .B1(_05755_),
    .B2(_04564_),
    .C1(_05756_),
    .C2(_16370_),
    .ZN(_05757_));
 XNOR2_X1 _28118_ (.A(_17618_),
    .B(_17946_),
    .ZN(_05758_));
 XNOR2_X2 _28119_ (.A(_18243_),
    .B(_05758_),
    .ZN(_05759_));
 XNOR2_X1 _28120_ (.A(_17673_),
    .B(_05759_),
    .ZN(_05760_));
 XNOR2_X1 _28121_ (.A(_18262_),
    .B(_05760_),
    .ZN(_05761_));
 XNOR2_X1 _28122_ (.A(_17798_),
    .B(_05761_),
    .ZN(_05762_));
 OAI21_X1 _28123_ (.A(_05757_),
    .B1(_05762_),
    .B2(_17204_),
    .ZN(_05763_));
 OAI22_X1 _28124_ (.A1(\core.dec_block.block_w0_reg[9] ),
    .A2(_16366_),
    .B1(_05754_),
    .B2(_05763_),
    .ZN(_05764_));
 INV_X1 _28125_ (.A(_05764_),
    .ZN(_00598_));
 AOI21_X1 _28126_ (.A(_16354_),
    .B1(_18568_),
    .B2(_16360_),
    .ZN(_05765_));
 NOR2_X1 _28127_ (.A1(_16258_),
    .A2(_05765_),
    .ZN(_05766_));
 NOR2_X1 _28128_ (.A1(_16353_),
    .A2(_05766_),
    .ZN(_05767_));
 CLKBUF_X3 _28129_ (.A(_05767_),
    .Z(_05768_));
 CLKBUF_X3 _28130_ (.A(_05768_),
    .Z(_05769_));
 OR2_X1 _28131_ (.A1(_16353_),
    .A2(_05766_),
    .ZN(_05770_));
 CLKBUF_X3 _28132_ (.A(_05770_),
    .Z(_05771_));
 BUF_X4 _28133_ (.A(_05771_),
    .Z(_05772_));
 XNOR2_X1 _28134_ (.A(\block_reg[2][0] ),
    .B(_17778_),
    .ZN(_05773_));
 BUF_X4 _28135_ (.A(_17709_),
    .Z(_05774_));
 OAI221_X1 _28136_ (.A(_05772_),
    .B1(_05773_),
    .B2(_05774_),
    .C1(_03525_),
    .C2(_04264_),
    .ZN(_05775_));
 XNOR2_X2 _28137_ (.A(_17618_),
    .B(_17906_),
    .ZN(_05776_));
 XNOR2_X1 _28138_ (.A(_18261_),
    .B(_05776_),
    .ZN(_05777_));
 XOR2_X1 _28139_ (.A(_17574_),
    .B(_17658_),
    .Z(_05778_));
 XNOR2_X1 _28140_ (.A(_17762_),
    .B(_05778_),
    .ZN(_05779_));
 XNOR2_X2 _28141_ (.A(_05777_),
    .B(_05779_),
    .ZN(_05780_));
 XNOR2_X2 _28142_ (.A(_17948_),
    .B(_05780_),
    .ZN(_05781_));
 CLKBUF_X3 _28143_ (.A(_17748_),
    .Z(_05782_));
 AOI21_X1 _28144_ (.A(_05775_),
    .B1(_05781_),
    .B2(_05782_),
    .ZN(_05783_));
 AOI22_X1 _28145_ (.A1(_03524_),
    .A2(_05769_),
    .B1(_05783_),
    .B2(_16851_),
    .ZN(_00599_));
 BUF_X4 _28146_ (.A(_05772_),
    .Z(_05784_));
 XNOR2_X1 _28147_ (.A(\block_reg[3][10] ),
    .B(_19411_),
    .ZN(_05785_));
 AOI21_X1 _28148_ (.A(_05768_),
    .B1(_05785_),
    .B2(_16372_),
    .ZN(_05786_));
 XOR2_X1 _28149_ (.A(_18982_),
    .B(_19016_),
    .Z(_05787_));
 XNOR2_X1 _28150_ (.A(_19224_),
    .B(_05787_),
    .ZN(_05788_));
 XNOR2_X1 _28151_ (.A(_03743_),
    .B(_05788_),
    .ZN(_05789_));
 XOR2_X1 _28152_ (.A(_19285_),
    .B(_19430_),
    .Z(_05790_));
 XNOR2_X1 _28153_ (.A(_03745_),
    .B(_05790_),
    .ZN(_05791_));
 XNOR2_X1 _28154_ (.A(_05789_),
    .B(_05791_),
    .ZN(_05792_));
 BUF_X4 _28155_ (.A(_17203_),
    .Z(_05793_));
 OAI221_X1 _28156_ (.A(_05786_),
    .B1(_05792_),
    .B2(_05793_),
    .C1(_16556_),
    .C2(_05158_),
    .ZN(_05794_));
 OAI22_X1 _28157_ (.A1(\core.dec_block.block_w1_reg[10] ),
    .A2(_05784_),
    .B1(_05794_),
    .B2(_17503_),
    .ZN(_05795_));
 INV_X1 _28158_ (.A(_05795_),
    .ZN(_00600_));
 XNOR2_X1 _28159_ (.A(_19274_),
    .B(_19299_),
    .ZN(_05796_));
 XNOR2_X2 _28160_ (.A(_03763_),
    .B(_05796_),
    .ZN(_05797_));
 XNOR2_X2 _28161_ (.A(_19027_),
    .B(_19441_),
    .ZN(_05798_));
 XOR2_X1 _28162_ (.A(_19261_),
    .B(_05798_),
    .Z(_05799_));
 XNOR2_X1 _28163_ (.A(_19003_),
    .B(_05799_),
    .ZN(_05800_));
 XNOR2_X1 _28164_ (.A(_05797_),
    .B(_05800_),
    .ZN(_05801_));
 XNOR2_X2 _28165_ (.A(_19229_),
    .B(_05801_),
    .ZN(_05802_));
 XNOR2_X2 _28166_ (.A(_19246_),
    .B(_03918_),
    .ZN(_05803_));
 XNOR2_X1 _28167_ (.A(_19413_),
    .B(_03742_),
    .ZN(_05804_));
 XNOR2_X1 _28168_ (.A(_05803_),
    .B(_05804_),
    .ZN(_05805_));
 XNOR2_X1 _28169_ (.A(_05802_),
    .B(_05805_),
    .ZN(_05806_));
 NOR2_X1 _28170_ (.A1(_17504_),
    .A2(_05806_),
    .ZN(_05807_));
 XNOR2_X2 _28171_ (.A(\block_reg[3][11] ),
    .B(_03343_),
    .ZN(_05808_));
 OAI221_X2 _28172_ (.A(_05772_),
    .B1(_05808_),
    .B2(_18078_),
    .C1(_05385_),
    .C2(_17741_),
    .ZN(_05809_));
 NOR3_X1 _28173_ (.A1(_18051_),
    .A2(_05807_),
    .A3(_05809_),
    .ZN(_05810_));
 AOI21_X1 _28174_ (.A(_05810_),
    .B1(_05769_),
    .B2(_17333_),
    .ZN(_00601_));
 XNOR2_X2 _28175_ (.A(_19224_),
    .B(_03921_),
    .ZN(_05811_));
 XNOR2_X1 _28176_ (.A(_19274_),
    .B(_03776_),
    .ZN(_05812_));
 XNOR2_X1 _28177_ (.A(_05811_),
    .B(_05812_),
    .ZN(_05813_));
 XNOR2_X1 _28178_ (.A(_03789_),
    .B(_05813_),
    .ZN(_05814_));
 XNOR2_X1 _28179_ (.A(_03784_),
    .B(_05814_),
    .ZN(_05815_));
 XNOR2_X1 _28180_ (.A(_03741_),
    .B(_05815_),
    .ZN(_05816_));
 NAND2_X1 _28181_ (.A1(_17749_),
    .A2(_05816_),
    .ZN(_05817_));
 XOR2_X2 _28182_ (.A(\block_reg[3][12] ),
    .B(_03774_),
    .Z(_05818_));
 OAI22_X1 _28183_ (.A1(_18052_),
    .A2(_05537_),
    .B1(_05818_),
    .B2(_18078_),
    .ZN(_05819_));
 NOR3_X1 _28184_ (.A1(_18228_),
    .A2(_05768_),
    .A3(_05819_),
    .ZN(_05820_));
 AOI22_X1 _28185_ (.A1(_05525_),
    .A2(_05769_),
    .B1(_05817_),
    .B2(_05820_),
    .ZN(_00602_));
 NOR2_X1 _28186_ (.A1(\core.dec_block.block_w1_reg[13] ),
    .A2(_05784_),
    .ZN(_05821_));
 XOR2_X2 _28187_ (.A(\block_reg[3][13] ),
    .B(_18969_),
    .Z(_05822_));
 OAI22_X1 _28188_ (.A1(_16556_),
    .A2(_17062_),
    .B1(_05822_),
    .B2(_04266_),
    .ZN(_05823_));
 NOR2_X1 _28189_ (.A1(_05768_),
    .A2(_05823_),
    .ZN(_05824_));
 XNOR2_X1 _28190_ (.A(_03326_),
    .B(_03333_),
    .ZN(_05825_));
 XNOR2_X2 _28191_ (.A(_19430_),
    .B(_05825_),
    .ZN(_05826_));
 XOR2_X2 _28192_ (.A(_03791_),
    .B(_05826_),
    .Z(_05827_));
 XNOR2_X1 _28193_ (.A(_18922_),
    .B(_03776_),
    .ZN(_05828_));
 XOR2_X1 _28194_ (.A(_19002_),
    .B(_03775_),
    .Z(_05829_));
 XNOR2_X1 _28195_ (.A(_05828_),
    .B(_05829_),
    .ZN(_05830_));
 XOR2_X1 _28196_ (.A(_19414_),
    .B(_03760_),
    .Z(_05831_));
 XNOR2_X1 _28197_ (.A(_05830_),
    .B(_05831_),
    .ZN(_05832_));
 XNOR2_X2 _28198_ (.A(_05827_),
    .B(_05832_),
    .ZN(_05833_));
 AOI21_X1 _28199_ (.A(_18398_),
    .B1(_05833_),
    .B2(_19031_),
    .ZN(_05834_));
 AOI21_X1 _28200_ (.A(_05821_),
    .B1(_05824_),
    .B2(_05834_),
    .ZN(_00603_));
 NOR2_X1 _28201_ (.A1(\core.dec_block.block_w1_reg[14] ),
    .A2(_05784_),
    .ZN(_05835_));
 OAI21_X1 _28202_ (.A(_05771_),
    .B1(_03596_),
    .B2(_16554_),
    .ZN(_05836_));
 XNOR2_X2 _28203_ (.A(_18970_),
    .B(_03775_),
    .ZN(_05837_));
 XNOR2_X2 _28204_ (.A(_18897_),
    .B(_03961_),
    .ZN(_05838_));
 XOR2_X2 _28205_ (.A(_05837_),
    .B(_05838_),
    .Z(_05839_));
 XNOR2_X2 _28206_ (.A(_18921_),
    .B(_18956_),
    .ZN(_05840_));
 XNOR2_X2 _28207_ (.A(_03919_),
    .B(_05840_),
    .ZN(_05841_));
 XNOR2_X2 _28208_ (.A(_05839_),
    .B(_05841_),
    .ZN(_05842_));
 XNOR2_X2 _28209_ (.A(_05803_),
    .B(_05842_),
    .ZN(_05843_));
 XNOR2_X2 _28210_ (.A(\block_reg[3][14] ),
    .B(_19223_),
    .ZN(_05844_));
 AOI221_X2 _28211_ (.A(_05836_),
    .B1(_05843_),
    .B2(_17748_),
    .C1(_16372_),
    .C2(_05844_),
    .ZN(_05845_));
 AOI21_X1 _28212_ (.A(_05835_),
    .B1(_05845_),
    .B2(_18465_),
    .ZN(_00604_));
 NOR2_X1 _28213_ (.A1(\core.dec_block.block_w1_reg[15] ),
    .A2(_05784_),
    .ZN(_05846_));
 BUF_X4 _28214_ (.A(_05771_),
    .Z(_05847_));
 XOR2_X2 _28215_ (.A(\block_reg[3][15] ),
    .B(_18941_),
    .Z(_05848_));
 OAI221_X1 _28216_ (.A(_05847_),
    .B1(_05848_),
    .B2(_18466_),
    .C1(_05115_),
    .C2(_18399_),
    .ZN(_05849_));
 XOR2_X1 _28217_ (.A(_19002_),
    .B(_03922_),
    .Z(_05850_));
 XNOR2_X1 _28218_ (.A(_03961_),
    .B(_05850_),
    .ZN(_05851_));
 XNOR2_X2 _28219_ (.A(_19260_),
    .B(_05837_),
    .ZN(_05852_));
 XNOR2_X2 _28220_ (.A(_05811_),
    .B(_05852_),
    .ZN(_05853_));
 XNOR2_X2 _28221_ (.A(_05851_),
    .B(_05853_),
    .ZN(_05854_));
 AOI21_X1 _28222_ (.A(_05849_),
    .B1(_05854_),
    .B2(_04370_),
    .ZN(_05855_));
 AOI21_X1 _28223_ (.A(_05846_),
    .B1(_05855_),
    .B2(_18526_),
    .ZN(_00605_));
 NOR2_X1 _28224_ (.A1(\core.dec_block.block_w1_reg[16] ),
    .A2(_05784_),
    .ZN(_05856_));
 XNOR2_X1 _28225_ (.A(\block_reg[0][16] ),
    .B(_18870_),
    .ZN(_05857_));
 OAI221_X1 _28226_ (.A(_05847_),
    .B1(_05857_),
    .B2(_18466_),
    .C1(_17139_),
    .C2(_18399_),
    .ZN(_05858_));
 XNOR2_X2 _28227_ (.A(_16551_),
    .B(_04263_),
    .ZN(_05859_));
 XOR2_X1 _28228_ (.A(_05188_),
    .B(_05859_),
    .Z(_05860_));
 XNOR2_X1 _28229_ (.A(_04590_),
    .B(_04812_),
    .ZN(_05861_));
 XNOR2_X1 _28230_ (.A(_05860_),
    .B(_05861_),
    .ZN(_05862_));
 XNOR2_X1 _28231_ (.A(_05265_),
    .B(_05862_),
    .ZN(_05863_));
 AOI21_X1 _28232_ (.A(_05858_),
    .B1(_05863_),
    .B2(_04370_),
    .ZN(_05864_));
 AOI21_X1 _28233_ (.A(_05856_),
    .B1(_05864_),
    .B2(_18848_),
    .ZN(_00606_));
 XNOR2_X2 _28234_ (.A(\block_reg[0][17] ),
    .B(_19191_),
    .ZN(_05865_));
 AOI21_X1 _28235_ (.A(_05767_),
    .B1(_05865_),
    .B2(_16371_),
    .ZN(_05866_));
 OAI21_X1 _28236_ (.A(_05866_),
    .B1(_03616_),
    .B2(_18479_),
    .ZN(_05867_));
 XNOR2_X2 _28237_ (.A(_18550_),
    .B(_03857_),
    .ZN(_05868_));
 XNOR2_X2 _28238_ (.A(_18871_),
    .B(_05868_),
    .ZN(_05869_));
 XNOR2_X2 _28239_ (.A(_04813_),
    .B(_05869_),
    .ZN(_05870_));
 XNOR2_X1 _28240_ (.A(_03510_),
    .B(_04812_),
    .ZN(_05871_));
 XOR2_X1 _28241_ (.A(_04811_),
    .B(_05871_),
    .Z(_05872_));
 XNOR2_X1 _28242_ (.A(_05870_),
    .B(_05872_),
    .ZN(_05873_));
 AOI21_X1 _28243_ (.A(_05867_),
    .B1(_05873_),
    .B2(_05782_),
    .ZN(_05874_));
 AOI22_X1 _28244_ (.A1(_03598_),
    .A2(_05769_),
    .B1(_05874_),
    .B2(_19179_),
    .ZN(_00607_));
 BUF_X4 _28245_ (.A(_05772_),
    .Z(_05875_));
 NOR2_X1 _28246_ (.A1(\core.dec_block.block_w1_reg[18] ),
    .A2(_05875_),
    .ZN(_05876_));
 XNOR2_X2 _28247_ (.A(\block_reg[0][18] ),
    .B(_19384_),
    .ZN(_05877_));
 OAI221_X1 _28248_ (.A(_05847_),
    .B1(_05877_),
    .B2(_18466_),
    .C1(_05176_),
    .C2(_18399_),
    .ZN(_05878_));
 XNOR2_X1 _28249_ (.A(_18871_),
    .B(_03915_),
    .ZN(_05879_));
 XNOR2_X1 _28250_ (.A(_16551_),
    .B(_05879_),
    .ZN(_05880_));
 XNOR2_X1 _28251_ (.A(_04924_),
    .B(_05880_),
    .ZN(_05881_));
 XNOR2_X2 _28252_ (.A(_19192_),
    .B(_04809_),
    .ZN(_05882_));
 XNOR2_X1 _28253_ (.A(_04589_),
    .B(_04699_),
    .ZN(_05883_));
 XNOR2_X1 _28254_ (.A(_05882_),
    .B(_05883_),
    .ZN(_05884_));
 XNOR2_X1 _28255_ (.A(_05881_),
    .B(_05884_),
    .ZN(_05885_));
 AOI21_X1 _28256_ (.A(_05878_),
    .B1(_05885_),
    .B2(_04370_),
    .ZN(_05886_));
 AOI21_X1 _28257_ (.A(_05876_),
    .B1(_05886_),
    .B2(_19371_),
    .ZN(_00608_));
 XOR2_X2 _28258_ (.A(\block_reg[0][19] ),
    .B(_03286_),
    .Z(_05887_));
 OAI221_X1 _28259_ (.A(_05772_),
    .B1(_05887_),
    .B2(_05774_),
    .C1(_05406_),
    .C2(_04264_),
    .ZN(_05888_));
 XNOR2_X1 _28260_ (.A(_04724_),
    .B(_05871_),
    .ZN(_05889_));
 XNOR2_X1 _28261_ (.A(_04366_),
    .B(_04593_),
    .ZN(_05890_));
 XNOR2_X2 _28262_ (.A(_05889_),
    .B(_05890_),
    .ZN(_05891_));
 XNOR2_X2 _28263_ (.A(_04819_),
    .B(_04941_),
    .ZN(_05892_));
 XNOR2_X1 _28264_ (.A(_04594_),
    .B(_05892_),
    .ZN(_05893_));
 XNOR2_X2 _28265_ (.A(_05891_),
    .B(_05893_),
    .ZN(_05894_));
 XOR2_X1 _28266_ (.A(_17740_),
    .B(_04834_),
    .Z(_05895_));
 XNOR2_X1 _28267_ (.A(_05869_),
    .B(_05895_),
    .ZN(_05896_));
 XNOR2_X1 _28268_ (.A(_05894_),
    .B(_05896_),
    .ZN(_05897_));
 AOI21_X1 _28269_ (.A(_05888_),
    .B1(_05897_),
    .B2(_05782_),
    .ZN(_05898_));
 AOI22_X1 _28270_ (.A1(_05394_),
    .A2(_05769_),
    .B1(_05898_),
    .B2(_19519_),
    .ZN(_00609_));
 NOR2_X1 _28271_ (.A1(\core.dec_block.block_w1_reg[1] ),
    .A2(_05875_),
    .ZN(_05899_));
 INV_X1 _28272_ (.A(\block_reg[2][1] ),
    .ZN(_05900_));
 XNOR2_X1 _28273_ (.A(_05900_),
    .B(_17671_),
    .ZN(_05901_));
 BUF_X4 _28274_ (.A(_16555_),
    .Z(_05902_));
 OAI221_X1 _28275_ (.A(_05847_),
    .B1(_05901_),
    .B2(_18466_),
    .C1(_05177_),
    .C2(_05902_),
    .ZN(_05903_));
 XOR2_X2 _28276_ (.A(_18247_),
    .B(_05719_),
    .Z(_05904_));
 XNOR2_X2 _28277_ (.A(_17761_),
    .B(_17779_),
    .ZN(_05905_));
 XNOR2_X1 _28278_ (.A(_17552_),
    .B(_17935_),
    .ZN(_05906_));
 XNOR2_X1 _28279_ (.A(_17643_),
    .B(_18259_),
    .ZN(_05907_));
 XNOR2_X1 _28280_ (.A(_05906_),
    .B(_05907_),
    .ZN(_05908_));
 XNOR2_X1 _28281_ (.A(_05905_),
    .B(_05908_),
    .ZN(_05909_));
 XNOR2_X2 _28282_ (.A(_05904_),
    .B(_05909_),
    .ZN(_05910_));
 AOI21_X1 _28283_ (.A(_05903_),
    .B1(_05910_),
    .B2(_04370_),
    .ZN(_05911_));
 AOI21_X1 _28284_ (.A(_05899_),
    .B1(_05911_),
    .B2(_03498_),
    .ZN(_00610_));
 NOR2_X1 _28285_ (.A1(\core.dec_block.block_w1_reg[20] ),
    .A2(_05875_),
    .ZN(_05912_));
 XNOR2_X2 _28286_ (.A(\block_reg[0][20] ),
    .B(_03723_),
    .ZN(_05913_));
 OAI221_X1 _28287_ (.A(_05847_),
    .B1(_05913_),
    .B2(_18466_),
    .C1(_05524_),
    .C2(_05902_),
    .ZN(_05914_));
 XNOR2_X2 _28288_ (.A(_04591_),
    .B(_04725_),
    .ZN(_05915_));
 XNOR2_X1 _28289_ (.A(_05183_),
    .B(_05262_),
    .ZN(_05916_));
 XNOR2_X1 _28290_ (.A(_04819_),
    .B(_05015_),
    .ZN(_05917_));
 XNOR2_X1 _28291_ (.A(_04918_),
    .B(_05917_),
    .ZN(_05918_));
 XNOR2_X1 _28292_ (.A(_05916_),
    .B(_05918_),
    .ZN(_05919_));
 XNOR2_X1 _28293_ (.A(_05915_),
    .B(_05919_),
    .ZN(_05920_));
 CLKBUF_X3 _28294_ (.A(_17748_),
    .Z(_05921_));
 AOI21_X1 _28295_ (.A(_05914_),
    .B1(_05920_),
    .B2(_05921_),
    .ZN(_05922_));
 AOI21_X1 _28296_ (.A(_05912_),
    .B1(_05922_),
    .B2(_03698_),
    .ZN(_00611_));
 XNOR2_X1 _28297_ (.A(\block_reg[0][21] ),
    .B(_03856_),
    .ZN(_05923_));
 OAI221_X1 _28298_ (.A(_05772_),
    .B1(_05923_),
    .B2(_17710_),
    .C1(_16943_),
    .C2(_18052_),
    .ZN(_05924_));
 XNOR2_X2 _28299_ (.A(_04312_),
    .B(_04365_),
    .ZN(_05925_));
 XNOR2_X1 _28300_ (.A(_04943_),
    .B(_05925_),
    .ZN(_05926_));
 XNOR2_X1 _28301_ (.A(_04684_),
    .B(_05008_),
    .ZN(_05927_));
 XNOR2_X1 _28302_ (.A(_05926_),
    .B(_05927_),
    .ZN(_05928_));
 XNOR2_X1 _28303_ (.A(_04724_),
    .B(_04919_),
    .ZN(_05929_));
 XNOR2_X1 _28304_ (.A(_18478_),
    .B(_05929_),
    .ZN(_05930_));
 XOR2_X2 _28305_ (.A(_04833_),
    .B(_04923_),
    .Z(_05931_));
 XOR2_X1 _28306_ (.A(_05930_),
    .B(_05931_),
    .Z(_05932_));
 XNOR2_X1 _28307_ (.A(_05928_),
    .B(_05932_),
    .ZN(_05933_));
 NOR2_X1 _28308_ (.A1(_05793_),
    .A2(_05933_),
    .ZN(_05934_));
 NOR3_X1 _28309_ (.A1(_03845_),
    .A2(_05924_),
    .A3(_05934_),
    .ZN(_05935_));
 AOI21_X1 _28310_ (.A(_05935_),
    .B1(_05769_),
    .B2(_16876_),
    .ZN(_00612_));
 XNOR2_X2 _28311_ (.A(\block_reg[0][22] ),
    .B(_03914_),
    .ZN(_05936_));
 OAI221_X1 _28312_ (.A(_05771_),
    .B1(_05936_),
    .B2(_05774_),
    .C1(_16978_),
    .C2(_04264_),
    .ZN(_05937_));
 XNOR2_X2 _28313_ (.A(_04723_),
    .B(_04833_),
    .ZN(_05938_));
 XNOR2_X1 _28314_ (.A(_04937_),
    .B(_05938_),
    .ZN(_05939_));
 XNOR2_X1 _28315_ (.A(_05892_),
    .B(_05939_),
    .ZN(_05940_));
 XNOR2_X2 _28316_ (.A(_04943_),
    .B(_05940_),
    .ZN(_05941_));
 XNOR2_X2 _28317_ (.A(_18478_),
    .B(_04589_),
    .ZN(_05942_));
 XOR2_X1 _28318_ (.A(_04311_),
    .B(_05015_),
    .Z(_05943_));
 XNOR2_X1 _28319_ (.A(_05942_),
    .B(_05943_),
    .ZN(_05944_));
 XNOR2_X1 _28320_ (.A(_05941_),
    .B(_05944_),
    .ZN(_05945_));
 AOI21_X1 _28321_ (.A(_05937_),
    .B1(_05945_),
    .B2(_05782_),
    .ZN(_05946_));
 AOI22_X1 _28322_ (.A1(_16944_),
    .A2(_05769_),
    .B1(_05946_),
    .B2(_03893_),
    .ZN(_00613_));
 OAI21_X1 _28323_ (.A(_05771_),
    .B1(_03627_),
    .B2(_16554_),
    .ZN(_05947_));
 XNOR2_X1 _28324_ (.A(\block_reg[0][23] ),
    .B(_03975_),
    .ZN(_05948_));
 AOI21_X1 _28325_ (.A(_05947_),
    .B1(_05948_),
    .B2(_16371_),
    .ZN(_05949_));
 XNOR2_X2 _28326_ (.A(_04349_),
    .B(_05016_),
    .ZN(_05950_));
 XNOR2_X1 _28327_ (.A(_05262_),
    .B(_05868_),
    .ZN(_05951_));
 XNOR2_X2 _28328_ (.A(_05950_),
    .B(_05951_),
    .ZN(_05952_));
 XNOR2_X1 _28329_ (.A(_04813_),
    .B(_05190_),
    .ZN(_05953_));
 XNOR2_X1 _28330_ (.A(_05952_),
    .B(_05953_),
    .ZN(_05954_));
 OAI21_X1 _28331_ (.A(_05949_),
    .B1(_05954_),
    .B2(_17504_),
    .ZN(_05955_));
 NOR2_X1 _28332_ (.A1(_03955_),
    .A2(_05955_),
    .ZN(_05956_));
 INV_X1 _28333_ (.A(_18577_),
    .ZN(_05957_));
 AOI21_X1 _28334_ (.A(_05956_),
    .B1(_05769_),
    .B2(_05957_),
    .ZN(_00614_));
 NOR2_X1 _28335_ (.A1(\core.dec_block.block_w1_reg[24] ),
    .A2(_05875_),
    .ZN(_05958_));
 INV_X1 _28336_ (.A(\block_reg[1][24] ),
    .ZN(_05959_));
 XNOR2_X1 _28337_ (.A(_05959_),
    .B(_17096_),
    .ZN(_05960_));
 BUF_X4 _28338_ (.A(_17709_),
    .Z(_05961_));
 OAI221_X1 _28339_ (.A(_04251_),
    .B1(_05960_),
    .B2(_05961_),
    .C1(_17097_),
    .C2(_05902_),
    .ZN(_05962_));
 XNOR2_X2 _28340_ (.A(_03542_),
    .B(_03596_),
    .ZN(_05963_));
 XOR2_X1 _28341_ (.A(_03523_),
    .B(_05162_),
    .Z(_05964_));
 XNOR2_X1 _28342_ (.A(_05351_),
    .B(_05964_),
    .ZN(_05965_));
 XNOR2_X1 _28343_ (.A(_05963_),
    .B(_05965_),
    .ZN(_05966_));
 AOI21_X1 _28344_ (.A(_05962_),
    .B1(_05966_),
    .B2(_05921_),
    .ZN(_05967_));
 AOI21_X1 _28345_ (.A(_05958_),
    .B1(_05967_),
    .B2(_05784_),
    .ZN(_00615_));
 NOR2_X1 _28346_ (.A1(\core.dec_block.block_w1_reg[25] ),
    .A2(_05875_),
    .ZN(_05968_));
 XNOR2_X1 _28347_ (.A(\block_reg[1][25] ),
    .B(_03555_),
    .ZN(_05969_));
 OAI221_X2 _28348_ (.A(_05847_),
    .B1(_05969_),
    .B2(_05961_),
    .C1(_03556_),
    .C2(_05902_),
    .ZN(_05970_));
 XNOR2_X2 _28349_ (.A(_03627_),
    .B(_05115_),
    .ZN(_05971_));
 XNOR2_X1 _28350_ (.A(_16943_),
    .B(_05971_),
    .ZN(_05972_));
 XNOR2_X1 _28351_ (.A(_03576_),
    .B(_05972_),
    .ZN(_05973_));
 XNOR2_X1 _28352_ (.A(_17141_),
    .B(_05973_),
    .ZN(_05974_));
 XNOR2_X1 _28353_ (.A(_05348_),
    .B(_05974_),
    .ZN(_05975_));
 AOI21_X1 _28354_ (.A(_05970_),
    .B1(_05975_),
    .B2(_05921_),
    .ZN(_05976_));
 AOI21_X1 _28355_ (.A(_05968_),
    .B1(_05976_),
    .B2(_04538_),
    .ZN(_00616_));
 XNOR2_X1 _28356_ (.A(_17012_),
    .B(_03596_),
    .ZN(_05977_));
 XNOR2_X2 _28357_ (.A(_17097_),
    .B(_03541_),
    .ZN(_05978_));
 XNOR2_X1 _28358_ (.A(_05977_),
    .B(_05978_),
    .ZN(_05979_));
 XNOR2_X2 _28359_ (.A(_05393_),
    .B(_05979_),
    .ZN(_05980_));
 XNOR2_X1 _28360_ (.A(_05158_),
    .B(_05592_),
    .ZN(_05981_));
 XNOR2_X1 _28361_ (.A(_05179_),
    .B(_05981_),
    .ZN(_05982_));
 XNOR2_X1 _28362_ (.A(_05345_),
    .B(_05982_),
    .ZN(_05983_));
 XNOR2_X1 _28363_ (.A(_05980_),
    .B(_05983_),
    .ZN(_05984_));
 NOR2_X1 _28364_ (.A1(_17504_),
    .A2(_05984_),
    .ZN(_05985_));
 XNOR2_X2 _28365_ (.A(\block_reg[1][26] ),
    .B(_05137_),
    .ZN(_05986_));
 OAI221_X2 _28366_ (.A(_05772_),
    .B1(_05986_),
    .B2(_18078_),
    .C1(_05138_),
    .C2(_17741_),
    .ZN(_05987_));
 NOR3_X1 _28367_ (.A1(_04657_),
    .A2(_05985_),
    .A3(_05987_),
    .ZN(_05988_));
 INV_X1 _28368_ (.A(\core.dec_block.block_w1_reg[26] ),
    .ZN(_05989_));
 AOI21_X1 _28369_ (.A(_05988_),
    .B1(_05769_),
    .B2(_05989_),
    .ZN(_00617_));
 NOR2_X1 _28370_ (.A1(\core.dec_block.block_w1_reg[27] ),
    .A2(_05875_),
    .ZN(_05990_));
 OAI21_X1 _28371_ (.A(_05847_),
    .B1(_05362_),
    .B2(_05021_),
    .ZN(_05991_));
 XOR2_X1 _28372_ (.A(\block_reg[1][27] ),
    .B(_05361_),
    .Z(_05992_));
 AOI21_X1 _28373_ (.A(_05991_),
    .B1(_05992_),
    .B2(_16372_),
    .ZN(_05993_));
 XNOR2_X2 _28374_ (.A(_16943_),
    .B(_05596_),
    .ZN(_05994_));
 XNOR2_X2 _28375_ (.A(_17012_),
    .B(_17139_),
    .ZN(_05995_));
 XNOR2_X1 _28376_ (.A(_05116_),
    .B(_05995_),
    .ZN(_05996_));
 XNOR2_X1 _28377_ (.A(_03576_),
    .B(_05996_),
    .ZN(_05997_));
 XNOR2_X1 _28378_ (.A(_05994_),
    .B(_05997_),
    .ZN(_05998_));
 XNOR2_X2 _28379_ (.A(_03558_),
    .B(_05998_),
    .ZN(_05999_));
 XOR2_X1 _28380_ (.A(_05407_),
    .B(_05540_),
    .Z(_06000_));
 XNOR2_X1 _28381_ (.A(_05385_),
    .B(_05592_),
    .ZN(_06001_));
 XNOR2_X1 _28382_ (.A(_06000_),
    .B(_06001_),
    .ZN(_06002_));
 XNOR2_X1 _28383_ (.A(_05999_),
    .B(_06002_),
    .ZN(_06003_));
 AOI21_X1 _28384_ (.A(_04792_),
    .B1(_06003_),
    .B2(_19031_),
    .ZN(_06004_));
 AOI21_X1 _28385_ (.A(_05990_),
    .B1(_05993_),
    .B2(_06004_),
    .ZN(_00618_));
 NOR2_X1 _28386_ (.A1(\core.dec_block.block_w1_reg[28] ),
    .A2(_05875_),
    .ZN(_06005_));
 XNOR2_X1 _28387_ (.A(\block_reg[1][28] ),
    .B(_05509_),
    .ZN(_06006_));
 OAI221_X1 _28388_ (.A(_05847_),
    .B1(_06006_),
    .B2(_05961_),
    .C1(_05510_),
    .C2(_05902_),
    .ZN(_06007_));
 XOR2_X2 _28389_ (.A(_05161_),
    .B(_05348_),
    .Z(_06008_));
 XNOR2_X2 _28390_ (.A(_05494_),
    .B(_06008_),
    .ZN(_06009_));
 XNOR2_X2 _28391_ (.A(_05537_),
    .B(_05608_),
    .ZN(_06010_));
 XNOR2_X1 _28392_ (.A(_05614_),
    .B(_06010_),
    .ZN(_06011_));
 XNOR2_X1 _28393_ (.A(_06009_),
    .B(_06011_),
    .ZN(_06012_));
 AOI21_X1 _28394_ (.A(_06007_),
    .B1(_06012_),
    .B2(_05921_),
    .ZN(_06013_));
 AOI21_X1 _28395_ (.A(_06005_),
    .B1(_06013_),
    .B2(_04902_),
    .ZN(_00619_));
 INV_X1 _28396_ (.A(\block_reg[1][29] ),
    .ZN(_06014_));
 XNOR2_X1 _28397_ (.A(_06014_),
    .B(_17078_),
    .ZN(_06015_));
 OAI22_X1 _28398_ (.A1(_19180_),
    .A2(_17079_),
    .B1(_06015_),
    .B2(_18552_),
    .ZN(_06016_));
 XNOR2_X2 _28399_ (.A(_16875_),
    .B(_05392_),
    .ZN(_06017_));
 XNOR2_X1 _28400_ (.A(_17062_),
    .B(_05524_),
    .ZN(_06018_));
 XNOR2_X2 _28401_ (.A(_05386_),
    .B(_06018_),
    .ZN(_06019_));
 XOR2_X1 _28402_ (.A(_06017_),
    .B(_06019_),
    .Z(_06020_));
 XNOR2_X1 _28403_ (.A(_05512_),
    .B(_06020_),
    .ZN(_06021_));
 XNOR2_X1 _28404_ (.A(_05594_),
    .B(_06021_),
    .ZN(_06022_));
 NOR2_X1 _28405_ (.A1(_17203_),
    .A2(_06022_),
    .ZN(_06023_));
 NOR4_X1 _28406_ (.A1(_05003_),
    .A2(_05768_),
    .A3(_06016_),
    .A4(_06023_),
    .ZN(_06024_));
 AOI21_X1 _28407_ (.A(_06024_),
    .B1(_05769_),
    .B2(_17065_),
    .ZN(_00620_));
 OAI21_X1 _28408_ (.A(_05772_),
    .B1(_05392_),
    .B2(_18479_),
    .ZN(_06025_));
 XNOR2_X1 _28409_ (.A(\block_reg[2][2] ),
    .B(_17534_),
    .ZN(_06026_));
 AOI21_X1 _28410_ (.A(_06025_),
    .B1(_06026_),
    .B2(_16372_),
    .ZN(_06027_));
 XNOR2_X1 _28411_ (.A(_17779_),
    .B(_17906_),
    .ZN(_06028_));
 XNOR2_X2 _28412_ (.A(_18245_),
    .B(_06028_),
    .ZN(_06029_));
 XOR2_X1 _28413_ (.A(_17563_),
    .B(_17796_),
    .Z(_06030_));
 XNOR2_X2 _28414_ (.A(_17574_),
    .B(_17702_),
    .ZN(_06031_));
 XNOR2_X1 _28415_ (.A(_06030_),
    .B(_06031_),
    .ZN(_06032_));
 XNOR2_X2 _28416_ (.A(_17673_),
    .B(_06032_),
    .ZN(_06033_));
 XNOR2_X2 _28417_ (.A(_06029_),
    .B(_06033_),
    .ZN(_06034_));
 AOI21_X1 _28418_ (.A(_05101_),
    .B1(_06034_),
    .B2(_18332_),
    .ZN(_06035_));
 AOI22_X1 _28419_ (.A1(_05391_),
    .A2(_05768_),
    .B1(_06027_),
    .B2(_06035_),
    .ZN(_00621_));
 NOR2_X1 _28420_ (.A1(\core.dec_block.block_w1_reg[30] ),
    .A2(_05875_),
    .ZN(_06036_));
 XNOR2_X2 _28421_ (.A(_05386_),
    .B(_05537_),
    .ZN(_06037_));
 XNOR2_X1 _28422_ (.A(_05363_),
    .B(_06037_),
    .ZN(_06038_));
 XOR2_X1 _28423_ (.A(_17079_),
    .B(_03596_),
    .Z(_06039_));
 XNOR2_X1 _28424_ (.A(_05540_),
    .B(_06039_),
    .ZN(_06040_));
 XNOR2_X1 _28425_ (.A(_05597_),
    .B(_06040_),
    .ZN(_06041_));
 XNOR2_X1 _28426_ (.A(_16980_),
    .B(_06041_),
    .ZN(_06042_));
 XNOR2_X1 _28427_ (.A(_06038_),
    .B(_06042_),
    .ZN(_06043_));
 NAND2_X1 _28428_ (.A1(_18333_),
    .A2(_06043_),
    .ZN(_06044_));
 XNOR2_X1 _28429_ (.A(\block_reg[1][30] ),
    .B(_03540_),
    .ZN(_06045_));
 OAI22_X1 _28430_ (.A1(_18399_),
    .A2(_03541_),
    .B1(_06045_),
    .B2(_18412_),
    .ZN(_06046_));
 NOR3_X1 _28431_ (.A1(_05227_),
    .A2(_05768_),
    .A3(_06046_),
    .ZN(_06047_));
 AOI21_X1 _28432_ (.A(_06036_),
    .B1(_06044_),
    .B2(_06047_),
    .ZN(_00622_));
 NOR2_X1 _28433_ (.A1(\core.dec_block.block_w1_reg[31] ),
    .A2(_05875_),
    .ZN(_06048_));
 XOR2_X2 _28434_ (.A(\block_reg[1][31] ),
    .B(_17168_),
    .Z(_06049_));
 OAI221_X1 _28435_ (.A(_05259_),
    .B1(_06049_),
    .B2(_05961_),
    .C1(_17169_),
    .C2(_05902_),
    .ZN(_06050_));
 XNOR2_X2 _28436_ (.A(_16978_),
    .B(_03627_),
    .ZN(_06051_));
 XNOR2_X1 _28437_ (.A(_17062_),
    .B(_06051_),
    .ZN(_06052_));
 XOR2_X1 _28438_ (.A(_17185_),
    .B(_05590_),
    .Z(_06053_));
 XNOR2_X1 _28439_ (.A(_05491_),
    .B(_06053_),
    .ZN(_06054_));
 XNOR2_X1 _28440_ (.A(_05679_),
    .B(_06054_),
    .ZN(_06055_));
 XNOR2_X1 _28441_ (.A(_06052_),
    .B(_06055_),
    .ZN(_06056_));
 AOI21_X1 _28442_ (.A(_06050_),
    .B1(_06056_),
    .B2(_05921_),
    .ZN(_06057_));
 AOI21_X1 _28443_ (.A(_06048_),
    .B1(_06057_),
    .B2(_05784_),
    .ZN(_00623_));
 INV_X1 _28444_ (.A(\block_reg[2][3] ),
    .ZN(_06058_));
 XNOR2_X1 _28445_ (.A(_06058_),
    .B(_17861_),
    .ZN(_06059_));
 OAI221_X1 _28446_ (.A(_05847_),
    .B1(_06059_),
    .B2(_04266_),
    .C1(_05539_),
    .C2(_05021_),
    .ZN(_06060_));
 XNOR2_X1 _28447_ (.A(_17673_),
    .B(_18260_),
    .ZN(_06061_));
 XNOR2_X2 _28448_ (.A(_17780_),
    .B(_06061_),
    .ZN(_06062_));
 XNOR2_X2 _28449_ (.A(_17950_),
    .B(_06062_),
    .ZN(_06063_));
 XNOR2_X1 _28450_ (.A(_17592_),
    .B(_17935_),
    .ZN(_06064_));
 XNOR2_X1 _28451_ (.A(_17811_),
    .B(_18267_),
    .ZN(_06065_));
 XNOR2_X1 _28452_ (.A(_06064_),
    .B(_06065_),
    .ZN(_06066_));
 XNOR2_X1 _28453_ (.A(_17850_),
    .B(_06066_),
    .ZN(_06067_));
 XNOR2_X1 _28454_ (.A(_17536_),
    .B(_06067_),
    .ZN(_06068_));
 XNOR2_X2 _28455_ (.A(_06063_),
    .B(_06068_),
    .ZN(_06069_));
 OAI21_X1 _28456_ (.A(_05344_),
    .B1(_06069_),
    .B2(_17204_),
    .ZN(_06070_));
 OAI22_X1 _28457_ (.A1(\core.dec_block.block_w1_reg[3] ),
    .A2(_05784_),
    .B1(_06060_),
    .B2(_06070_),
    .ZN(_06071_));
 INV_X1 _28458_ (.A(_06071_),
    .ZN(_00624_));
 XNOR2_X1 _28459_ (.A(\block_reg[2][4] ),
    .B(_18281_),
    .ZN(_06072_));
 AOI21_X1 _28460_ (.A(_05768_),
    .B1(_06072_),
    .B2(_16372_),
    .ZN(_06073_));
 XNOR2_X2 _28461_ (.A(_17574_),
    .B(_17891_),
    .ZN(_06074_));
 XNOR2_X1 _28462_ (.A(_18259_),
    .B(_06074_),
    .ZN(_06075_));
 XNOR2_X1 _28463_ (.A(_18560_),
    .B(_06075_),
    .ZN(_06076_));
 XNOR2_X2 _28464_ (.A(_18247_),
    .B(_06076_),
    .ZN(_06077_));
 XNOR2_X2 _28465_ (.A(_18334_),
    .B(_06077_),
    .ZN(_06078_));
 XOR2_X2 _28466_ (.A(_17922_),
    .B(_18338_),
    .Z(_06079_));
 XNOR2_X2 _28467_ (.A(_18265_),
    .B(_06079_),
    .ZN(_06080_));
 XNOR2_X1 _28468_ (.A(_18283_),
    .B(_18311_),
    .ZN(_06081_));
 XNOR2_X1 _28469_ (.A(_06080_),
    .B(_06081_),
    .ZN(_06082_));
 XNOR2_X1 _28470_ (.A(_06078_),
    .B(_06082_),
    .ZN(_06083_));
 OAI221_X1 _28471_ (.A(_06073_),
    .B1(_06083_),
    .B2(_05793_),
    .C1(_16556_),
    .C2(_05590_),
    .ZN(_06084_));
 OAI22_X1 _28472_ (.A1(\core.dec_block.block_w1_reg[4] ),
    .A2(_05784_),
    .B1(_06084_),
    .B2(_05477_),
    .ZN(_06085_));
 INV_X1 _28473_ (.A(_06085_),
    .ZN(_00625_));
 NOR2_X1 _28474_ (.A1(\core.dec_block.block_w1_reg[5] ),
    .A2(_05875_),
    .ZN(_06086_));
 XNOR2_X2 _28475_ (.A(\block_reg[2][5] ),
    .B(_17760_),
    .ZN(_06087_));
 OAI221_X1 _28476_ (.A(_05772_),
    .B1(_06087_),
    .B2(_05961_),
    .C1(_17198_),
    .C2(_05902_),
    .ZN(_06088_));
 XOR2_X1 _28477_ (.A(_18482_),
    .B(_18557_),
    .Z(_06089_));
 XNOR2_X1 _28478_ (.A(_05719_),
    .B(_06089_),
    .ZN(_06090_));
 XNOR2_X1 _28479_ (.A(_18284_),
    .B(_06090_),
    .ZN(_06091_));
 XOR2_X1 _28480_ (.A(_18245_),
    .B(_18334_),
    .Z(_06092_));
 XNOR2_X1 _28481_ (.A(_06091_),
    .B(_06092_),
    .ZN(_06093_));
 AOI21_X1 _28482_ (.A(_06088_),
    .B1(_06093_),
    .B2(_05921_),
    .ZN(_06094_));
 AOI21_X1 _28483_ (.A(_06086_),
    .B1(_06094_),
    .B2(_05589_),
    .ZN(_00626_));
 NOR2_X1 _28484_ (.A1(\core.dec_block.block_w1_reg[6] ),
    .A2(_05847_),
    .ZN(_06095_));
 XNOR2_X1 _28485_ (.A(\block_reg[2][6] ),
    .B(_17657_),
    .ZN(_06096_));
 OAI221_X1 _28486_ (.A(_05772_),
    .B1(_06096_),
    .B2(_05961_),
    .C1(_16875_),
    .C2(_05902_),
    .ZN(_06097_));
 XNOR2_X2 _28487_ (.A(_17811_),
    .B(_18555_),
    .ZN(_06098_));
 XNOR2_X1 _28488_ (.A(_18343_),
    .B(_06098_),
    .ZN(_06099_));
 XOR2_X1 _28489_ (.A(_17604_),
    .B(_06031_),
    .Z(_06100_));
 XNOR2_X1 _28490_ (.A(_18284_),
    .B(_06100_),
    .ZN(_06101_));
 XNOR2_X1 _28491_ (.A(_06099_),
    .B(_06101_),
    .ZN(_06102_));
 XNOR2_X2 _28492_ (.A(_18481_),
    .B(_06102_),
    .ZN(_06103_));
 AOI21_X1 _28493_ (.A(_06097_),
    .B1(_06103_),
    .B2(_05921_),
    .ZN(_06104_));
 AOI21_X1 _28494_ (.A(_06095_),
    .B1(_06104_),
    .B2(_05650_),
    .ZN(_00627_));
 INV_X1 _28495_ (.A(\block_reg[2][7] ),
    .ZN(_06105_));
 XNOR2_X1 _28496_ (.A(_06105_),
    .B(_17517_),
    .ZN(_06106_));
 OAI221_X1 _28497_ (.A(_05771_),
    .B1(_06106_),
    .B2(_05774_),
    .C1(_17185_),
    .C2(_04264_),
    .ZN(_06107_));
 XOR2_X2 _28498_ (.A(_17658_),
    .B(_18489_),
    .Z(_06108_));
 XNOR2_X1 _28499_ (.A(_18555_),
    .B(_05721_),
    .ZN(_06109_));
 XNOR2_X2 _28500_ (.A(_06108_),
    .B(_06109_),
    .ZN(_06110_));
 XNOR2_X2 _28501_ (.A(_18340_),
    .B(_06110_),
    .ZN(_06111_));
 AOI21_X1 _28502_ (.A(_06107_),
    .B1(_06111_),
    .B2(_05782_),
    .ZN(_06112_));
 AOI22_X1 _28503_ (.A1(_17170_),
    .A2(_05768_),
    .B1(_06112_),
    .B2(_05674_),
    .ZN(_00628_));
 XNOR2_X1 _28504_ (.A(\block_reg[3][8] ),
    .B(_19015_),
    .ZN(_06113_));
 OAI221_X1 _28505_ (.A(_05771_),
    .B1(_06113_),
    .B2(_05774_),
    .C1(_17012_),
    .C2(_04264_),
    .ZN(_06114_));
 XOR2_X1 _28506_ (.A(_19027_),
    .B(_19224_),
    .Z(_06115_));
 XNOR2_X1 _28507_ (.A(_03925_),
    .B(_06115_),
    .ZN(_06116_));
 XNOR2_X1 _28508_ (.A(_19262_),
    .B(_06116_),
    .ZN(_06117_));
 XNOR2_X2 _28509_ (.A(_03301_),
    .B(_06117_),
    .ZN(_06118_));
 AOI21_X1 _28510_ (.A(_06114_),
    .B1(_06118_),
    .B2(_05782_),
    .ZN(_06119_));
 AOI22_X1 _28511_ (.A1(_16981_),
    .A2(_05768_),
    .B1(_06119_),
    .B2(_05715_),
    .ZN(_00629_));
 XNOR2_X2 _28512_ (.A(\block_reg[3][9] ),
    .B(_19273_),
    .ZN(_06120_));
 AOI21_X1 _28513_ (.A(_05767_),
    .B1(_06120_),
    .B2(_16372_),
    .ZN(_06121_));
 XNOR2_X2 _28514_ (.A(_18923_),
    .B(_03302_),
    .ZN(_06122_));
 XOR2_X1 _28515_ (.A(_18970_),
    .B(_19002_),
    .Z(_06123_));
 XOR2_X1 _28516_ (.A(_19300_),
    .B(_19445_),
    .Z(_06124_));
 XNOR2_X1 _28517_ (.A(_05798_),
    .B(_06124_),
    .ZN(_06125_));
 XNOR2_X1 _28518_ (.A(_06123_),
    .B(_06125_),
    .ZN(_06126_));
 XNOR2_X2 _28519_ (.A(_06122_),
    .B(_06126_),
    .ZN(_06127_));
 OAI221_X1 _28520_ (.A(_06121_),
    .B1(_06127_),
    .B2(_05793_),
    .C1(_03575_),
    .C2(_05021_),
    .ZN(_06128_));
 OAI22_X1 _28521_ (.A1(\core.dec_block.block_w1_reg[9] ),
    .A2(_05784_),
    .B1(_06128_),
    .B2(_05754_),
    .ZN(_06129_));
 INV_X1 _28522_ (.A(_06129_),
    .ZN(_00630_));
 AOI21_X1 _28523_ (.A(_16354_),
    .B1(_18569_),
    .B2(_16360_),
    .ZN(_06130_));
 NOR2_X1 _28524_ (.A1(_16258_),
    .A2(_06130_),
    .ZN(_06131_));
 OR2_X1 _28525_ (.A1(_16353_),
    .A2(_06131_),
    .ZN(_06132_));
 CLKBUF_X3 _28526_ (.A(_06132_),
    .Z(_06133_));
 BUF_X4 _28527_ (.A(_06133_),
    .Z(_06134_));
 BUF_X4 _28528_ (.A(_06134_),
    .Z(_06135_));
 BUF_X4 _28529_ (.A(_06133_),
    .Z(_06136_));
 XNOR2_X1 _28530_ (.A(\block_reg[3][0] ),
    .B(_19026_),
    .ZN(_06137_));
 OAI221_X2 _28531_ (.A(_06136_),
    .B1(_06137_),
    .B2(_04266_),
    .C1(_17779_),
    .C2(_05021_),
    .ZN(_06138_));
 XNOR2_X1 _28532_ (.A(_03301_),
    .B(_06122_),
    .ZN(_06139_));
 XNOR2_X1 _28533_ (.A(_19441_),
    .B(_06139_),
    .ZN(_06140_));
 OAI21_X1 _28534_ (.A(_16851_),
    .B1(_06140_),
    .B2(_17504_),
    .ZN(_06141_));
 OAI22_X1 _28535_ (.A1(\core.dec_block.block_w2_reg[0] ),
    .A2(_06135_),
    .B1(_06138_),
    .B2(_06141_),
    .ZN(_06142_));
 INV_X1 _28536_ (.A(_06142_),
    .ZN(_00631_));
 XOR2_X1 _28537_ (.A(_03510_),
    .B(_04679_),
    .Z(_06143_));
 XNOR2_X1 _28538_ (.A(_04809_),
    .B(_06143_),
    .ZN(_06144_));
 XNOR2_X1 _28539_ (.A(_04728_),
    .B(_06144_),
    .ZN(_06145_));
 NOR2_X1 _28540_ (.A1(_17504_),
    .A2(_06145_),
    .ZN(_06146_));
 XNOR2_X1 _28541_ (.A(\block_reg[0][10] ),
    .B(_17739_),
    .ZN(_06147_));
 OAI221_X1 _28542_ (.A(_06134_),
    .B1(_06147_),
    .B2(_18078_),
    .C1(_17865_),
    .C2(_17741_),
    .ZN(_06148_));
 NOR3_X1 _28543_ (.A1(_17503_),
    .A2(_06146_),
    .A3(_06148_),
    .ZN(_06149_));
 NOR2_X2 _28544_ (.A1(_16353_),
    .A2(_06131_),
    .ZN(_06150_));
 BUF_X4 _28545_ (.A(_06150_),
    .Z(_06151_));
 BUF_X4 _28546_ (.A(_06151_),
    .Z(_06152_));
 AOI21_X1 _28547_ (.A(_06149_),
    .B1(_06152_),
    .B2(_17864_),
    .ZN(_00632_));
 XOR2_X1 _28548_ (.A(_17740_),
    .B(_05184_),
    .Z(_06153_));
 XNOR2_X1 _28549_ (.A(_05008_),
    .B(_06153_),
    .ZN(_06154_));
 XNOR2_X1 _28550_ (.A(_04818_),
    .B(_06154_),
    .ZN(_06155_));
 NAND2_X1 _28551_ (.A1(_17749_),
    .A2(_06155_),
    .ZN(_06156_));
 XOR2_X1 _28552_ (.A(\block_reg[0][11] ),
    .B(_18063_),
    .Z(_06157_));
 OAI22_X1 _28553_ (.A1(_17741_),
    .A2(_18267_),
    .B1(_06157_),
    .B2(_18078_),
    .ZN(_06158_));
 NOR3_X1 _28554_ (.A1(_18051_),
    .A2(_06151_),
    .A3(_06158_),
    .ZN(_06159_));
 AOI22_X1 _28555_ (.A1(_18266_),
    .A2(_06152_),
    .B1(_06156_),
    .B2(_06159_),
    .ZN(_00633_));
 INV_X1 _28556_ (.A(\block_reg[0][12] ),
    .ZN(_06160_));
 XNOR2_X1 _28557_ (.A(_06160_),
    .B(_18325_),
    .ZN(_06161_));
 AOI21_X1 _28558_ (.A(_06151_),
    .B1(_06161_),
    .B2(_16371_),
    .ZN(_06162_));
 XOR2_X1 _28559_ (.A(_05016_),
    .B(_05938_),
    .Z(_06163_));
 XNOR2_X1 _28560_ (.A(_04940_),
    .B(_06163_),
    .ZN(_06164_));
 XNOR2_X1 _28561_ (.A(_05918_),
    .B(_06164_),
    .ZN(_06165_));
 OAI221_X1 _28562_ (.A(_06162_),
    .B1(_06165_),
    .B2(_05793_),
    .C1(_16556_),
    .C2(_18337_),
    .ZN(_06166_));
 OAI22_X1 _28563_ (.A1(\core.dec_block.block_w2_reg[12] ),
    .A2(_06135_),
    .B1(_06166_),
    .B2(_18228_),
    .ZN(_06167_));
 INV_X1 _28564_ (.A(_06167_),
    .ZN(_00634_));
 NOR2_X1 _28565_ (.A1(\core.dec_block.block_w2_reg[13] ),
    .A2(_06135_),
    .ZN(_06168_));
 XOR2_X1 _28566_ (.A(_05188_),
    .B(_05262_),
    .Z(_06169_));
 XNOR2_X1 _28567_ (.A(_05014_),
    .B(_06169_),
    .ZN(_06170_));
 NAND2_X1 _28568_ (.A1(_18333_),
    .A2(_06170_),
    .ZN(_06171_));
 XNOR2_X1 _28569_ (.A(\block_reg[0][13] ),
    .B(_18409_),
    .ZN(_06172_));
 OAI22_X1 _28570_ (.A1(_18399_),
    .A2(_17824_),
    .B1(_06172_),
    .B2(_18412_),
    .ZN(_06173_));
 NOR3_X1 _28571_ (.A1(_18398_),
    .A2(_06151_),
    .A3(_06173_),
    .ZN(_06174_));
 AOI21_X1 _28572_ (.A(_06168_),
    .B1(_06171_),
    .B2(_06174_),
    .ZN(_00635_));
 NOR2_X1 _28573_ (.A1(\core.dec_block.block_w2_reg[14] ),
    .A2(_06135_),
    .ZN(_06175_));
 XNOR2_X1 _28574_ (.A(\block_reg[0][14] ),
    .B(_18477_),
    .ZN(_06176_));
 OAI221_X2 _28575_ (.A(_06136_),
    .B1(_06176_),
    .B2(_05961_),
    .C1(_17702_),
    .C2(_05902_),
    .ZN(_06177_));
 XNOR2_X1 _28576_ (.A(_03915_),
    .B(_04723_),
    .ZN(_06178_));
 XNOR2_X1 _28577_ (.A(_04919_),
    .B(_06178_),
    .ZN(_06179_));
 XNOR2_X1 _28578_ (.A(_05007_),
    .B(_06179_),
    .ZN(_06180_));
 XNOR2_X1 _28579_ (.A(_05187_),
    .B(_06180_),
    .ZN(_06181_));
 AOI21_X1 _28580_ (.A(_06177_),
    .B1(_06181_),
    .B2(_05921_),
    .ZN(_06182_));
 AOI21_X1 _28581_ (.A(_06175_),
    .B1(_06182_),
    .B2(_18465_),
    .ZN(_00636_));
 NOR2_X1 _28582_ (.A1(\core.dec_block.block_w2_reg[15] ),
    .A2(_06135_),
    .ZN(_06183_));
 XNOR2_X2 _28583_ (.A(\block_reg[0][15] ),
    .B(_18549_),
    .ZN(_06184_));
 OAI221_X2 _28584_ (.A(_06136_),
    .B1(_06184_),
    .B2(_05961_),
    .C1(_17848_),
    .C2(_05902_),
    .ZN(_06185_));
 XOR2_X1 _28585_ (.A(_03976_),
    .B(_04289_),
    .Z(_06186_));
 XNOR2_X1 _28586_ (.A(_04937_),
    .B(_06186_),
    .ZN(_06187_));
 XNOR2_X1 _28587_ (.A(_05950_),
    .B(_06187_),
    .ZN(_06188_));
 XNOR2_X1 _28588_ (.A(_05930_),
    .B(_06188_),
    .ZN(_06189_));
 AOI21_X1 _28589_ (.A(_06185_),
    .B1(_06189_),
    .B2(_05921_),
    .ZN(_06190_));
 AOI21_X1 _28590_ (.A(_06183_),
    .B1(_06190_),
    .B2(_18526_),
    .ZN(_00637_));
 XNOR2_X1 _28591_ (.A(\block_reg[1][16] ),
    .B(_17138_),
    .ZN(_06191_));
 OAI221_X2 _28592_ (.A(_06133_),
    .B1(_06191_),
    .B2(_05774_),
    .C1(_17906_),
    .C2(_04264_),
    .ZN(_06192_));
 XOR2_X1 _28593_ (.A(_03527_),
    .B(_05971_),
    .Z(_06193_));
 XNOR2_X1 _28594_ (.A(_17064_),
    .B(_06193_),
    .ZN(_06194_));
 AOI21_X1 _28595_ (.A(_06192_),
    .B1(_06194_),
    .B2(_05782_),
    .ZN(_06195_));
 AOI22_X1 _28596_ (.A1(_17892_),
    .A2(_06152_),
    .B1(_06195_),
    .B2(_18848_),
    .ZN(_00638_));
 NOR2_X1 _28597_ (.A1(\core.dec_block.block_w2_reg[17] ),
    .A2(_06135_),
    .ZN(_06196_));
 INV_X1 _28598_ (.A(\block_reg[1][17] ),
    .ZN(_06197_));
 XNOR2_X1 _28599_ (.A(_06197_),
    .B(_03615_),
    .ZN(_06198_));
 BUF_X4 _28600_ (.A(_16555_),
    .Z(_06199_));
 OAI221_X2 _28601_ (.A(_06136_),
    .B1(_06198_),
    .B2(_05961_),
    .C1(_18259_),
    .C2(_06199_),
    .ZN(_06200_));
 XNOR2_X1 _28602_ (.A(_05115_),
    .B(_05177_),
    .ZN(_06201_));
 XNOR2_X1 _28603_ (.A(_05995_),
    .B(_06201_),
    .ZN(_06202_));
 XNOR2_X1 _28604_ (.A(_17199_),
    .B(_06202_),
    .ZN(_06203_));
 XNOR2_X1 _28605_ (.A(_05494_),
    .B(_06203_),
    .ZN(_06204_));
 AOI21_X1 _28606_ (.A(_06200_),
    .B1(_06204_),
    .B2(_05921_),
    .ZN(_06205_));
 AOI21_X1 _28607_ (.A(_06196_),
    .B1(_06205_),
    .B2(_19179_),
    .ZN(_00639_));
 NOR2_X1 _28608_ (.A1(\core.dec_block.block_w2_reg[18] ),
    .A2(_06135_),
    .ZN(_06206_));
 XNOR2_X1 _28609_ (.A(\block_reg[1][18] ),
    .B(_05175_),
    .ZN(_06207_));
 OAI221_X2 _28610_ (.A(_06136_),
    .B1(_06207_),
    .B2(_05961_),
    .C1(_17563_),
    .C2(_06199_),
    .ZN(_06208_));
 XOR2_X1 _28611_ (.A(_03575_),
    .B(_03616_),
    .Z(_06209_));
 XNOR2_X1 _28612_ (.A(_06017_),
    .B(_06209_),
    .ZN(_06210_));
 XNOR2_X1 _28613_ (.A(_05164_),
    .B(_06210_),
    .ZN(_06211_));
 BUF_X4 _28614_ (.A(_17748_),
    .Z(_06212_));
 AOI21_X1 _28615_ (.A(_06208_),
    .B1(_06211_),
    .B2(_06212_),
    .ZN(_06213_));
 AOI21_X1 _28616_ (.A(_06206_),
    .B1(_06213_),
    .B2(_19371_),
    .ZN(_00640_));
 XNOR2_X1 _28617_ (.A(\block_reg[1][19] ),
    .B(_05405_),
    .ZN(_06214_));
 AOI21_X1 _28618_ (.A(_06150_),
    .B1(_06214_),
    .B2(_16371_),
    .ZN(_06215_));
 OAI21_X1 _28619_ (.A(_06215_),
    .B1(_17811_),
    .B2(_18052_),
    .ZN(_06216_));
 XNOR2_X1 _28620_ (.A(_05115_),
    .B(_05539_),
    .ZN(_06217_));
 XNOR2_X2 _28621_ (.A(_05158_),
    .B(_06217_),
    .ZN(_06218_));
 XNOR2_X1 _28622_ (.A(_05592_),
    .B(_06218_),
    .ZN(_06219_));
 XNOR2_X1 _28623_ (.A(_05390_),
    .B(_06219_),
    .ZN(_06220_));
 AOI21_X1 _28624_ (.A(_06216_),
    .B1(_06220_),
    .B2(_05782_),
    .ZN(_06221_));
 AOI22_X1 _28625_ (.A1(_17799_),
    .A2(_06152_),
    .B1(_06221_),
    .B2(_19519_),
    .ZN(_00641_));
 BUF_X4 _28626_ (.A(_06134_),
    .Z(_06222_));
 NOR2_X1 _28627_ (.A1(\core.dec_block.block_w2_reg[1] ),
    .A2(_06222_),
    .ZN(_06223_));
 XNOR2_X2 _28628_ (.A(\block_reg[3][1] ),
    .B(_19284_),
    .ZN(_06224_));
 BUF_X4 _28629_ (.A(_17709_),
    .Z(_06225_));
 OAI221_X2 _28630_ (.A(_03498_),
    .B1(_06224_),
    .B2(_06225_),
    .C1(_17672_),
    .C2(_06199_),
    .ZN(_06226_));
 XNOR2_X1 _28631_ (.A(_18896_),
    .B(_18956_),
    .ZN(_06227_));
 XNOR2_X1 _28632_ (.A(_05798_),
    .B(_06227_),
    .ZN(_06228_));
 XOR2_X1 _28633_ (.A(_19003_),
    .B(_06228_),
    .Z(_06229_));
 XNOR2_X1 _28634_ (.A(_19299_),
    .B(_19446_),
    .ZN(_06230_));
 XNOR2_X1 _28635_ (.A(_03926_),
    .B(_06230_),
    .ZN(_06231_));
 XNOR2_X1 _28636_ (.A(_06229_),
    .B(_06231_),
    .ZN(_06232_));
 AOI21_X1 _28637_ (.A(_06226_),
    .B1(_06232_),
    .B2(_06212_),
    .ZN(_06233_));
 AOI21_X1 _28638_ (.A(_06223_),
    .B1(_06233_),
    .B2(_06135_),
    .ZN(_00642_));
 XNOR2_X1 _28639_ (.A(\block_reg[1][20] ),
    .B(_05523_),
    .ZN(_06234_));
 OAI221_X2 _28640_ (.A(_06133_),
    .B1(_06234_),
    .B2(_05774_),
    .C1(_18297_),
    .C2(_04264_),
    .ZN(_06235_));
 XNOR2_X1 _28641_ (.A(_17199_),
    .B(_05590_),
    .ZN(_06236_));
 XNOR2_X1 _28642_ (.A(_06037_),
    .B(_06236_),
    .ZN(_06237_));
 XNOR2_X1 _28643_ (.A(_05597_),
    .B(_06237_),
    .ZN(_06238_));
 XNOR2_X1 _28644_ (.A(_05498_),
    .B(_06238_),
    .ZN(_06239_));
 AOI21_X1 _28645_ (.A(_06235_),
    .B1(_06239_),
    .B2(_05782_),
    .ZN(_06240_));
 AOI22_X1 _28646_ (.A1(_18285_),
    .A2(_06152_),
    .B1(_06240_),
    .B2(_03698_),
    .ZN(_00643_));
 NOR2_X1 _28647_ (.A1(\core.dec_block.block_w2_reg[21] ),
    .A2(_06222_),
    .ZN(_06241_));
 XOR2_X1 _28648_ (.A(\block_reg[1][21] ),
    .B(_16942_),
    .Z(_06242_));
 OAI22_X1 _28649_ (.A1(_16556_),
    .A2(_17891_),
    .B1(_06242_),
    .B2(_04266_),
    .ZN(_06243_));
 NOR2_X1 _28650_ (.A1(_06151_),
    .A2(_06243_),
    .ZN(_06244_));
 XNOR2_X1 _28651_ (.A(_05138_),
    .B(_06051_),
    .ZN(_06245_));
 XNOR2_X1 _28652_ (.A(_05538_),
    .B(_05598_),
    .ZN(_06246_));
 XNOR2_X1 _28653_ (.A(_17198_),
    .B(_05176_),
    .ZN(_06247_));
 XNOR2_X1 _28654_ (.A(_05596_),
    .B(_06247_),
    .ZN(_06248_));
 XNOR2_X1 _28655_ (.A(_06246_),
    .B(_06248_),
    .ZN(_06249_));
 XNOR2_X1 _28656_ (.A(_06245_),
    .B(_06249_),
    .ZN(_06250_));
 XOR2_X1 _28657_ (.A(_06017_),
    .B(_06218_),
    .Z(_06251_));
 XNOR2_X1 _28658_ (.A(_05963_),
    .B(_06251_),
    .ZN(_06252_));
 XNOR2_X1 _28659_ (.A(_06250_),
    .B(_06252_),
    .ZN(_06253_));
 AOI21_X1 _28660_ (.A(_03845_),
    .B1(_06253_),
    .B2(_19031_),
    .ZN(_06254_));
 AOI21_X1 _28661_ (.A(_06241_),
    .B1(_06244_),
    .B2(_06254_),
    .ZN(_00644_));
 NOR2_X1 _28662_ (.A1(\core.dec_block.block_w2_reg[22] ),
    .A2(_06222_),
    .ZN(_06255_));
 XOR2_X2 _28663_ (.A(\block_reg[1][22] ),
    .B(_16977_),
    .Z(_06256_));
 OAI221_X2 _28664_ (.A(_06136_),
    .B1(_06256_),
    .B2(_06225_),
    .C1(_17574_),
    .C2(_06199_),
    .ZN(_06257_));
 XNOR2_X1 _28665_ (.A(_05994_),
    .B(_06019_),
    .ZN(_06258_));
 XNOR2_X1 _28666_ (.A(_05963_),
    .B(_06258_),
    .ZN(_06259_));
 XOR2_X1 _28667_ (.A(_05362_),
    .B(_05591_),
    .Z(_06260_));
 XNOR2_X1 _28668_ (.A(_05540_),
    .B(_06260_),
    .ZN(_06261_));
 XNOR2_X2 _28669_ (.A(_06259_),
    .B(_06261_),
    .ZN(_06262_));
 AOI21_X1 _28670_ (.A(_06257_),
    .B1(_06262_),
    .B2(_06212_),
    .ZN(_06263_));
 AOI21_X1 _28671_ (.A(_06255_),
    .B1(_06263_),
    .B2(_03893_),
    .ZN(_00645_));
 XOR2_X2 _28672_ (.A(\block_reg[1][23] ),
    .B(_03626_),
    .Z(_06264_));
 AOI21_X2 _28673_ (.A(_06150_),
    .B1(_06264_),
    .B2(_16371_),
    .ZN(_06265_));
 XNOR2_X1 _28674_ (.A(_05613_),
    .B(_06010_),
    .ZN(_06266_));
 XNOR2_X2 _28675_ (.A(_17169_),
    .B(_05510_),
    .ZN(_06267_));
 XNOR2_X1 _28676_ (.A(_16979_),
    .B(_06267_),
    .ZN(_06268_));
 XNOR2_X2 _28677_ (.A(_06266_),
    .B(_06268_),
    .ZN(_06269_));
 OAI221_X2 _28678_ (.A(_06265_),
    .B1(_06269_),
    .B2(_05793_),
    .C1(_16556_),
    .C2(_17552_),
    .ZN(_06270_));
 OAI22_X1 _28679_ (.A1(_17537_),
    .A2(_06135_),
    .B1(_06270_),
    .B2(_03955_),
    .ZN(_06271_));
 INV_X1 _28680_ (.A(_06271_),
    .ZN(_00646_));
 NOR2_X1 _28681_ (.A1(\core.dec_block.block_w2_reg[24] ),
    .A2(_06222_),
    .ZN(_06272_));
 XNOR2_X1 _28682_ (.A(\block_reg[2][24] ),
    .B(_17642_),
    .ZN(_06273_));
 OAI221_X1 _28683_ (.A(_06136_),
    .B1(_06273_),
    .B2(_06225_),
    .C1(_17643_),
    .C2(_06199_),
    .ZN(_06274_));
 XOR2_X1 _28684_ (.A(_18560_),
    .B(_05905_),
    .Z(_06275_));
 XNOR2_X1 _28685_ (.A(_05759_),
    .B(_06275_),
    .ZN(_06276_));
 XNOR2_X1 _28686_ (.A(_17908_),
    .B(_06276_),
    .ZN(_06277_));
 AOI21_X1 _28687_ (.A(_06274_),
    .B1(_06277_),
    .B2(_06212_),
    .ZN(_06278_));
 AOI21_X1 _28688_ (.A(_06272_),
    .B1(_06278_),
    .B2(_04251_),
    .ZN(_00647_));
 NOR2_X1 _28689_ (.A1(\core.dec_block.block_w2_reg[25] ),
    .A2(_06222_),
    .ZN(_06279_));
 XNOR2_X1 _28690_ (.A(\block_reg[2][25] ),
    .B(_17795_),
    .ZN(_06280_));
 OAI221_X1 _28691_ (.A(_06136_),
    .B1(_06280_),
    .B2(_06225_),
    .C1(_17796_),
    .C2(_06199_),
    .ZN(_06281_));
 XNOR2_X1 _28692_ (.A(_17552_),
    .B(_17947_),
    .ZN(_06282_));
 XOR2_X1 _28693_ (.A(_17689_),
    .B(_17848_),
    .Z(_06283_));
 XNOR2_X1 _28694_ (.A(_17906_),
    .B(_06283_),
    .ZN(_06284_));
 XNOR2_X1 _28695_ (.A(_06282_),
    .B(_06284_),
    .ZN(_06285_));
 XNOR2_X1 _28696_ (.A(_18262_),
    .B(_18265_),
    .ZN(_06286_));
 XNOR2_X1 _28697_ (.A(_06285_),
    .B(_06286_),
    .ZN(_06287_));
 AOI21_X1 _28698_ (.A(_06281_),
    .B1(_06287_),
    .B2(_06212_),
    .ZN(_06288_));
 AOI21_X1 _28699_ (.A(_06279_),
    .B1(_06288_),
    .B2(_04538_),
    .ZN(_00648_));
 NOR2_X1 _28700_ (.A1(\core.dec_block.block_w2_reg[26] ),
    .A2(_06222_),
    .ZN(_06289_));
 OAI21_X1 _28701_ (.A(_06136_),
    .B1(_17592_),
    .B2(_05021_),
    .ZN(_06290_));
 XOR2_X1 _28702_ (.A(\block_reg[2][26] ),
    .B(_17591_),
    .Z(_06291_));
 AOI21_X1 _28703_ (.A(_06290_),
    .B1(_06291_),
    .B2(_16372_),
    .ZN(_06292_));
 XOR2_X1 _28704_ (.A(_17618_),
    .B(_17865_),
    .Z(_06293_));
 XNOR2_X1 _28705_ (.A(_05907_),
    .B(_06293_),
    .ZN(_06294_));
 XNOR2_X1 _28706_ (.A(_17797_),
    .B(_06294_),
    .ZN(_06295_));
 XNOR2_X1 _28707_ (.A(_18335_),
    .B(_06295_),
    .ZN(_06296_));
 AOI21_X1 _28708_ (.A(_04657_),
    .B1(_06296_),
    .B2(_05782_),
    .ZN(_06297_));
 AOI21_X1 _28709_ (.A(_06289_),
    .B1(_06292_),
    .B2(_06297_),
    .ZN(_00649_));
 XOR2_X1 _28710_ (.A(\block_reg[2][27] ),
    .B(_17921_),
    .Z(_06298_));
 OAI221_X1 _28711_ (.A(_06134_),
    .B1(_06298_),
    .B2(_18078_),
    .C1(_17922_),
    .C2(_18052_),
    .ZN(_06299_));
 XNOR2_X1 _28712_ (.A(_17907_),
    .B(_17947_),
    .ZN(_06300_));
 XNOR2_X1 _28713_ (.A(_17592_),
    .B(_06300_),
    .ZN(_06301_));
 XNOR2_X1 _28714_ (.A(_17563_),
    .B(_18267_),
    .ZN(_06302_));
 XNOR2_X1 _28715_ (.A(_17863_),
    .B(_06302_),
    .ZN(_06303_));
 XNOR2_X1 _28716_ (.A(_06301_),
    .B(_06303_),
    .ZN(_06304_));
 XNOR2_X1 _28717_ (.A(_17813_),
    .B(_06304_),
    .ZN(_06305_));
 NOR2_X1 _28718_ (.A1(_05793_),
    .A2(_06305_),
    .ZN(_06306_));
 NOR3_X1 _28719_ (.A1(_04792_),
    .A2(_06299_),
    .A3(_06306_),
    .ZN(_06307_));
 AOI21_X1 _28720_ (.A(_06307_),
    .B1(_06152_),
    .B2(_17909_),
    .ZN(_00650_));
 NOR2_X1 _28721_ (.A1(\core.dec_block.block_w2_reg[28] ),
    .A2(_06222_),
    .ZN(_06308_));
 XNOR2_X1 _28722_ (.A(\block_reg[2][28] ),
    .B(_18309_),
    .ZN(_06309_));
 OAI221_X1 _28723_ (.A(_06134_),
    .B1(_06309_),
    .B2(_06225_),
    .C1(_18310_),
    .C2(_06199_),
    .ZN(_06310_));
 XNOR2_X1 _28724_ (.A(_18282_),
    .B(_06098_),
    .ZN(_06311_));
 XNOR2_X2 _28725_ (.A(_06080_),
    .B(_06311_),
    .ZN(_06312_));
 XNOR2_X2 _28726_ (.A(_18264_),
    .B(_06312_),
    .ZN(_06313_));
 AOI21_X1 _28727_ (.A(_06310_),
    .B1(_06313_),
    .B2(_06212_),
    .ZN(_06314_));
 AOI21_X1 _28728_ (.A(_06308_),
    .B1(_06314_),
    .B2(_04902_),
    .ZN(_00651_));
 NOR2_X1 _28729_ (.A1(\core.dec_block.block_w2_reg[29] ),
    .A2(_06222_),
    .ZN(_06315_));
 XOR2_X1 _28730_ (.A(_17761_),
    .B(_18261_),
    .Z(_06316_));
 XNOR2_X1 _28731_ (.A(_18311_),
    .B(_06316_),
    .ZN(_06317_));
 XNOR2_X1 _28732_ (.A(_18481_),
    .B(_06317_),
    .ZN(_06318_));
 XNOR2_X1 _28733_ (.A(_18336_),
    .B(_06318_),
    .ZN(_06319_));
 NAND2_X1 _28734_ (.A1(_18333_),
    .A2(_06319_),
    .ZN(_06320_));
 XNOR2_X1 _28735_ (.A(\block_reg[2][29] ),
    .B(_17945_),
    .ZN(_06321_));
 OAI22_X1 _28736_ (.A1(_18399_),
    .A2(_17946_),
    .B1(_06321_),
    .B2(_18466_),
    .ZN(_06322_));
 NOR3_X1 _28737_ (.A1(_05003_),
    .A2(_06151_),
    .A3(_06322_),
    .ZN(_06323_));
 AOI21_X1 _28738_ (.A(_06315_),
    .B1(_06320_),
    .B2(_06323_),
    .ZN(_00652_));
 XNOR2_X1 _28739_ (.A(\block_reg[3][2] ),
    .B(_19457_),
    .ZN(_06324_));
 OAI22_X1 _28740_ (.A1(_03858_),
    .A2(_17535_),
    .B1(_06324_),
    .B2(_18553_),
    .ZN(_06325_));
 NOR2_X1 _28741_ (.A1(_06151_),
    .A2(_06325_),
    .ZN(_06326_));
 XOR2_X1 _28742_ (.A(_19300_),
    .B(_03332_),
    .Z(_06327_));
 XNOR2_X1 _28743_ (.A(_19444_),
    .B(_06327_),
    .ZN(_06328_));
 AOI21_X1 _28744_ (.A(_05101_),
    .B1(_06328_),
    .B2(_18332_),
    .ZN(_06329_));
 AOI22_X1 _28745_ (.A1(_17519_),
    .A2(_06152_),
    .B1(_06326_),
    .B2(_06329_),
    .ZN(_00653_));
 XOR2_X1 _28746_ (.A(_17702_),
    .B(_18337_),
    .Z(_06330_));
 XNOR2_X1 _28747_ (.A(_06074_),
    .B(_06330_),
    .ZN(_06331_));
 XNOR2_X1 _28748_ (.A(_18557_),
    .B(_06331_),
    .ZN(_06332_));
 XNOR2_X1 _28749_ (.A(_18485_),
    .B(_06332_),
    .ZN(_06333_));
 NOR2_X1 _28750_ (.A1(_05793_),
    .A2(_06333_),
    .ZN(_06334_));
 XNOR2_X2 _28751_ (.A(\block_reg[2][30] ),
    .B(_17603_),
    .ZN(_06335_));
 OAI221_X1 _28752_ (.A(_06134_),
    .B1(_06335_),
    .B2(_18078_),
    .C1(_17604_),
    .C2(_04264_),
    .ZN(_06336_));
 NOR3_X1 _28753_ (.A1(_05227_),
    .A2(_06334_),
    .A3(_06336_),
    .ZN(_06337_));
 INV_X1 _28754_ (.A(\core.dec_block.block_w2_reg[30] ),
    .ZN(_06338_));
 AOI21_X1 _28755_ (.A(_06337_),
    .B1(_06152_),
    .B2(_06338_),
    .ZN(_00654_));
 XOR2_X2 _28756_ (.A(\block_reg[2][31] ),
    .B(_17934_),
    .Z(_06339_));
 OAI221_X1 _28757_ (.A(_06133_),
    .B1(_06339_),
    .B2(_05774_),
    .C1(_17935_),
    .C2(_04264_),
    .ZN(_06340_));
 XOR2_X2 _28758_ (.A(_18488_),
    .B(_05721_),
    .Z(_06341_));
 XNOR2_X2 _28759_ (.A(_18559_),
    .B(_06341_),
    .ZN(_06342_));
 AOI21_X1 _28760_ (.A(_06340_),
    .B1(_06342_),
    .B2(_18332_),
    .ZN(_06343_));
 AOI22_X1 _28761_ (.A1(_17923_),
    .A2(_06152_),
    .B1(_06343_),
    .B2(_05259_),
    .ZN(_00655_));
 XNOR2_X1 _28762_ (.A(\block_reg[3][3] ),
    .B(_03357_),
    .ZN(_06344_));
 OAI221_X1 _28763_ (.A(_06136_),
    .B1(_06344_),
    .B2(_04266_),
    .C1(_17862_),
    .C2(_05021_),
    .ZN(_06345_));
 XNOR2_X1 _28764_ (.A(_19429_),
    .B(_05798_),
    .ZN(_06346_));
 XNOR2_X1 _28765_ (.A(_03919_),
    .B(_06346_),
    .ZN(_06347_));
 XNOR2_X1 _28766_ (.A(_03791_),
    .B(_06347_),
    .ZN(_06348_));
 XNOR2_X1 _28767_ (.A(_03331_),
    .B(_06348_),
    .ZN(_06349_));
 OAI21_X1 _28768_ (.A(_05344_),
    .B1(_06349_),
    .B2(_17504_),
    .ZN(_06350_));
 OAI22_X1 _28769_ (.A1(\core.dec_block.block_w2_reg[3] ),
    .A2(_06135_),
    .B1(_06345_),
    .B2(_06350_),
    .ZN(_06351_));
 INV_X1 _28770_ (.A(_06351_),
    .ZN(_00656_));
 XNOR2_X1 _28771_ (.A(_19224_),
    .B(_03327_),
    .ZN(_06352_));
 XNOR2_X1 _28772_ (.A(_03783_),
    .B(_05837_),
    .ZN(_06353_));
 XNOR2_X1 _28773_ (.A(_06352_),
    .B(_06353_),
    .ZN(_06354_));
 XNOR2_X1 _28774_ (.A(_03790_),
    .B(_06354_),
    .ZN(_06355_));
 XNOR2_X1 _28775_ (.A(_03747_),
    .B(_06355_),
    .ZN(_06356_));
 NAND2_X1 _28776_ (.A1(_17749_),
    .A2(_06356_),
    .ZN(_06357_));
 XNOR2_X1 _28777_ (.A(\block_reg[3][4] ),
    .B(_03759_),
    .ZN(_06358_));
 OAI221_X2 _28778_ (.A(_06134_),
    .B1(_06358_),
    .B2(_17710_),
    .C1(_18282_),
    .C2(_18052_),
    .ZN(_06359_));
 NOR2_X1 _28779_ (.A1(_05477_),
    .A2(_06359_),
    .ZN(_06360_));
 AOI22_X1 _28780_ (.A1(_18270_),
    .A2(_06151_),
    .B1(_06357_),
    .B2(_06360_),
    .ZN(_00657_));
 NOR2_X1 _28781_ (.A1(\core.dec_block.block_w2_reg[5] ),
    .A2(_06222_),
    .ZN(_06361_));
 INV_X1 _28782_ (.A(\block_reg[3][5] ),
    .ZN(_06362_));
 XNOR2_X1 _28783_ (.A(_06362_),
    .B(_18895_),
    .ZN(_06363_));
 OAI221_X2 _28784_ (.A(_06134_),
    .B1(_06363_),
    .B2(_06225_),
    .C1(_17761_),
    .C2(_06199_),
    .ZN(_06364_));
 XNOR2_X1 _28785_ (.A(_18909_),
    .B(_03739_),
    .ZN(_06365_));
 XNOR2_X1 _28786_ (.A(_19413_),
    .B(_06365_),
    .ZN(_06366_));
 XNOR2_X1 _28787_ (.A(_03761_),
    .B(_06366_),
    .ZN(_06367_));
 XNOR2_X1 _28788_ (.A(_03743_),
    .B(_06367_),
    .ZN(_06368_));
 XNOR2_X1 _28789_ (.A(_03788_),
    .B(_06368_),
    .ZN(_06369_));
 AOI21_X1 _28790_ (.A(_06364_),
    .B1(_06369_),
    .B2(_06212_),
    .ZN(_06370_));
 AOI21_X1 _28791_ (.A(_06361_),
    .B1(_06370_),
    .B2(_05589_),
    .ZN(_00658_));
 NOR2_X1 _28792_ (.A1(_16589_),
    .A2(_06222_),
    .ZN(_06371_));
 XNOR2_X1 _28793_ (.A(\block_reg[3][6] ),
    .B(_18883_),
    .ZN(_06372_));
 OAI221_X2 _28794_ (.A(_06134_),
    .B1(_06372_),
    .B2(_06225_),
    .C1(_17658_),
    .C2(_06199_),
    .ZN(_06373_));
 XOR2_X1 _28795_ (.A(_18896_),
    .B(_19247_),
    .Z(_06374_));
 XNOR2_X1 _28796_ (.A(_03327_),
    .B(_03783_),
    .ZN(_06375_));
 XNOR2_X1 _28797_ (.A(_06374_),
    .B(_06375_),
    .ZN(_06376_));
 XNOR2_X1 _28798_ (.A(_05811_),
    .B(_06376_),
    .ZN(_06377_));
 XNOR2_X1 _28799_ (.A(_05841_),
    .B(_06377_),
    .ZN(_06378_));
 AOI21_X1 _28800_ (.A(_06373_),
    .B1(_06378_),
    .B2(_06212_),
    .ZN(_06379_));
 AOI21_X1 _28801_ (.A(_06371_),
    .B1(_06379_),
    .B2(_05650_),
    .ZN(_00659_));
 XNOR2_X1 _28802_ (.A(\block_reg[3][7] ),
    .B(_19259_),
    .ZN(_06380_));
 AOI21_X1 _28803_ (.A(_06150_),
    .B1(_06380_),
    .B2(_16371_),
    .ZN(_06381_));
 OAI21_X1 _28804_ (.A(_06381_),
    .B1(_17518_),
    .B2(_18052_),
    .ZN(_06382_));
 XOR2_X2 _28805_ (.A(_18957_),
    .B(_03925_),
    .Z(_06383_));
 XNOR2_X2 _28806_ (.A(_05838_),
    .B(_06383_),
    .ZN(_06384_));
 XNOR2_X2 _28807_ (.A(_03959_),
    .B(_06384_),
    .ZN(_06385_));
 AOI21_X1 _28808_ (.A(_06382_),
    .B1(_06385_),
    .B2(_18332_),
    .ZN(_06386_));
 AOI22_X1 _28809_ (.A1(_17505_),
    .A2(_06151_),
    .B1(_06386_),
    .B2(_05674_),
    .ZN(_00660_));
 XNOR2_X1 _28810_ (.A(\block_reg[0][8] ),
    .B(_04326_),
    .ZN(_06387_));
 OAI221_X1 _28811_ (.A(_06133_),
    .B1(_06387_),
    .B2(_05774_),
    .C1(_17618_),
    .C2(_19180_),
    .ZN(_06388_));
 XOR2_X1 _28812_ (.A(_04314_),
    .B(_05870_),
    .Z(_06389_));
 XNOR2_X1 _28813_ (.A(_05859_),
    .B(_06389_),
    .ZN(_06390_));
 AOI21_X1 _28814_ (.A(_06388_),
    .B1(_06390_),
    .B2(_18332_),
    .ZN(_06391_));
 AOI22_X1 _28815_ (.A1(_17606_),
    .A2(_06151_),
    .B1(_06391_),
    .B2(_05715_),
    .ZN(_00661_));
 XNOR2_X1 _28816_ (.A(\block_reg[0][9] ),
    .B(_04563_),
    .ZN(_06392_));
 OAI221_X1 _28817_ (.A(_06134_),
    .B1(_06392_),
    .B2(_18078_),
    .C1(_17689_),
    .C2(_18052_),
    .ZN(_06393_));
 XNOR2_X2 _28818_ (.A(_04349_),
    .B(_04552_),
    .ZN(_06394_));
 XNOR2_X1 _28819_ (.A(_05188_),
    .B(_06394_),
    .ZN(_06395_));
 XNOR2_X1 _28820_ (.A(_05891_),
    .B(_06395_),
    .ZN(_06396_));
 NOR2_X1 _28821_ (.A1(_05793_),
    .A2(_06396_),
    .ZN(_06397_));
 NOR3_X1 _28822_ (.A1(_05754_),
    .A2(_06393_),
    .A3(_06397_),
    .ZN(_06398_));
 INV_X1 _28823_ (.A(\core.dec_block.block_w2_reg[9] ),
    .ZN(_06399_));
 AOI21_X1 _28824_ (.A(_06398_),
    .B1(_06152_),
    .B2(_06399_),
    .ZN(_00662_));
 OAI21_X1 _28825_ (.A(_16351_),
    .B1(_16269_),
    .B2(_16260_),
    .ZN(_06400_));
 AND2_X1 _28826_ (.A1(_16259_),
    .A2(_06400_),
    .ZN(_06401_));
 OR2_X1 _28827_ (.A1(_16353_),
    .A2(_06401_),
    .ZN(_06402_));
 BUF_X2 _28828_ (.A(_06402_),
    .Z(_06403_));
 BUF_X4 _28829_ (.A(_06403_),
    .Z(_06404_));
 BUF_X4 _28830_ (.A(_06404_),
    .Z(_06405_));
 NOR2_X1 _28831_ (.A1(\core.dec_block.block_w3_reg[0] ),
    .A2(_06405_),
    .ZN(_06406_));
 BUF_X4 _28832_ (.A(_06403_),
    .Z(_06407_));
 XNOR2_X1 _28833_ (.A(\block_reg[0][0] ),
    .B(_16550_),
    .ZN(_06408_));
 OAI221_X1 _28834_ (.A(_06407_),
    .B1(_06408_),
    .B2(_06225_),
    .C1(_19027_),
    .C2(_06199_),
    .ZN(_06409_));
 XOR2_X1 _28835_ (.A(_04589_),
    .B(_05879_),
    .Z(_06410_));
 XNOR2_X1 _28836_ (.A(_05188_),
    .B(_06410_),
    .ZN(_06411_));
 XNOR2_X2 _28837_ (.A(_04816_),
    .B(_06411_),
    .ZN(_06412_));
 AOI21_X1 _28838_ (.A(_06409_),
    .B1(_06412_),
    .B2(_06212_),
    .ZN(_06413_));
 AOI21_X1 _28839_ (.A(_06406_),
    .B1(_06413_),
    .B2(_16851_),
    .ZN(_00663_));
 XNOR2_X1 _28840_ (.A(\block_reg[1][10] ),
    .B(_05157_),
    .ZN(_06414_));
 OAI22_X1 _28841_ (.A1(_16555_),
    .A2(_19412_),
    .B1(_06414_),
    .B2(_18552_),
    .ZN(_06415_));
 NOR2_X1 _28842_ (.A1(_17503_),
    .A2(_06415_),
    .ZN(_06416_));
 XNOR2_X1 _28843_ (.A(_03575_),
    .B(_05178_),
    .ZN(_06417_));
 XNOR2_X1 _28844_ (.A(_16875_),
    .B(_06417_),
    .ZN(_06418_));
 XNOR2_X1 _28845_ (.A(_06245_),
    .B(_06418_),
    .ZN(_06419_));
 XNOR2_X1 _28846_ (.A(_05980_),
    .B(_06419_),
    .ZN(_06420_));
 OAI21_X1 _28847_ (.A(_06416_),
    .B1(_06420_),
    .B2(_17204_),
    .ZN(_06421_));
 CLKBUF_X3 _28848_ (.A(_06404_),
    .Z(_06422_));
 MUX2_X1 _28849_ (.A(\core.dec_block.block_w3_reg[10] ),
    .B(_06421_),
    .S(_06422_),
    .Z(_00664_));
 XNOR2_X1 _28850_ (.A(_05362_),
    .B(_05392_),
    .ZN(_06423_));
 XNOR2_X1 _28851_ (.A(_06218_),
    .B(_06423_),
    .ZN(_06424_));
 XNOR2_X1 _28852_ (.A(_05999_),
    .B(_06424_),
    .ZN(_06425_));
 NOR2_X1 _28853_ (.A1(_17504_),
    .A2(_06425_),
    .ZN(_06426_));
 XNOR2_X1 _28854_ (.A(\block_reg[1][11] ),
    .B(_05384_),
    .ZN(_06427_));
 OAI221_X1 _28855_ (.A(_06404_),
    .B1(_06427_),
    .B2(_05774_),
    .C1(_03344_),
    .C2(_19180_),
    .ZN(_06428_));
 OAI33_X1 _28856_ (.A1(_17216_),
    .A2(_16353_),
    .A3(_06401_),
    .B1(_06426_),
    .B2(_06428_),
    .B3(_18051_),
    .ZN(_06429_));
 INV_X1 _28857_ (.A(_06429_),
    .ZN(_00665_));
 NOR2_X1 _28858_ (.A1(\core.dec_block.block_w3_reg[12] ),
    .A2(_06405_),
    .ZN(_06430_));
 XNOR2_X1 _28859_ (.A(_05540_),
    .B(_05608_),
    .ZN(_06431_));
 XNOR2_X1 _28860_ (.A(_05386_),
    .B(_05510_),
    .ZN(_06432_));
 XNOR2_X1 _28861_ (.A(_06431_),
    .B(_06432_),
    .ZN(_06433_));
 XNOR2_X1 _28862_ (.A(_06009_),
    .B(_06433_),
    .ZN(_06434_));
 NAND2_X1 _28863_ (.A1(_18333_),
    .A2(_06434_),
    .ZN(_06435_));
 CLKBUF_X3 _28864_ (.A(_06403_),
    .Z(_06436_));
 INV_X1 _28865_ (.A(\block_reg[1][12] ),
    .ZN(_06437_));
 XNOR2_X2 _28866_ (.A(_06437_),
    .B(_05536_),
    .ZN(_06438_));
 OAI221_X2 _28867_ (.A(_06436_),
    .B1(_06438_),
    .B2(_18553_),
    .C1(_03775_),
    .C2(_03858_),
    .ZN(_06439_));
 NOR2_X1 _28868_ (.A1(_18228_),
    .A2(_06439_),
    .ZN(_06440_));
 AOI21_X1 _28869_ (.A(_06430_),
    .B1(_06435_),
    .B2(_06440_),
    .ZN(_00666_));
 XOR2_X2 _28870_ (.A(_03523_),
    .B(_05393_),
    .Z(_06441_));
 XNOR2_X1 _28871_ (.A(_06038_),
    .B(_06441_),
    .ZN(_06442_));
 XNOR2_X1 _28872_ (.A(_05595_),
    .B(_06442_),
    .ZN(_06443_));
 NOR2_X1 _28873_ (.A1(_17504_),
    .A2(_06443_),
    .ZN(_06444_));
 XNOR2_X2 _28874_ (.A(\block_reg[1][13] ),
    .B(_17061_),
    .ZN(_06445_));
 OAI221_X2 _28875_ (.A(_06403_),
    .B1(_06445_),
    .B2(_18552_),
    .C1(_18970_),
    .C2(_19180_),
    .ZN(_06446_));
 OAI33_X1 _28876_ (.A1(\core.dec_block.block_w3_reg[13] ),
    .A2(_16353_),
    .A3(_06401_),
    .B1(_06444_),
    .B2(_06446_),
    .B3(_18398_),
    .ZN(_06447_));
 INV_X1 _28877_ (.A(_06447_),
    .ZN(_00667_));
 NOR2_X1 _28878_ (.A1(_17248_),
    .A2(_06405_),
    .ZN(_06448_));
 XNOR2_X2 _28879_ (.A(\block_reg[1][14] ),
    .B(_03595_),
    .ZN(_06449_));
 CLKBUF_X3 _28880_ (.A(_16554_),
    .Z(_06450_));
 OAI221_X2 _28881_ (.A(_06407_),
    .B1(_06449_),
    .B2(_06225_),
    .C1(_19224_),
    .C2(_06450_),
    .ZN(_06451_));
 XOR2_X1 _28882_ (.A(_03541_),
    .B(_05406_),
    .Z(_06452_));
 XNOR2_X1 _28883_ (.A(_16875_),
    .B(_05539_),
    .ZN(_06453_));
 XNOR2_X1 _28884_ (.A(_06452_),
    .B(_06453_),
    .ZN(_06454_));
 XNOR2_X1 _28885_ (.A(_06037_),
    .B(_06454_),
    .ZN(_06455_));
 XNOR2_X1 _28886_ (.A(_06052_),
    .B(_06455_),
    .ZN(_06456_));
 XNOR2_X1 _28887_ (.A(_05512_),
    .B(_06456_),
    .ZN(_06457_));
 AOI21_X1 _28888_ (.A(_06451_),
    .B1(_06457_),
    .B2(_06212_),
    .ZN(_06458_));
 AOI21_X1 _28889_ (.A(_06448_),
    .B1(_06458_),
    .B2(_18465_),
    .ZN(_00668_));
 NOR2_X1 _28890_ (.A1(\core.dec_block.block_w3_reg[15] ),
    .A2(_06405_),
    .ZN(_06459_));
 XNOR2_X2 _28891_ (.A(\block_reg[1][15] ),
    .B(_05114_),
    .ZN(_06460_));
 OAI221_X2 _28892_ (.A(_06407_),
    .B1(_06460_),
    .B2(_06225_),
    .C1(_18942_),
    .C2(_06450_),
    .ZN(_06461_));
 XNOR2_X1 _28893_ (.A(_05591_),
    .B(_06267_),
    .ZN(_06462_));
 XOR2_X1 _28894_ (.A(_03596_),
    .B(_03627_),
    .Z(_06463_));
 XNOR2_X1 _28895_ (.A(_17185_),
    .B(_06463_),
    .ZN(_06464_));
 XNOR2_X1 _28896_ (.A(_06462_),
    .B(_06464_),
    .ZN(_06465_));
 XNOR2_X1 _28897_ (.A(_06246_),
    .B(_06465_),
    .ZN(_06466_));
 CLKBUF_X3 _28898_ (.A(_17748_),
    .Z(_06467_));
 AOI21_X1 _28899_ (.A(_06461_),
    .B1(_06466_),
    .B2(_06467_),
    .ZN(_06468_));
 AOI21_X1 _28900_ (.A(_06459_),
    .B1(_06468_),
    .B2(_18526_),
    .ZN(_00669_));
 NOR2_X1 _28901_ (.A1(\core.dec_block.block_w3_reg[16] ),
    .A2(_06405_),
    .ZN(_06469_));
 XOR2_X2 _28902_ (.A(\block_reg[2][16] ),
    .B(_17905_),
    .Z(_06470_));
 CLKBUF_X3 _28903_ (.A(_17709_),
    .Z(_06471_));
 OAI221_X1 _28904_ (.A(_06407_),
    .B1(_06470_),
    .B2(_06471_),
    .C1(_19226_),
    .C2(_06450_),
    .ZN(_06472_));
 XOR2_X1 _28905_ (.A(_17658_),
    .B(_06074_),
    .Z(_06473_));
 XNOR2_X1 _28906_ (.A(_05905_),
    .B(_06473_),
    .ZN(_06474_));
 XNOR2_X1 _28907_ (.A(_17850_),
    .B(_06282_),
    .ZN(_06475_));
 XNOR2_X2 _28908_ (.A(_06474_),
    .B(_06475_),
    .ZN(_06476_));
 AOI21_X1 _28909_ (.A(_06472_),
    .B1(_06476_),
    .B2(_06467_),
    .ZN(_06477_));
 AOI21_X1 _28910_ (.A(_06469_),
    .B1(_06477_),
    .B2(_18848_),
    .ZN(_00670_));
 NOR2_X1 _28911_ (.A1(\core.dec_block.block_w3_reg[17] ),
    .A2(_06405_),
    .ZN(_06478_));
 XNOR2_X2 _28912_ (.A(_17848_),
    .B(_17762_),
    .ZN(_06479_));
 XOR2_X1 _28913_ (.A(_17672_),
    .B(_05776_),
    .Z(_06480_));
 XNOR2_X1 _28914_ (.A(_06479_),
    .B(_06480_),
    .ZN(_06481_));
 XNOR2_X2 _28915_ (.A(_05904_),
    .B(_06481_),
    .ZN(_06482_));
 NOR2_X1 _28916_ (.A1(_17204_),
    .A2(_06482_),
    .ZN(_06483_));
 XNOR2_X2 _28917_ (.A(\block_reg[2][17] ),
    .B(_18258_),
    .ZN(_06484_));
 OAI221_X1 _28918_ (.A(_06436_),
    .B1(_06484_),
    .B2(_18553_),
    .C1(_19445_),
    .C2(_05021_),
    .ZN(_06485_));
 NOR2_X1 _28919_ (.A1(_06483_),
    .A2(_06485_),
    .ZN(_06486_));
 AOI21_X1 _28920_ (.A(_06478_),
    .B1(_06486_),
    .B2(_19179_),
    .ZN(_00671_));
 NOR2_X1 _28921_ (.A1(\core.dec_block.block_w3_reg[18] ),
    .A2(_06405_),
    .ZN(_06487_));
 XNOR2_X2 _28922_ (.A(\block_reg[2][18] ),
    .B(_17562_),
    .ZN(_06488_));
 OAI221_X1 _28923_ (.A(_06407_),
    .B1(_06488_),
    .B2(_06471_),
    .C1(_03332_),
    .C2(_06450_),
    .ZN(_06489_));
 XOR2_X1 _28924_ (.A(_17535_),
    .B(_17658_),
    .Z(_06490_));
 XNOR2_X1 _28925_ (.A(_18260_),
    .B(_06490_),
    .ZN(_06491_));
 XNOR2_X1 _28926_ (.A(_17703_),
    .B(_06491_),
    .ZN(_06492_));
 XNOR2_X2 _28927_ (.A(_06029_),
    .B(_06492_),
    .ZN(_06493_));
 AOI21_X1 _28928_ (.A(_06489_),
    .B1(_06493_),
    .B2(_06467_),
    .ZN(_06494_));
 AOI21_X1 _28929_ (.A(_06487_),
    .B1(_06494_),
    .B2(_19371_),
    .ZN(_00672_));
 NOR2_X1 _28930_ (.A1(\core.dec_block.block_w3_reg[19] ),
    .A2(_06405_),
    .ZN(_06495_));
 XOR2_X2 _28931_ (.A(\block_reg[2][19] ),
    .B(_17810_),
    .Z(_06496_));
 OAI221_X1 _28932_ (.A(_06407_),
    .B1(_06496_),
    .B2(_06471_),
    .C1(_03762_),
    .C2(_06450_),
    .ZN(_06497_));
 XOR2_X1 _28933_ (.A(_17552_),
    .B(_17866_),
    .Z(_06498_));
 XNOR2_X1 _28934_ (.A(_06303_),
    .B(_06498_),
    .ZN(_06499_));
 XNOR2_X2 _28935_ (.A(_06063_),
    .B(_06499_),
    .ZN(_06500_));
 AOI21_X1 _28936_ (.A(_06497_),
    .B1(_06500_),
    .B2(_06467_),
    .ZN(_06501_));
 AOI21_X1 _28937_ (.A(_06495_),
    .B1(_06501_),
    .B2(_19519_),
    .ZN(_00673_));
 BUF_X4 _28938_ (.A(_06404_),
    .Z(_06502_));
 NOR2_X1 _28939_ (.A1(\core.dec_block.block_w3_reg[1] ),
    .A2(_06502_),
    .ZN(_06503_));
 INV_X1 _28940_ (.A(\block_reg[0][1] ),
    .ZN(_06504_));
 XNOR2_X2 _28941_ (.A(_06504_),
    .B(_03509_),
    .ZN(_06505_));
 OAI221_X1 _28942_ (.A(_03498_),
    .B1(_06505_),
    .B2(_06471_),
    .C1(_19285_),
    .C2(_06450_),
    .ZN(_06506_));
 XOR2_X1 _28943_ (.A(_03976_),
    .B(_05015_),
    .Z(_06507_));
 XNOR2_X1 _28944_ (.A(_05859_),
    .B(_06394_),
    .ZN(_06508_));
 XNOR2_X1 _28945_ (.A(_06507_),
    .B(_06508_),
    .ZN(_06509_));
 XNOR2_X1 _28946_ (.A(_05882_),
    .B(_05925_),
    .ZN(_06510_));
 XNOR2_X2 _28947_ (.A(_06509_),
    .B(_06510_),
    .ZN(_06511_));
 AOI21_X1 _28948_ (.A(_06506_),
    .B1(_06511_),
    .B2(_06467_),
    .ZN(_06512_));
 AOI21_X1 _28949_ (.A(_06503_),
    .B1(_06512_),
    .B2(_06405_),
    .ZN(_00674_));
 NOR2_X1 _28950_ (.A1(\core.dec_block.block_w3_reg[20] ),
    .A2(_06502_),
    .ZN(_06513_));
 XOR2_X2 _28951_ (.A(\block_reg[2][20] ),
    .B(_18296_),
    .Z(_06514_));
 OAI221_X1 _28952_ (.A(_06407_),
    .B1(_06514_),
    .B2(_06471_),
    .C1(_03790_),
    .C2(_06450_),
    .ZN(_06515_));
 XOR2_X1 _28953_ (.A(_18310_),
    .B(_18337_),
    .Z(_06516_));
 XNOR2_X1 _28954_ (.A(_18482_),
    .B(_06516_),
    .ZN(_06517_));
 XNOR2_X1 _28955_ (.A(_18282_),
    .B(_06517_),
    .ZN(_06518_));
 XNOR2_X1 _28956_ (.A(_18269_),
    .B(_06518_),
    .ZN(_06519_));
 XNOR2_X2 _28957_ (.A(_06078_),
    .B(_06519_),
    .ZN(_06520_));
 AOI21_X1 _28958_ (.A(_06515_),
    .B1(_06520_),
    .B2(_06467_),
    .ZN(_06521_));
 AOI21_X1 _28959_ (.A(_06513_),
    .B1(_06521_),
    .B2(_03698_),
    .ZN(_00675_));
 NOR2_X1 _28960_ (.A1(\core.dec_block.block_w3_reg[21] ),
    .A2(_06502_),
    .ZN(_06522_));
 XOR2_X1 _28961_ (.A(_18283_),
    .B(_18487_),
    .Z(_06523_));
 XNOR2_X1 _28962_ (.A(_06099_),
    .B(_06523_),
    .ZN(_06524_));
 XNOR2_X1 _28963_ (.A(_18336_),
    .B(_06524_),
    .ZN(_06525_));
 NAND2_X2 _28964_ (.A1(_18333_),
    .A2(_06525_),
    .ZN(_06526_));
 XNOR2_X2 _28965_ (.A(\block_reg[2][21] ),
    .B(_17890_),
    .ZN(_06527_));
 OAI221_X1 _28966_ (.A(_06436_),
    .B1(_06527_),
    .B2(_18553_),
    .C1(_18909_),
    .C2(_03858_),
    .ZN(_06528_));
 NOR2_X1 _28967_ (.A1(_03845_),
    .A2(_06528_),
    .ZN(_06529_));
 AOI21_X1 _28968_ (.A(_06522_),
    .B1(_06526_),
    .B2(_06529_),
    .ZN(_00676_));
 NOR2_X1 _28969_ (.A1(\core.dec_block.block_w3_reg[22] ),
    .A2(_06502_),
    .ZN(_06530_));
 XNOR2_X1 _28970_ (.A(\block_reg[2][22] ),
    .B(_17573_),
    .ZN(_06531_));
 OAI221_X1 _28971_ (.A(_06407_),
    .B1(_06531_),
    .B2(_06471_),
    .C1(_18921_),
    .C2(_06450_),
    .ZN(_06532_));
 XOR2_X2 _28972_ (.A(_18282_),
    .B(_18297_),
    .Z(_06533_));
 XNOR2_X2 _28973_ (.A(_05719_),
    .B(_06533_),
    .ZN(_06534_));
 XNOR2_X2 _28974_ (.A(_18486_),
    .B(_06534_),
    .ZN(_06535_));
 AOI21_X1 _28975_ (.A(_06532_),
    .B1(_06535_),
    .B2(_06467_),
    .ZN(_06536_));
 AOI21_X1 _28976_ (.A(_06530_),
    .B1(_06536_),
    .B2(_03893_),
    .ZN(_00677_));
 NOR2_X1 _28977_ (.A1(_18576_),
    .A2(_06502_),
    .ZN(_06537_));
 XOR2_X1 _28978_ (.A(_18311_),
    .B(_06031_),
    .Z(_06538_));
 XNOR2_X1 _28979_ (.A(_06479_),
    .B(_06538_),
    .ZN(_06539_));
 XNOR2_X1 _28980_ (.A(_18340_),
    .B(_06539_),
    .ZN(_06540_));
 NAND2_X1 _28981_ (.A1(_18333_),
    .A2(_06540_),
    .ZN(_06541_));
 INV_X1 _28982_ (.A(\block_reg[2][23] ),
    .ZN(_06542_));
 XNOR2_X1 _28983_ (.A(_06542_),
    .B(_17551_),
    .ZN(_06543_));
 OAI221_X1 _28984_ (.A(_06436_),
    .B1(_06543_),
    .B2(_18412_),
    .C1(_18956_),
    .C2(_03858_),
    .ZN(_06544_));
 NOR2_X1 _28985_ (.A1(_03955_),
    .A2(_06544_),
    .ZN(_06545_));
 AOI21_X1 _28986_ (.A(_06537_),
    .B1(_06541_),
    .B2(_06545_),
    .ZN(_00678_));
 INV_X1 _28987_ (.A(\block_reg[3][24] ),
    .ZN(_06546_));
 XNOR2_X1 _28988_ (.A(_06546_),
    .B(_18981_),
    .ZN(_06547_));
 OAI221_X1 _28989_ (.A(_06436_),
    .B1(_06547_),
    .B2(_04266_),
    .C1(_18982_),
    .C2(_05021_),
    .ZN(_06548_));
 XOR2_X1 _28990_ (.A(_19248_),
    .B(_06228_),
    .Z(_06549_));
 OAI21_X1 _28991_ (.A(_04251_),
    .B1(_06549_),
    .B2(_17504_),
    .ZN(_06550_));
 OAI22_X1 _28992_ (.A1(\core.dec_block.block_w3_reg[24] ),
    .A2(_06405_),
    .B1(_06548_),
    .B2(_06550_),
    .ZN(_06551_));
 INV_X1 _28993_ (.A(_06551_),
    .ZN(_00679_));
 NOR2_X1 _28994_ (.A1(\core.dec_block.block_w3_reg[25] ),
    .A2(_06502_),
    .ZN(_06552_));
 XNOR2_X1 _28995_ (.A(\block_reg[3][25] ),
    .B(_19298_),
    .ZN(_06553_));
 OAI221_X1 _28996_ (.A(_06407_),
    .B1(_06553_),
    .B2(_06471_),
    .C1(_19299_),
    .C2(_06450_),
    .ZN(_06554_));
 XOR2_X1 _28997_ (.A(_19285_),
    .B(_19446_),
    .Z(_06555_));
 XNOR2_X1 _28998_ (.A(_18958_),
    .B(_06555_),
    .ZN(_06556_));
 XNOR2_X1 _28999_ (.A(_03301_),
    .B(_06556_),
    .ZN(_06557_));
 AOI21_X1 _29000_ (.A(_06554_),
    .B1(_06557_),
    .B2(_06467_),
    .ZN(_06558_));
 AOI21_X1 _29001_ (.A(_06552_),
    .B1(_06558_),
    .B2(_04538_),
    .ZN(_00680_));
 NOR2_X1 _29002_ (.A1(\core.dec_block.block_w3_reg[26] ),
    .A2(_06502_),
    .ZN(_06559_));
 XNOR2_X1 _29003_ (.A(_19246_),
    .B(_05840_),
    .ZN(_06560_));
 XNOR2_X1 _29004_ (.A(_19412_),
    .B(_19445_),
    .ZN(_06561_));
 XNOR2_X1 _29005_ (.A(_19299_),
    .B(_03332_),
    .ZN(_06562_));
 XNOR2_X1 _29006_ (.A(_06561_),
    .B(_06562_),
    .ZN(_06563_));
 XNOR2_X1 _29007_ (.A(_06560_),
    .B(_06563_),
    .ZN(_06564_));
 XNOR2_X1 _29008_ (.A(_05789_),
    .B(_06564_),
    .ZN(_06565_));
 NAND2_X1 _29009_ (.A1(_18333_),
    .A2(_06565_),
    .ZN(_06566_));
 XNOR2_X1 _29010_ (.A(\block_reg[3][26] ),
    .B(_19428_),
    .ZN(_06567_));
 OAI221_X1 _29011_ (.A(_06436_),
    .B1(_06567_),
    .B2(_18412_),
    .C1(_19429_),
    .C2(_03858_),
    .ZN(_06568_));
 NOR2_X1 _29012_ (.A1(_04657_),
    .A2(_06568_),
    .ZN(_06569_));
 AOI21_X1 _29013_ (.A(_06559_),
    .B1(_06566_),
    .B2(_06569_),
    .ZN(_00681_));
 XNOR2_X1 _29014_ (.A(\block_reg[3][27] ),
    .B(_03325_),
    .ZN(_06570_));
 OAI22_X1 _29015_ (.A1(_16555_),
    .A2(_03326_),
    .B1(_06570_),
    .B2(_18552_),
    .ZN(_06571_));
 NOR2_X1 _29016_ (.A1(_04792_),
    .A2(_06571_),
    .ZN(_06572_));
 XOR2_X1 _29017_ (.A(_03345_),
    .B(_03784_),
    .Z(_06573_));
 XNOR2_X1 _29018_ (.A(_05802_),
    .B(_06573_),
    .ZN(_06574_));
 OAI21_X1 _29019_ (.A(_06572_),
    .B1(_06574_),
    .B2(_17204_),
    .ZN(_06575_));
 MUX2_X1 _29020_ (.A(\core.dec_block.block_w3_reg[27] ),
    .B(_06575_),
    .S(_06422_),
    .Z(_00682_));
 NOR2_X1 _29021_ (.A1(\core.dec_block.block_w3_reg[28] ),
    .A2(_06502_),
    .ZN(_06576_));
 XNOR2_X1 _29022_ (.A(\block_reg[3][28] ),
    .B(_03738_),
    .ZN(_06577_));
 OAI221_X1 _29023_ (.A(_06407_),
    .B1(_06577_),
    .B2(_06471_),
    .C1(_03739_),
    .C2(_06450_),
    .ZN(_06578_));
 XOR2_X1 _29024_ (.A(_05797_),
    .B(_06352_),
    .Z(_06579_));
 XNOR2_X1 _29025_ (.A(_19442_),
    .B(_03959_),
    .ZN(_06580_));
 XNOR2_X1 _29026_ (.A(_06579_),
    .B(_06580_),
    .ZN(_06581_));
 XNOR2_X1 _29027_ (.A(_03727_),
    .B(_03789_),
    .ZN(_06582_));
 XNOR2_X1 _29028_ (.A(_06581_),
    .B(_06582_),
    .ZN(_06583_));
 AOI21_X1 _29029_ (.A(_06578_),
    .B1(_06583_),
    .B2(_06467_),
    .ZN(_06584_));
 AOI21_X1 _29030_ (.A(_06576_),
    .B1(_06584_),
    .B2(_04902_),
    .ZN(_00683_));
 NOR2_X1 _29031_ (.A1(\core.dec_block.block_w3_reg[29] ),
    .A2(_06502_),
    .ZN(_06585_));
 XOR2_X1 _29032_ (.A(_03739_),
    .B(_05828_),
    .Z(_06586_));
 XNOR2_X1 _29033_ (.A(_05826_),
    .B(_06586_),
    .ZN(_06587_));
 XNOR2_X1 _29034_ (.A(_03793_),
    .B(_06587_),
    .ZN(_06588_));
 NAND2_X1 _29035_ (.A1(_18333_),
    .A2(_06588_),
    .ZN(_06589_));
 XOR2_X1 _29036_ (.A(\block_reg[3][29] ),
    .B(_19001_),
    .Z(_06590_));
 OAI221_X1 _29037_ (.A(_06436_),
    .B1(_06590_),
    .B2(_18412_),
    .C1(_19002_),
    .C2(_03858_),
    .ZN(_06591_));
 NOR2_X1 _29038_ (.A1(_05003_),
    .A2(_06591_),
    .ZN(_06592_));
 AOI21_X1 _29039_ (.A(_06585_),
    .B1(_06589_),
    .B2(_06592_),
    .ZN(_00684_));
 NOR2_X1 _29040_ (.A1(\core.dec_block.block_w3_reg[2] ),
    .A2(_06502_),
    .ZN(_06593_));
 XNOR2_X1 _29041_ (.A(_19385_),
    .B(_03510_),
    .ZN(_06594_));
 XNOR2_X1 _29042_ (.A(_04552_),
    .B(_06594_),
    .ZN(_06595_));
 XNOR2_X1 _29043_ (.A(_05942_),
    .B(_06595_),
    .ZN(_06596_));
 XNOR2_X1 _29044_ (.A(_05881_),
    .B(_06596_),
    .ZN(_06597_));
 NAND2_X1 _29045_ (.A1(_04370_),
    .A2(_06597_),
    .ZN(_06598_));
 XNOR2_X2 _29046_ (.A(\block_reg[0][2] ),
    .B(_04698_),
    .ZN(_06599_));
 OAI221_X1 _29047_ (.A(_06436_),
    .B1(_06599_),
    .B2(_18412_),
    .C1(_19458_),
    .C2(_03858_),
    .ZN(_06600_));
 NOR2_X1 _29048_ (.A1(_05101_),
    .A2(_06600_),
    .ZN(_06601_));
 AOI21_X1 _29049_ (.A(_06593_),
    .B1(_06598_),
    .B2(_06601_),
    .ZN(_00685_));
 NOR2_X1 _29050_ (.A1(\core.dec_block.block_w3_reg[30] ),
    .A2(_06422_),
    .ZN(_06602_));
 XNOR2_X1 _29051_ (.A(_18884_),
    .B(_03763_),
    .ZN(_06603_));
 XNOR2_X1 _29052_ (.A(_03962_),
    .B(_06603_),
    .ZN(_06604_));
 XNOR2_X1 _29053_ (.A(_03918_),
    .B(_06604_),
    .ZN(_06605_));
 XNOR2_X1 _29054_ (.A(_05830_),
    .B(_06605_),
    .ZN(_06606_));
 NAND2_X1 _29055_ (.A1(_04370_),
    .A2(_06606_),
    .ZN(_06607_));
 XNOR2_X1 _29056_ (.A(\block_reg[3][30] ),
    .B(_19245_),
    .ZN(_06608_));
 OAI221_X1 _29057_ (.A(_06436_),
    .B1(_06608_),
    .B2(_18412_),
    .C1(_19246_),
    .C2(_18399_),
    .ZN(_06609_));
 NOR2_X1 _29058_ (.A1(_05227_),
    .A2(_06609_),
    .ZN(_06610_));
 AOI21_X1 _29059_ (.A(_06602_),
    .B1(_06607_),
    .B2(_06610_),
    .ZN(_00686_));
 NOR2_X1 _29060_ (.A1(\core.dec_block.block_w3_reg[31] ),
    .A2(_06422_),
    .ZN(_06611_));
 XNOR2_X1 _29061_ (.A(\block_reg[3][31] ),
    .B(_19440_),
    .ZN(_06612_));
 OAI221_X1 _29062_ (.A(_06404_),
    .B1(_06612_),
    .B2(_06471_),
    .C1(_19441_),
    .C2(_18479_),
    .ZN(_06613_));
 XNOR2_X1 _29063_ (.A(_19247_),
    .B(_03921_),
    .ZN(_06614_));
 XOR2_X1 _29064_ (.A(_18921_),
    .B(_03739_),
    .Z(_06615_));
 XNOR2_X1 _29065_ (.A(_18957_),
    .B(_06615_),
    .ZN(_06616_));
 XNOR2_X1 _29066_ (.A(_06614_),
    .B(_06616_),
    .ZN(_06617_));
 XNOR2_X1 _29067_ (.A(_05852_),
    .B(_06617_),
    .ZN(_06618_));
 AOI21_X1 _29068_ (.A(_06613_),
    .B1(_06618_),
    .B2(_06467_),
    .ZN(_06619_));
 AOI21_X1 _29069_ (.A(_06611_),
    .B1(_06619_),
    .B2(_05259_),
    .ZN(_00687_));
 NOR2_X1 _29070_ (.A1(\core.dec_block.block_w3_reg[3] ),
    .A2(_06422_),
    .ZN(_06620_));
 XNOR2_X1 _29071_ (.A(\block_reg[0][3] ),
    .B(_04832_),
    .ZN(_06621_));
 OAI221_X1 _29072_ (.A(_06404_),
    .B1(_06621_),
    .B2(_06471_),
    .C1(_03358_),
    .C2(_18479_),
    .ZN(_06622_));
 XNOR2_X1 _29073_ (.A(_04807_),
    .B(_05009_),
    .ZN(_06623_));
 XNOR2_X2 _29074_ (.A(_05894_),
    .B(_06623_),
    .ZN(_06624_));
 AOI21_X1 _29075_ (.A(_06622_),
    .B1(_06624_),
    .B2(_17749_),
    .ZN(_06625_));
 AOI21_X1 _29076_ (.A(_06620_),
    .B1(_06625_),
    .B2(_05344_),
    .ZN(_00688_));
 NOR2_X1 _29077_ (.A1(\core.dec_block.block_w3_reg[4] ),
    .A2(_06422_),
    .ZN(_06626_));
 XNOR2_X1 _29078_ (.A(_04723_),
    .B(_05184_),
    .ZN(_06627_));
 XNOR2_X1 _29079_ (.A(_05950_),
    .B(_06627_),
    .ZN(_06628_));
 XNOR2_X1 _29080_ (.A(_04921_),
    .B(_06628_),
    .ZN(_06629_));
 XNOR2_X2 _29081_ (.A(_05915_),
    .B(_06629_),
    .ZN(_06630_));
 NAND2_X1 _29082_ (.A1(_04370_),
    .A2(_06630_),
    .ZN(_06631_));
 INV_X1 _29083_ (.A(\block_reg[0][4] ),
    .ZN(_06632_));
 XNOR2_X1 _29084_ (.A(_06632_),
    .B(_04936_),
    .ZN(_06633_));
 OAI221_X1 _29085_ (.A(_06436_),
    .B1(_06633_),
    .B2(_18412_),
    .C1(_03760_),
    .C2(_18399_),
    .ZN(_06634_));
 NOR2_X1 _29086_ (.A1(_05477_),
    .A2(_06634_),
    .ZN(_06635_));
 AOI21_X1 _29087_ (.A(_06626_),
    .B1(_06631_),
    .B2(_06635_),
    .ZN(_00689_));
 NOR2_X1 _29088_ (.A1(\core.dec_block.block_w3_reg[5] ),
    .A2(_06422_),
    .ZN(_06636_));
 XNOR2_X1 _29089_ (.A(\block_reg[0][5] ),
    .B(_04364_),
    .ZN(_06637_));
 OAI221_X1 _29090_ (.A(_06404_),
    .B1(_06637_),
    .B2(_17710_),
    .C1(_18896_),
    .C2(_18479_),
    .ZN(_06638_));
 XOR2_X1 _29091_ (.A(_03857_),
    .B(_04937_),
    .Z(_06639_));
 XNOR2_X1 _29092_ (.A(_05942_),
    .B(_06639_),
    .ZN(_06640_));
 XNOR2_X1 _29093_ (.A(_04313_),
    .B(_06640_),
    .ZN(_06641_));
 XNOR2_X1 _29094_ (.A(_05183_),
    .B(_06641_),
    .ZN(_06642_));
 XOR2_X2 _29095_ (.A(_04700_),
    .B(_05931_),
    .Z(_06643_));
 XNOR2_X2 _29096_ (.A(_06642_),
    .B(_06643_),
    .ZN(_06644_));
 AOI21_X1 _29097_ (.A(_06638_),
    .B1(_06644_),
    .B2(_17749_),
    .ZN(_06645_));
 AOI21_X1 _29098_ (.A(_06636_),
    .B1(_06645_),
    .B2(_05589_),
    .ZN(_00690_));
 NOR2_X1 _29099_ (.A1(\core.dec_block.block_w3_reg[6] ),
    .A2(_06422_),
    .ZN(_06646_));
 XNOR2_X1 _29100_ (.A(\block_reg[0][6] ),
    .B(_04588_),
    .ZN(_06647_));
 OAI221_X1 _29101_ (.A(_06404_),
    .B1(_06647_),
    .B2(_17710_),
    .C1(_18884_),
    .C2(_18479_),
    .ZN(_06648_));
 XOR2_X2 _29102_ (.A(_05190_),
    .B(_05925_),
    .Z(_06649_));
 XNOR2_X2 _29103_ (.A(_05941_),
    .B(_06649_),
    .ZN(_06650_));
 AOI21_X1 _29104_ (.A(_06648_),
    .B1(_06650_),
    .B2(_17749_),
    .ZN(_06651_));
 AOI21_X1 _29105_ (.A(_06646_),
    .B1(_06651_),
    .B2(_05650_),
    .ZN(_00691_));
 NOR2_X1 _29106_ (.A1(\core.dec_block.block_w3_reg[7] ),
    .A2(_06422_),
    .ZN(_06652_));
 XNOR2_X1 _29107_ (.A(\block_reg[0][7] ),
    .B(_04722_),
    .ZN(_06653_));
 OAI221_X1 _29108_ (.A(_06404_),
    .B1(_06653_),
    .B2(_17710_),
    .C1(_19260_),
    .C2(_18479_),
    .ZN(_06654_));
 XOR2_X2 _29109_ (.A(_03976_),
    .B(_05007_),
    .Z(_06655_));
 XNOR2_X2 _29110_ (.A(_05952_),
    .B(_06655_),
    .ZN(_06656_));
 AOI21_X1 _29111_ (.A(_06654_),
    .B1(_06656_),
    .B2(_17749_),
    .ZN(_06657_));
 AOI21_X1 _29112_ (.A(_06652_),
    .B1(_06657_),
    .B2(_05674_),
    .ZN(_00692_));
 NOR2_X1 _29113_ (.A1(\core.dec_block.block_w3_reg[8] ),
    .A2(_06422_),
    .ZN(_06658_));
 OAI21_X1 _29114_ (.A(_06403_),
    .B1(_19016_),
    .B2(_16554_),
    .ZN(_06659_));
 XOR2_X1 _29115_ (.A(_05598_),
    .B(_05978_),
    .Z(_06660_));
 XNOR2_X1 _29116_ (.A(_16943_),
    .B(_05162_),
    .ZN(_06661_));
 XNOR2_X1 _29117_ (.A(_06660_),
    .B(_06661_),
    .ZN(_06662_));
 XNOR2_X2 _29118_ (.A(_05613_),
    .B(_06662_),
    .ZN(_06663_));
 XNOR2_X1 _29119_ (.A(\block_reg[1][8] ),
    .B(_17011_),
    .ZN(_06664_));
 AOI221_X2 _29120_ (.A(_06659_),
    .B1(_06663_),
    .B2(_17747_),
    .C1(_16372_),
    .C2(_06664_),
    .ZN(_06665_));
 AOI21_X1 _29121_ (.A(_06658_),
    .B1(_06665_),
    .B2(_05715_),
    .ZN(_00693_));
 XOR2_X2 _29122_ (.A(\block_reg[1][9] ),
    .B(_03574_),
    .Z(_06666_));
 OAI221_X2 _29123_ (.A(_06404_),
    .B1(_06666_),
    .B2(_17710_),
    .C1(_19274_),
    .C2(_18052_),
    .ZN(_06667_));
 XOR2_X1 _29124_ (.A(_17063_),
    .B(_03542_),
    .Z(_06668_));
 XNOR2_X1 _29125_ (.A(_05493_),
    .B(_06668_),
    .ZN(_06669_));
 XNOR2_X1 _29126_ (.A(_05350_),
    .B(_06669_),
    .ZN(_06670_));
 NOR2_X1 _29127_ (.A1(_05793_),
    .A2(_06670_),
    .ZN(_06671_));
 OAI33_X1 _29128_ (.A1(\core.dec_block.block_w3_reg[9] ),
    .A2(_16353_),
    .A3(_06401_),
    .B1(_06667_),
    .B2(_06671_),
    .B3(_05754_),
    .ZN(_06672_));
 INV_X1 _29129_ (.A(_06672_),
    .ZN(_00694_));
 NAND2_X1 _29130_ (.A1(\core.dec_block.ready ),
    .A2(_16264_),
    .ZN(_06673_));
 OAI21_X1 _29131_ (.A(_06673_),
    .B1(_16552_),
    .B2(_16259_),
    .ZN(_00695_));
 XNOR2_X1 _29132_ (.A(_16878_),
    .B(_16269_),
    .ZN(_06674_));
 AOI21_X1 _29133_ (.A(_06674_),
    .B1(_16263_),
    .B2(\core.dec_block.dec_ctrl_reg[0] ),
    .ZN(_00696_));
 MUX2_X1 _29134_ (.A(_22129_),
    .B(_16412_),
    .S(_16269_),
    .Z(_06675_));
 NAND2_X1 _29135_ (.A1(_16264_),
    .A2(_06675_),
    .ZN(_00697_));
 BUF_X4 _29136_ (.A(_16219_),
    .Z(_06676_));
 BUF_X4 _29137_ (.A(_06676_),
    .Z(_06677_));
 BUF_X8 _29138_ (.A(_06677_),
    .Z(_06678_));
 BUF_X4 _29139_ (.A(_06678_),
    .Z(_06679_));
 BUF_X8 _29140_ (.A(_06679_),
    .Z(_06680_));
 NAND3_X1 _29141_ (.A1(\core.dec_block.dec_ctrl_reg[1] ),
    .A2(_22128_),
    .A3(_16268_),
    .ZN(_06681_));
 XNOR2_X1 _29142_ (.A(_16272_),
    .B(_06681_),
    .ZN(_06682_));
 MUX2_X1 _29143_ (.A(_06680_),
    .B(_06682_),
    .S(_16264_),
    .Z(_00698_));
 NOR4_X1 _29144_ (.A1(_16272_),
    .A2(_16375_),
    .A3(_16376_),
    .A4(_16269_),
    .ZN(_06683_));
 XNOR2_X1 _29145_ (.A(_16273_),
    .B(_06683_),
    .ZN(_06684_));
 NAND2_X1 _29146_ (.A1(_16264_),
    .A2(_06684_),
    .ZN(_00699_));
 NOR3_X1 _29147_ (.A1(_16278_),
    .A2(_16260_),
    .A3(\core.dec_block.sword_ctr_reg[0] ),
    .ZN(_06685_));
 AOI21_X1 _29148_ (.A(_06685_),
    .B1(\core.dec_block.sword_ctr_reg[0] ),
    .B2(_16260_),
    .ZN(_06686_));
 NOR3_X1 _29149_ (.A1(_16258_),
    .A2(_16271_),
    .A3(_06686_),
    .ZN(_00700_));
 AND2_X1 _29150_ (.A1(_16260_),
    .A2(\core.dec_block.sword_ctr_reg[1] ),
    .ZN(_06687_));
 AOI21_X1 _29151_ (.A(_06687_),
    .B1(_22133_),
    .B2(_16261_),
    .ZN(_06688_));
 NOR3_X1 _29152_ (.A1(_16258_),
    .A2(_16271_),
    .A3(_06688_),
    .ZN(_00701_));
 INV_X1 _29153_ (.A(\core.enc_block.block_w0_reg[0] ),
    .ZN(_06689_));
 BUF_X4 _29154_ (.A(_00329_),
    .Z(_06690_));
 AOI21_X2 _29155_ (.A(_16246_),
    .B1(_06690_),
    .B2(_16239_),
    .ZN(_06691_));
 AOI21_X4 _29156_ (.A(_06691_),
    .B1(_06690_),
    .B2(_16235_),
    .ZN(_06692_));
 INV_X1 _29157_ (.A(_16243_),
    .ZN(_06693_));
 INV_X4 _29158_ (.A(_06690_),
    .ZN(_06694_));
 NOR4_X4 _29159_ (.A1(_16234_),
    .A2(_06693_),
    .A3(_16239_),
    .A4(_06694_),
    .ZN(_06695_));
 BUF_X4 _29160_ (.A(_06695_),
    .Z(_06696_));
 BUF_X4 _29161_ (.A(_06696_),
    .Z(_06697_));
 BUF_X8 _29162_ (.A(_06697_),
    .Z(_06698_));
 BUF_X4 _29163_ (.A(_22118_),
    .Z(_06699_));
 BUF_X8 _29164_ (.A(_06699_),
    .Z(_06700_));
 BUF_X4 _29165_ (.A(_06700_),
    .Z(_06701_));
 BUF_X4 _29166_ (.A(_06701_),
    .Z(_06702_));
 AOI21_X4 _29167_ (.A(_06692_),
    .B1(_06698_),
    .B2(_06702_),
    .ZN(_06703_));
 BUF_X4 _29168_ (.A(_06703_),
    .Z(_06704_));
 BUF_X4 _29169_ (.A(_06704_),
    .Z(_06705_));
 NAND4_X4 _29170_ (.A1(_16235_),
    .A2(_16243_),
    .A3(_16240_),
    .A4(_06690_),
    .ZN(_06706_));
 BUF_X8 _29171_ (.A(_06706_),
    .Z(_06707_));
 CLKBUF_X3 _29172_ (.A(_00368_),
    .Z(_06708_));
 NOR2_X2 _29173_ (.A1(_16200_),
    .A2(_16212_),
    .ZN(_06709_));
 BUF_X4 _29174_ (.A(_06709_),
    .Z(_06710_));
 BUF_X8 _29175_ (.A(_06710_),
    .Z(_06711_));
 NOR2_X4 _29176_ (.A1(_06708_),
    .A2(_06711_),
    .ZN(_06712_));
 CLKBUF_X3 _29177_ (.A(_22118_),
    .Z(_06713_));
 CLKBUF_X3 _29178_ (.A(\core.enc_block.block_w2_reg[3] ),
    .Z(_06714_));
 BUF_X2 _29179_ (.A(_22120_),
    .Z(_06715_));
 CLKBUF_X3 _29180_ (.A(_06715_),
    .Z(_06716_));
 AOI21_X1 _29181_ (.A(_06713_),
    .B1(_06714_),
    .B2(_06716_),
    .ZN(_06717_));
 BUF_X2 _29182_ (.A(_22122_),
    .Z(_06718_));
 INV_X1 _29183_ (.A(_06718_),
    .ZN(_06719_));
 BUF_X4 _29184_ (.A(_06719_),
    .Z(_06720_));
 BUF_X2 _29185_ (.A(\core.enc_block.block_w1_reg[3] ),
    .Z(_06721_));
 INV_X1 _29186_ (.A(_06721_),
    .ZN(_06722_));
 BUF_X4 _29187_ (.A(_16250_),
    .Z(_06723_));
 OAI221_X2 _29188_ (.A(_06717_),
    .B1(_06720_),
    .B2(_06722_),
    .C1(_00370_),
    .C2(_06723_),
    .ZN(_06724_));
 BUF_X4 _29189_ (.A(_06699_),
    .Z(_06725_));
 NAND2_X2 _29190_ (.A1(_06725_),
    .A2(_00369_),
    .ZN(_06726_));
 AND4_X2 _29191_ (.A1(_06696_),
    .A2(_06710_),
    .A3(_06724_),
    .A4(_06726_),
    .ZN(_06727_));
 BUF_X4 _29192_ (.A(_06727_),
    .Z(_06728_));
 NOR2_X1 _29193_ (.A1(_06712_),
    .A2(_06728_),
    .ZN(_06729_));
 BUF_X4 _29194_ (.A(_06729_),
    .Z(_06730_));
 BUF_X4 _29195_ (.A(_06730_),
    .Z(_06731_));
 BUF_X4 _29196_ (.A(_06695_),
    .Z(_06732_));
 BUF_X16 _29197_ (.A(_06732_),
    .Z(_06733_));
 BUF_X4 _29198_ (.A(_06709_),
    .Z(_06734_));
 BUF_X8 _29199_ (.A(_06734_),
    .Z(_06735_));
 NAND2_X2 _29200_ (.A1(_06701_),
    .A2(_00358_),
    .ZN(_06736_));
 BUF_X4 _29201_ (.A(\core.enc_block.block_w2_reg[7] ),
    .Z(_06737_));
 BUF_X4 _29202_ (.A(_06715_),
    .Z(_06738_));
 AOI21_X1 _29203_ (.A(_06713_),
    .B1(_06737_),
    .B2(_06738_),
    .ZN(_06739_));
 CLKBUF_X3 _29204_ (.A(\core.enc_block.block_w1_reg[7] ),
    .Z(_06740_));
 INV_X1 _29205_ (.A(_06740_),
    .ZN(_06741_));
 BUF_X2 _29206_ (.A(_00359_),
    .Z(_06742_));
 OAI221_X2 _29207_ (.A(_06739_),
    .B1(_06720_),
    .B2(_06741_),
    .C1(_06742_),
    .C2(_06723_),
    .ZN(_06743_));
 NAND4_X4 _29208_ (.A1(_06733_),
    .A2(_06735_),
    .A3(_06736_),
    .A4(_06743_),
    .ZN(_06744_));
 BUF_X8 _29209_ (.A(_06734_),
    .Z(_06745_));
 NOR2_X4 _29210_ (.A1(_00354_),
    .A2(_06745_),
    .ZN(_06746_));
 NAND2_X2 _29211_ (.A1(_06700_),
    .A2(_00355_),
    .ZN(_06747_));
 CLKBUF_X3 _29212_ (.A(\core.enc_block.block_w2_reg[6] ),
    .Z(_06748_));
 AOI21_X1 _29213_ (.A(_06699_),
    .B1(_06748_),
    .B2(_06738_),
    .ZN(_06749_));
 BUF_X4 _29214_ (.A(_06719_),
    .Z(_06750_));
 CLKBUF_X3 _29215_ (.A(\core.enc_block.block_w1_reg[6] ),
    .Z(_06751_));
 INV_X1 _29216_ (.A(_06751_),
    .ZN(_06752_));
 OAI221_X2 _29217_ (.A(_06749_),
    .B1(_06750_),
    .B2(_06752_),
    .C1(_00356_),
    .C2(_16250_),
    .ZN(_06753_));
 AND4_X1 _29218_ (.A1(_06732_),
    .A2(_06734_),
    .A3(_06747_),
    .A4(_06753_),
    .ZN(_06754_));
 BUF_X4 _29219_ (.A(_06754_),
    .Z(_06755_));
 INV_X2 _29220_ (.A(\core.keymem.prev_key1_reg[7] ),
    .ZN(_06756_));
 BUF_X8 _29221_ (.A(_06735_),
    .Z(_06757_));
 OAI221_X2 _29222_ (.A(_06744_),
    .B1(_06746_),
    .B2(_06755_),
    .C1(_06756_),
    .C2(_06757_),
    .ZN(_06758_));
 BUF_X4 _29223_ (.A(_06758_),
    .Z(_06759_));
 BUF_X4 _29224_ (.A(_06695_),
    .Z(_06760_));
 BUF_X4 _29225_ (.A(\core.enc_block.block_w2_reg[5] ),
    .Z(_06761_));
 AOI21_X1 _29226_ (.A(_06713_),
    .B1(_06761_),
    .B2(_06716_),
    .ZN(_06762_));
 CLKBUF_X3 _29227_ (.A(\core.enc_block.block_w1_reg[5] ),
    .Z(_06763_));
 INV_X1 _29228_ (.A(_06763_),
    .ZN(_06764_));
 OAI221_X2 _29229_ (.A(_06762_),
    .B1(_06720_),
    .B2(_06764_),
    .C1(_00353_),
    .C2(_06723_),
    .ZN(_06765_));
 NAND2_X2 _29230_ (.A1(_06701_),
    .A2(_00352_),
    .ZN(_06766_));
 NAND4_X4 _29231_ (.A1(_06760_),
    .A2(_06745_),
    .A3(_06765_),
    .A4(_06766_),
    .ZN(_06767_));
 BUF_X4 _29232_ (.A(\core.enc_block.block_w2_reg[4] ),
    .Z(_06768_));
 AOI21_X1 _29233_ (.A(_06699_),
    .B1(_06768_),
    .B2(_06738_),
    .ZN(_06769_));
 CLKBUF_X3 _29234_ (.A(\core.enc_block.block_w1_reg[4] ),
    .Z(_06770_));
 INV_X1 _29235_ (.A(_06770_),
    .ZN(_06771_));
 OAI221_X2 _29236_ (.A(_06769_),
    .B1(_06750_),
    .B2(_06771_),
    .C1(_00350_),
    .C2(_06723_),
    .ZN(_06772_));
 NAND2_X2 _29237_ (.A1(_06725_),
    .A2(_00349_),
    .ZN(_06773_));
 AND4_X4 _29238_ (.A1(_06732_),
    .A2(_06734_),
    .A3(_06772_),
    .A4(_06773_),
    .ZN(_06774_));
 BUF_X4 _29239_ (.A(\core.keymem.prev_key1_reg[4] ),
    .Z(_06775_));
 INV_X4 _29240_ (.A(_06775_),
    .ZN(_06776_));
 NOR2_X4 _29241_ (.A1(_06776_),
    .A2(_06710_),
    .ZN(_06777_));
 BUF_X4 _29242_ (.A(_00351_),
    .Z(_06778_));
 BUF_X8 _29243_ (.A(_06735_),
    .Z(_06779_));
 OAI221_X2 _29244_ (.A(_06767_),
    .B1(_06774_),
    .B2(_06777_),
    .C1(_06778_),
    .C2(_06779_),
    .ZN(_06780_));
 BUF_X4 _29245_ (.A(_06780_),
    .Z(_06781_));
 NOR2_X2 _29246_ (.A1(_06759_),
    .A2(_06781_),
    .ZN(_06782_));
 BUF_X4 _29247_ (.A(_00365_),
    .Z(_06783_));
 INV_X1 _29248_ (.A(_06783_),
    .ZN(_06784_));
 OR2_X1 _29249_ (.A1(_16200_),
    .A2(_16212_),
    .ZN(_06785_));
 BUF_X8 _29250_ (.A(_06785_),
    .Z(_06786_));
 NAND2_X4 _29251_ (.A1(_06784_),
    .A2(_06786_),
    .ZN(_06787_));
 CLKBUF_X3 _29252_ (.A(\core.enc_block.block_w2_reg[2] ),
    .Z(_06788_));
 AOI21_X1 _29253_ (.A(_06713_),
    .B1(_06788_),
    .B2(_06738_),
    .ZN(_06789_));
 CLKBUF_X3 _29254_ (.A(\core.enc_block.block_w1_reg[2] ),
    .Z(_06790_));
 INV_X1 _29255_ (.A(_06790_),
    .ZN(_06791_));
 OAI221_X2 _29256_ (.A(_06789_),
    .B1(_06720_),
    .B2(_06791_),
    .C1(_00367_),
    .C2(_06723_),
    .ZN(_06792_));
 NAND2_X2 _29257_ (.A1(_06725_),
    .A2(_00366_),
    .ZN(_06793_));
 NAND4_X4 _29258_ (.A1(_06733_),
    .A2(_06735_),
    .A3(_06792_),
    .A4(_06793_),
    .ZN(_06794_));
 NAND2_X4 _29259_ (.A1(_06787_),
    .A2(_06794_),
    .ZN(_06795_));
 BUF_X4 _29260_ (.A(_00362_),
    .Z(_06796_));
 INV_X1 _29261_ (.A(_06796_),
    .ZN(_06797_));
 NAND2_X2 _29262_ (.A1(_06797_),
    .A2(_06786_),
    .ZN(_06798_));
 BUF_X8 _29263_ (.A(_06798_),
    .Z(_06799_));
 CLKBUF_X3 _29264_ (.A(\core.enc_block.block_w2_reg[1] ),
    .Z(_06800_));
 AOI21_X1 _29265_ (.A(_06713_),
    .B1(_06800_),
    .B2(_06716_),
    .ZN(_06801_));
 CLKBUF_X3 _29266_ (.A(\core.enc_block.block_w1_reg[1] ),
    .Z(_06802_));
 INV_X1 _29267_ (.A(_06802_),
    .ZN(_06803_));
 OAI221_X2 _29268_ (.A(_06801_),
    .B1(_06720_),
    .B2(_06803_),
    .C1(_00364_),
    .C2(_16251_),
    .ZN(_06804_));
 NAND2_X2 _29269_ (.A1(_06701_),
    .A2(_00363_),
    .ZN(_06805_));
 NAND4_X4 _29270_ (.A1(_06733_),
    .A2(_06735_),
    .A3(_06804_),
    .A4(_06805_),
    .ZN(_06806_));
 NAND2_X4 _29271_ (.A1(_06799_),
    .A2(_06806_),
    .ZN(_06807_));
 BUF_X4 _29272_ (.A(_06807_),
    .Z(_06808_));
 NOR2_X2 _29273_ (.A1(_06795_),
    .A2(_06808_),
    .ZN(_06809_));
 BUF_X8 _29274_ (.A(_06786_),
    .Z(_06810_));
 NAND2_X4 _29275_ (.A1(_06775_),
    .A2(_06810_),
    .ZN(_06811_));
 NAND4_X4 _29276_ (.A1(_06733_),
    .A2(_06735_),
    .A3(_06772_),
    .A4(_06773_),
    .ZN(_06812_));
 INV_X1 _29277_ (.A(_06778_),
    .ZN(_06813_));
 NAND2_X4 _29278_ (.A1(_06813_),
    .A2(_06810_),
    .ZN(_06814_));
 NAND4_X4 _29279_ (.A1(_06811_),
    .A2(_06812_),
    .A3(_06814_),
    .A4(_06767_),
    .ZN(_06815_));
 AND4_X4 _29280_ (.A1(_06696_),
    .A2(_06710_),
    .A3(_06736_),
    .A4(_06743_),
    .ZN(_06816_));
 NOR2_X4 _29281_ (.A1(_00357_),
    .A2(_06745_),
    .ZN(_06817_));
 OAI22_X4 _29282_ (.A1(_06755_),
    .A2(_06746_),
    .B1(_06816_),
    .B2(_06817_),
    .ZN(_06818_));
 NOR2_X2 _29283_ (.A1(_06815_),
    .A2(_06818_),
    .ZN(_06819_));
 BUF_X8 _29284_ (.A(_06710_),
    .Z(_06820_));
 NAND4_X4 _29285_ (.A1(_06733_),
    .A2(_06820_),
    .A3(_06747_),
    .A4(_06753_),
    .ZN(_06821_));
 BUF_X4 _29286_ (.A(_06779_),
    .Z(_06822_));
 CLKBUF_X3 _29287_ (.A(\core.keymem.prev_key1_reg[6] ),
    .Z(_06823_));
 INV_X1 _29288_ (.A(_06823_),
    .ZN(_06824_));
 OAI221_X2 _29289_ (.A(_06821_),
    .B1(_06816_),
    .B2(_06817_),
    .C1(_06822_),
    .C2(_06824_),
    .ZN(_06825_));
 BUF_X4 _29290_ (.A(_06825_),
    .Z(_06826_));
 NOR2_X4 _29291_ (.A1(_06781_),
    .A2(_06826_),
    .ZN(_06827_));
 AOI221_X2 _29292_ (.A(_06782_),
    .B1(_06809_),
    .B2(_06819_),
    .C1(_06827_),
    .C2(_06795_),
    .ZN(_06828_));
 NOR2_X4 _29293_ (.A1(_06815_),
    .A2(_06759_),
    .ZN(_06829_));
 NOR2_X4 _29294_ (.A1(_06783_),
    .A2(_06820_),
    .ZN(_06830_));
 AND4_X1 _29295_ (.A1(_06732_),
    .A2(_06710_),
    .A3(_06792_),
    .A4(_06793_),
    .ZN(_06831_));
 BUF_X4 _29296_ (.A(_06831_),
    .Z(_06832_));
 NOR4_X4 _29297_ (.A1(_06712_),
    .A2(_06728_),
    .A3(_06830_),
    .A4(_06832_),
    .ZN(_06833_));
 NOR2_X4 _29298_ (.A1(_06778_),
    .A2(_06745_),
    .ZN(_06834_));
 BUF_X4 _29299_ (.A(_06734_),
    .Z(_06835_));
 AND4_X4 _29300_ (.A1(_06696_),
    .A2(_06835_),
    .A3(_06765_),
    .A4(_06766_),
    .ZN(_06836_));
 BUF_X8 _29301_ (.A(_06820_),
    .Z(_06837_));
 OAI221_X2 _29302_ (.A(_06812_),
    .B1(_06834_),
    .B2(_06836_),
    .C1(_06837_),
    .C2(_06776_),
    .ZN(_06838_));
 NOR2_X4 _29303_ (.A1(_06818_),
    .A2(_06838_),
    .ZN(_06839_));
 INV_X1 _29304_ (.A(_06708_),
    .ZN(_06840_));
 BUF_X8 _29305_ (.A(_06810_),
    .Z(_06841_));
 NAND2_X4 _29306_ (.A1(_06840_),
    .A2(_06841_),
    .ZN(_06842_));
 BUF_X8 _29307_ (.A(_06760_),
    .Z(_06843_));
 NAND4_X4 _29308_ (.A1(_06843_),
    .A2(_06779_),
    .A3(_06724_),
    .A4(_06726_),
    .ZN(_06844_));
 BUF_X8 _29309_ (.A(_06794_),
    .Z(_06845_));
 AOI22_X4 _29310_ (.A1(_06842_),
    .A2(_06844_),
    .B1(_06787_),
    .B2(_06845_),
    .ZN(_06846_));
 BUF_X4 _29311_ (.A(_06846_),
    .Z(_06847_));
 AOI22_X1 _29312_ (.A1(_06829_),
    .A2(_06833_),
    .B1(_06839_),
    .B2(_06847_),
    .ZN(_06848_));
 NOR2_X4 _29313_ (.A1(_06796_),
    .A2(_06820_),
    .ZN(_06849_));
 AND4_X1 _29314_ (.A1(_06696_),
    .A2(_06710_),
    .A3(_06804_),
    .A4(_06805_),
    .ZN(_06850_));
 BUF_X4 _29315_ (.A(_06850_),
    .Z(_06851_));
 NOR2_X4 _29316_ (.A1(_06849_),
    .A2(_06851_),
    .ZN(_06852_));
 BUF_X4 _29317_ (.A(_06852_),
    .Z(_06853_));
 OAI22_X2 _29318_ (.A1(_06731_),
    .A2(_06828_),
    .B1(_06848_),
    .B2(_06853_),
    .ZN(_06854_));
 BUF_X4 _29319_ (.A(_06815_),
    .Z(_06855_));
 BUF_X4 _29320_ (.A(_06826_),
    .Z(_06856_));
 NOR2_X4 _29321_ (.A1(_06855_),
    .A2(_06856_),
    .ZN(_06857_));
 BUF_X4 _29322_ (.A(\core.keymem.prev_key1_reg[0] ),
    .Z(_06858_));
 INV_X2 _29323_ (.A(_06858_),
    .ZN(_06859_));
 NOR2_X4 _29324_ (.A1(_06859_),
    .A2(_06779_),
    .ZN(_06860_));
 CLKBUF_X3 _29325_ (.A(\core.enc_block.block_w2_reg[0] ),
    .Z(_06861_));
 AOI21_X1 _29326_ (.A(_06700_),
    .B1(_06861_),
    .B2(_06716_),
    .ZN(_06862_));
 CLKBUF_X3 _29327_ (.A(\core.enc_block.block_w1_reg[0] ),
    .Z(_06863_));
 INV_X1 _29328_ (.A(_06863_),
    .ZN(_06864_));
 OAI221_X2 _29329_ (.A(_06862_),
    .B1(_06720_),
    .B2(_06864_),
    .C1(_00361_),
    .C2(_16251_),
    .ZN(_06865_));
 BUF_X4 _29330_ (.A(_06700_),
    .Z(_06866_));
 BUF_X2 _29331_ (.A(_00360_),
    .Z(_06867_));
 NAND2_X1 _29332_ (.A1(_06866_),
    .A2(_06867_),
    .ZN(_06868_));
 AND4_X1 _29333_ (.A1(_06760_),
    .A2(_06835_),
    .A3(_06865_),
    .A4(_06868_),
    .ZN(_06869_));
 BUF_X4 _29334_ (.A(_06869_),
    .Z(_06870_));
 NOR2_X4 _29335_ (.A1(_06860_),
    .A2(_06870_),
    .ZN(_06871_));
 BUF_X4 _29336_ (.A(_06871_),
    .Z(_06872_));
 AOI21_X1 _29337_ (.A(_06847_),
    .B1(_06833_),
    .B2(_06872_),
    .ZN(_06873_));
 BUF_X4 _29338_ (.A(_06852_),
    .Z(_06874_));
 OAI21_X1 _29339_ (.A(_06857_),
    .B1(_06873_),
    .B2(_06874_),
    .ZN(_06875_));
 BUF_X4 _29340_ (.A(_06759_),
    .Z(_06876_));
 OAI22_X4 _29341_ (.A1(_06712_),
    .A2(_06728_),
    .B1(_06849_),
    .B2(_06851_),
    .ZN(_06877_));
 NOR3_X1 _29342_ (.A1(_06855_),
    .A2(_06876_),
    .A3(_06877_),
    .ZN(_06878_));
 NOR2_X2 _29343_ (.A1(_06834_),
    .A2(_06836_),
    .ZN(_06879_));
 CLKBUF_X3 _29344_ (.A(_06879_),
    .Z(_06880_));
 NAND2_X2 _29345_ (.A1(\core.keymem.prev_key1_reg[7] ),
    .A2(_06810_),
    .ZN(_06881_));
 NAND2_X2 _29346_ (.A1(_06823_),
    .A2(_06810_),
    .ZN(_06882_));
 NAND4_X4 _29347_ (.A1(_06821_),
    .A2(_06744_),
    .A3(_06881_),
    .A4(_06882_),
    .ZN(_06883_));
 BUF_X4 _29348_ (.A(_06883_),
    .Z(_06884_));
 BUF_X4 _29349_ (.A(_06884_),
    .Z(_06885_));
 BUF_X4 _29350_ (.A(_06837_),
    .Z(_06886_));
 BUF_X4 _29351_ (.A(_06886_),
    .Z(_06887_));
 BUF_X4 _29352_ (.A(_06887_),
    .Z(_06888_));
 OAI221_X2 _29353_ (.A(_06767_),
    .B1(_06755_),
    .B2(_06746_),
    .C1(_06888_),
    .C2(_06778_),
    .ZN(_06889_));
 NOR2_X1 _29354_ (.A1(_06816_),
    .A2(_06817_),
    .ZN(_06890_));
 CLKBUF_X3 _29355_ (.A(_06890_),
    .Z(_06891_));
 OAI22_X1 _29356_ (.A1(_06880_),
    .A2(_06885_),
    .B1(_06889_),
    .B2(_06891_),
    .ZN(_06892_));
 NAND2_X4 _29357_ (.A1(_06842_),
    .A2(_06844_),
    .ZN(_06893_));
 BUF_X4 _29358_ (.A(_06893_),
    .Z(_06894_));
 NAND2_X1 _29359_ (.A1(_06811_),
    .A2(_06812_),
    .ZN(_06895_));
 NOR2_X1 _29360_ (.A1(_06894_),
    .A2(_06895_),
    .ZN(_06896_));
 AOI21_X1 _29361_ (.A(_06878_),
    .B1(_06892_),
    .B2(_06896_),
    .ZN(_06897_));
 NOR2_X4 _29362_ (.A1(_06830_),
    .A2(_06832_),
    .ZN(_06898_));
 BUF_X4 _29363_ (.A(_06898_),
    .Z(_06899_));
 BUF_X4 _29364_ (.A(_06899_),
    .Z(_06900_));
 OAI21_X1 _29365_ (.A(_06875_),
    .B1(_06897_),
    .B2(_06900_),
    .ZN(_06901_));
 BUF_X4 _29366_ (.A(_06781_),
    .Z(_06902_));
 NOR4_X1 _29367_ (.A1(_06730_),
    .A2(_06852_),
    .A3(_06902_),
    .A4(_06884_),
    .ZN(_06903_));
 BUF_X4 _29368_ (.A(_06838_),
    .Z(_06904_));
 NOR2_X1 _29369_ (.A1(_06826_),
    .A2(_06904_),
    .ZN(_06905_));
 BUF_X4 _29370_ (.A(_06905_),
    .Z(_06906_));
 AOI21_X1 _29371_ (.A(_06903_),
    .B1(_06906_),
    .B2(_06730_),
    .ZN(_06907_));
 OAI22_X4 _29372_ (.A1(_06777_),
    .A2(_06774_),
    .B1(_06834_),
    .B2(_06836_),
    .ZN(_06908_));
 BUF_X4 _29373_ (.A(_06908_),
    .Z(_06909_));
 NOR2_X4 _29374_ (.A1(_06818_),
    .A2(_06909_),
    .ZN(_06910_));
 NOR2_X1 _29375_ (.A1(_06899_),
    .A2(_06910_),
    .ZN(_06911_));
 NOR3_X1 _29376_ (.A1(_06808_),
    .A2(_06904_),
    .A3(_06885_),
    .ZN(_06912_));
 NAND2_X2 _29377_ (.A1(_06814_),
    .A2(_06767_),
    .ZN(_06913_));
 CLKBUF_X3 _29378_ (.A(_06818_),
    .Z(_06914_));
 OAI21_X1 _29379_ (.A(_06730_),
    .B1(_06913_),
    .B2(_06914_),
    .ZN(_06915_));
 OAI22_X1 _29380_ (.A1(_06730_),
    .A2(_06910_),
    .B1(_06912_),
    .B2(_06915_),
    .ZN(_06916_));
 AOI22_X1 _29381_ (.A1(_06907_),
    .A2(_06911_),
    .B1(_06916_),
    .B2(_06900_),
    .ZN(_06917_));
 OR3_X2 _29382_ (.A1(_06854_),
    .A2(_06901_),
    .A3(_06917_),
    .ZN(_06918_));
 BUF_X4 _29383_ (.A(_06757_),
    .Z(_06919_));
 OAI221_X2 _29384_ (.A(_06844_),
    .B1(_06830_),
    .B2(_06832_),
    .C1(_06919_),
    .C2(_06708_),
    .ZN(_06920_));
 BUF_X4 _29385_ (.A(_06920_),
    .Z(_06921_));
 BUF_X4 _29386_ (.A(_06921_),
    .Z(_06922_));
 NAND2_X4 _29387_ (.A1(_06858_),
    .A2(_06841_),
    .ZN(_06923_));
 NAND4_X4 _29388_ (.A1(_06843_),
    .A2(_06779_),
    .A3(_06865_),
    .A4(_06868_),
    .ZN(_06924_));
 NAND2_X2 _29389_ (.A1(_06923_),
    .A2(_06924_),
    .ZN(_06925_));
 NOR3_X1 _29390_ (.A1(_06902_),
    .A2(_06914_),
    .A3(_06925_),
    .ZN(_06926_));
 OAI21_X1 _29391_ (.A(_06874_),
    .B1(_06829_),
    .B2(_06926_),
    .ZN(_06927_));
 BUF_X4 _29392_ (.A(_06925_),
    .Z(_06928_));
 NOR3_X2 _29393_ (.A1(_06855_),
    .A2(_06759_),
    .A3(_06928_),
    .ZN(_06929_));
 NOR2_X1 _29394_ (.A1(_06827_),
    .A2(_06929_),
    .ZN(_06930_));
 AOI21_X1 _29395_ (.A(_06922_),
    .B1(_06927_),
    .B2(_06930_),
    .ZN(_06931_));
 NAND2_X4 _29396_ (.A1(_06821_),
    .A2(_06882_),
    .ZN(_06932_));
 NOR2_X1 _29397_ (.A1(_06730_),
    .A2(_06932_),
    .ZN(_06933_));
 BUF_X4 _29398_ (.A(_06822_),
    .Z(_06934_));
 OAI221_X2 _29399_ (.A(_06744_),
    .B1(_06836_),
    .B2(_06834_),
    .C1(_06756_),
    .C2(_06934_),
    .ZN(_06935_));
 BUF_X8 _29400_ (.A(_06810_),
    .Z(_06936_));
 AOI221_X2 _29401_ (.A(_06832_),
    .B1(_06811_),
    .B2(_06812_),
    .C1(_06936_),
    .C2(_06784_),
    .ZN(_06937_));
 BUF_X8 _29402_ (.A(_06810_),
    .Z(_06938_));
 AOI221_X2 _29403_ (.A(_06774_),
    .B1(_06794_),
    .B2(_06787_),
    .C1(_06775_),
    .C2(_06938_),
    .ZN(_06939_));
 OAI33_X1 _29404_ (.A1(_06852_),
    .A2(_06891_),
    .A3(_06904_),
    .B1(_06935_),
    .B2(_06937_),
    .B3(_06939_),
    .ZN(_06940_));
 NOR2_X2 _29405_ (.A1(_06815_),
    .A2(_06884_),
    .ZN(_06941_));
 OAI221_X2 _29406_ (.A(_06794_),
    .B1(_06728_),
    .B2(_06712_),
    .C1(_06783_),
    .C2(_06919_),
    .ZN(_06942_));
 BUF_X4 _29407_ (.A(_06942_),
    .Z(_06943_));
 NAND4_X4 _29408_ (.A1(_06799_),
    .A2(_06806_),
    .A3(_06923_),
    .A4(_06924_),
    .ZN(_06944_));
 NOR2_X4 _29409_ (.A1(_06943_),
    .A2(_06944_),
    .ZN(_06945_));
 OAI22_X4 _29410_ (.A1(_06849_),
    .A2(_06851_),
    .B1(_06860_),
    .B2(_06870_),
    .ZN(_06946_));
 NOR2_X4 _29411_ (.A1(_06921_),
    .A2(_06946_),
    .ZN(_06947_));
 AOI222_X2 _29412_ (.A1(_06933_),
    .A2(_06940_),
    .B1(_06941_),
    .B2(_06945_),
    .C1(_06947_),
    .C2(_06829_),
    .ZN(_06948_));
 NOR3_X1 _29413_ (.A1(_06921_),
    .A2(_06913_),
    .A3(_06884_),
    .ZN(_06949_));
 NOR2_X2 _29414_ (.A1(_06893_),
    .A2(_06807_),
    .ZN(_06950_));
 NAND4_X4 _29415_ (.A1(_06842_),
    .A2(_06844_),
    .A3(_06787_),
    .A4(_06845_),
    .ZN(_06951_));
 NOR3_X1 _29416_ (.A1(_06781_),
    .A2(_06826_),
    .A3(_06951_),
    .ZN(_06952_));
 BUF_X4 _29417_ (.A(_06806_),
    .Z(_06953_));
 OAI221_X2 _29418_ (.A(_06953_),
    .B1(_06860_),
    .B2(_06870_),
    .C1(_06886_),
    .C2(_06796_),
    .ZN(_06954_));
 BUF_X4 _29419_ (.A(_06954_),
    .Z(_06955_));
 AOI221_X2 _29420_ (.A(_06949_),
    .B1(_06839_),
    .B2(_06950_),
    .C1(_06952_),
    .C2(_06955_),
    .ZN(_06956_));
 NOR2_X4 _29421_ (.A1(_06730_),
    .A2(_06808_),
    .ZN(_06957_));
 NOR3_X1 _29422_ (.A1(_06898_),
    .A2(_06914_),
    .A3(_06904_),
    .ZN(_06958_));
 NOR3_X1 _29423_ (.A1(_06795_),
    .A2(_06902_),
    .A3(_06856_),
    .ZN(_06959_));
 OAI21_X1 _29424_ (.A(_06957_),
    .B1(_06958_),
    .B2(_06959_),
    .ZN(_06960_));
 NAND3_X1 _29425_ (.A1(_06948_),
    .A2(_06956_),
    .A3(_06960_),
    .ZN(_06961_));
 OAI22_X4 _29426_ (.A1(_06712_),
    .A2(_06727_),
    .B1(_06830_),
    .B2(_06832_),
    .ZN(_06962_));
 NOR4_X1 _29427_ (.A1(_06807_),
    .A2(_06815_),
    .A3(_06759_),
    .A4(_06962_),
    .ZN(_06963_));
 NOR2_X4 _29428_ (.A1(_06795_),
    .A2(_06852_),
    .ZN(_06964_));
 NOR3_X1 _29429_ (.A1(_06807_),
    .A2(_06781_),
    .A3(_06883_),
    .ZN(_06965_));
 AOI221_X1 _29430_ (.A(_06963_),
    .B1(_06964_),
    .B2(_06839_),
    .C1(_06846_),
    .C2(_06965_),
    .ZN(_06966_));
 OAI221_X2 _29431_ (.A(_06924_),
    .B1(_06851_),
    .B2(_06849_),
    .C1(_06859_),
    .C2(_06919_),
    .ZN(_06967_));
 BUF_X4 _29432_ (.A(_06967_),
    .Z(_06968_));
 NOR4_X2 _29433_ (.A1(_06893_),
    .A2(_06884_),
    .A3(_06908_),
    .A4(_06968_),
    .ZN(_06969_));
 OAI22_X1 _29434_ (.A1(_06893_),
    .A2(_06759_),
    .B1(_06826_),
    .B2(_06879_),
    .ZN(_06970_));
 BUF_X4 _29435_ (.A(_06895_),
    .Z(_06971_));
 AOI21_X1 _29436_ (.A(_06969_),
    .B1(_06970_),
    .B2(_06971_),
    .ZN(_06972_));
 NOR2_X4 _29437_ (.A1(_06884_),
    .A2(_06909_),
    .ZN(_06973_));
 BUF_X4 _29438_ (.A(_06946_),
    .Z(_06974_));
 NOR4_X1 _29439_ (.A1(_06730_),
    .A2(_06759_),
    .A3(_06974_),
    .A4(_06909_),
    .ZN(_06975_));
 OAI21_X1 _29440_ (.A(_06899_),
    .B1(_06973_),
    .B2(_06975_),
    .ZN(_06976_));
 NOR2_X2 _29441_ (.A1(_06824_),
    .A2(_06757_),
    .ZN(_06977_));
 NOR4_X2 _29442_ (.A1(_06777_),
    .A2(_06774_),
    .A3(_06755_),
    .A4(_06977_),
    .ZN(_06978_));
 NAND4_X2 _29443_ (.A1(_06799_),
    .A2(_06953_),
    .A3(_06811_),
    .A4(_06812_),
    .ZN(_06979_));
 OR2_X2 _29444_ (.A1(_00354_),
    .A2(_06820_),
    .ZN(_06980_));
 NAND2_X1 _29445_ (.A1(_06821_),
    .A2(_06980_),
    .ZN(_06981_));
 AOI21_X1 _29446_ (.A(_06978_),
    .B1(_06979_),
    .B2(_06981_),
    .ZN(_06982_));
 OR4_X1 _29447_ (.A1(_06893_),
    .A2(_06879_),
    .A3(_06891_),
    .A4(_06982_),
    .ZN(_06983_));
 NAND4_X1 _29448_ (.A1(_06966_),
    .A2(_06972_),
    .A3(_06976_),
    .A4(_06983_),
    .ZN(_06984_));
 NOR2_X4 _29449_ (.A1(_06781_),
    .A2(_06883_),
    .ZN(_06985_));
 NOR2_X1 _29450_ (.A1(_06807_),
    .A2(_06815_),
    .ZN(_06986_));
 AOI221_X2 _29451_ (.A(_06816_),
    .B1(_06980_),
    .B2(_06821_),
    .C1(\core.keymem.prev_key1_reg[7] ),
    .C2(_06936_),
    .ZN(_06987_));
 AOI221_X2 _29452_ (.A(_06795_),
    .B1(_06807_),
    .B2(_06985_),
    .C1(_06986_),
    .C2(_06987_),
    .ZN(_06988_));
 NOR2_X4 _29453_ (.A1(_06759_),
    .A2(_06904_),
    .ZN(_06989_));
 OAI21_X2 _29454_ (.A(_06730_),
    .B1(_06898_),
    .B2(_06989_),
    .ZN(_06990_));
 NOR2_X4 _29455_ (.A1(_06781_),
    .A2(_06818_),
    .ZN(_06991_));
 AOI21_X2 _29456_ (.A(_06991_),
    .B1(_06941_),
    .B2(_06944_),
    .ZN(_06992_));
 OAI22_X4 _29457_ (.A1(_06988_),
    .A2(_06990_),
    .B1(_06992_),
    .B2(_06943_),
    .ZN(_06993_));
 OR4_X2 _29458_ (.A1(_06931_),
    .A2(_06961_),
    .A3(_06984_),
    .A4(_06993_),
    .ZN(_06994_));
 NOR3_X2 _29459_ (.A1(_06852_),
    .A2(_06902_),
    .A3(_06856_),
    .ZN(_06995_));
 NOR3_X2 _29460_ (.A1(_06808_),
    .A2(_06876_),
    .A3(_06909_),
    .ZN(_06996_));
 OAI21_X1 _29461_ (.A(_06899_),
    .B1(_06995_),
    .B2(_06996_),
    .ZN(_06997_));
 NOR3_X1 _29462_ (.A1(_06898_),
    .A2(_06904_),
    .A3(_06884_),
    .ZN(_06998_));
 NOR2_X4 _29463_ (.A1(_06759_),
    .A2(_06908_),
    .ZN(_06999_));
 AOI221_X2 _29464_ (.A(_06870_),
    .B1(_06806_),
    .B2(_06798_),
    .C1(_06858_),
    .C2(_06938_),
    .ZN(_07000_));
 BUF_X4 _29465_ (.A(_07000_),
    .Z(_07001_));
 AOI221_X2 _29466_ (.A(_06998_),
    .B1(_06999_),
    .B2(_07001_),
    .C1(_06898_),
    .C2(_06829_),
    .ZN(_07002_));
 AOI21_X2 _29467_ (.A(_06731_),
    .B1(_06997_),
    .B2(_07002_),
    .ZN(_07003_));
 BUF_X4 _29468_ (.A(_06951_),
    .Z(_07004_));
 BUF_X4 _29469_ (.A(_06941_),
    .Z(_07005_));
 NAND2_X2 _29470_ (.A1(_07005_),
    .A2(_06944_),
    .ZN(_07006_));
 NOR2_X1 _29471_ (.A1(_06893_),
    .A2(_07001_),
    .ZN(_07007_));
 AOI22_X4 _29472_ (.A1(_06894_),
    .A2(_06999_),
    .B1(_07007_),
    .B2(_06973_),
    .ZN(_07008_));
 OAI22_X4 _29473_ (.A1(_07004_),
    .A2(_07006_),
    .B1(_07008_),
    .B2(_06899_),
    .ZN(_07009_));
 OR2_X2 _29474_ (.A1(_07003_),
    .A2(_07009_),
    .ZN(_07010_));
 NOR2_X4 _29475_ (.A1(_06777_),
    .A2(_06774_),
    .ZN(_07011_));
 NAND2_X1 _29476_ (.A1(_07011_),
    .A2(_06981_),
    .ZN(_07012_));
 OAI21_X1 _29477_ (.A(_06935_),
    .B1(_06891_),
    .B2(_06913_),
    .ZN(_07013_));
 NAND3_X1 _29478_ (.A1(_06898_),
    .A2(_06852_),
    .A3(_06880_),
    .ZN(_07014_));
 NAND2_X1 _29479_ (.A1(_07013_),
    .A2(_07014_),
    .ZN(_07015_));
 OAI221_X2 _29480_ (.A(_06845_),
    .B1(_06849_),
    .B2(_06851_),
    .C1(_06887_),
    .C2(_06783_),
    .ZN(_07016_));
 BUF_X4 _29481_ (.A(_07016_),
    .Z(_07017_));
 NOR2_X1 _29482_ (.A1(_06880_),
    .A2(_07017_),
    .ZN(_07018_));
 NOR4_X1 _29483_ (.A1(_06731_),
    .A2(_07012_),
    .A3(_07015_),
    .A4(_07018_),
    .ZN(_07019_));
 NOR4_X4 _29484_ (.A1(_06849_),
    .A2(_06851_),
    .A3(_06860_),
    .A4(_06870_),
    .ZN(_07020_));
 NOR2_X1 _29485_ (.A1(_06921_),
    .A2(_07020_),
    .ZN(_07021_));
 AOI22_X2 _29486_ (.A1(_07005_),
    .A2(_06846_),
    .B1(_07021_),
    .B2(_06991_),
    .ZN(_07022_));
 NOR2_X4 _29487_ (.A1(_06904_),
    .A2(_06884_),
    .ZN(_07023_));
 AOI21_X1 _29488_ (.A(_06965_),
    .B1(_07023_),
    .B2(_06808_),
    .ZN(_07024_));
 NAND2_X2 _29489_ (.A1(_06744_),
    .A2(_06881_),
    .ZN(_07025_));
 MUX2_X1 _29490_ (.A(_07025_),
    .B(_06890_),
    .S(_06852_),
    .Z(_07026_));
 OR3_X1 _29491_ (.A1(_06879_),
    .A2(_07012_),
    .A3(_07026_),
    .ZN(_07027_));
 BUF_X4 _29492_ (.A(_06943_),
    .Z(_07028_));
 OAI221_X2 _29493_ (.A(_07022_),
    .B1(_07024_),
    .B2(_07004_),
    .C1(_07027_),
    .C2(_07028_),
    .ZN(_07029_));
 NOR2_X4 _29494_ (.A1(_06955_),
    .A2(_06951_),
    .ZN(_07030_));
 AOI222_X2 _29495_ (.A1(_06787_),
    .A2(_06845_),
    .B1(_06811_),
    .B2(_06812_),
    .C1(_06821_),
    .C2(_06980_),
    .ZN(_07031_));
 MUX2_X1 _29496_ (.A(_06978_),
    .B(_07031_),
    .S(_06879_),
    .Z(_07032_));
 NOR3_X1 _29497_ (.A1(_06729_),
    .A2(_06808_),
    .A3(_06891_),
    .ZN(_07033_));
 NOR2_X1 _29498_ (.A1(_06795_),
    .A2(_07025_),
    .ZN(_07034_));
 NOR2_X4 _29499_ (.A1(_06755_),
    .A2(_06746_),
    .ZN(_07035_));
 OAI221_X1 _29500_ (.A(_06767_),
    .B1(_06728_),
    .B2(_06712_),
    .C1(_06778_),
    .C2(_06886_),
    .ZN(_07036_));
 OAI33_X1 _29501_ (.A1(_06893_),
    .A2(_07035_),
    .A3(_06838_),
    .B1(_07036_),
    .B2(_06932_),
    .B3(_07011_),
    .ZN(_07037_));
 AOI222_X2 _29502_ (.A1(_06827_),
    .A2(_07030_),
    .B1(_07032_),
    .B2(_07033_),
    .C1(_07034_),
    .C2(_07037_),
    .ZN(_07038_));
 NOR3_X2 _29503_ (.A1(_06815_),
    .A2(_06925_),
    .A3(_06826_),
    .ZN(_07039_));
 OAI22_X1 _29504_ (.A1(_06902_),
    .A2(_06914_),
    .B1(_06826_),
    .B2(_06815_),
    .ZN(_07040_));
 AOI22_X1 _29505_ (.A1(_06833_),
    .A2(_07039_),
    .B1(_07040_),
    .B2(_06846_),
    .ZN(_07041_));
 OAI21_X1 _29506_ (.A(_07038_),
    .B1(_07041_),
    .B2(_06853_),
    .ZN(_07042_));
 OR3_X2 _29507_ (.A1(_07019_),
    .A2(_07029_),
    .A3(_07042_),
    .ZN(_07043_));
 NOR4_X4 _29508_ (.A1(_06918_),
    .A2(_06994_),
    .A3(_07010_),
    .A4(_07043_),
    .ZN(_07044_));
 BUF_X4 _29509_ (.A(_06910_),
    .Z(_07045_));
 BUF_X4 _29510_ (.A(_06944_),
    .Z(_07046_));
 NOR2_X2 _29511_ (.A1(_07046_),
    .A2(_06962_),
    .ZN(_07047_));
 NOR2_X4 _29512_ (.A1(_06943_),
    .A2(_06955_),
    .ZN(_07048_));
 AOI222_X2 _29513_ (.A1(_07045_),
    .A2(_07030_),
    .B1(_07047_),
    .B2(_07023_),
    .C1(_07048_),
    .C2(_06857_),
    .ZN(_07049_));
 BUF_X4 _29514_ (.A(_06876_),
    .Z(_07050_));
 BUF_X4 _29515_ (.A(_06955_),
    .Z(_07051_));
 BUF_X4 _29516_ (.A(_06909_),
    .Z(_07052_));
 CLKBUF_X3 _29517_ (.A(_07052_),
    .Z(_07053_));
 NOR3_X1 _29518_ (.A1(_07050_),
    .A2(_07051_),
    .A3(_07053_),
    .ZN(_07054_));
 NOR2_X4 _29519_ (.A1(_06856_),
    .A2(_07052_),
    .ZN(_07055_));
 AOI21_X1 _29520_ (.A(_07054_),
    .B1(_07055_),
    .B2(_07051_),
    .ZN(_07056_));
 BUF_X4 _29521_ (.A(_06795_),
    .Z(_07057_));
 BUF_X4 _29522_ (.A(_07057_),
    .Z(_07058_));
 BUF_X4 _29523_ (.A(_06928_),
    .Z(_07059_));
 BUF_X4 _29524_ (.A(_07059_),
    .Z(_07060_));
 BUF_X4 _29525_ (.A(_06874_),
    .Z(_07061_));
 BUF_X4 _29526_ (.A(_07061_),
    .Z(_07062_));
 BUF_X4 _29527_ (.A(_06855_),
    .Z(_07063_));
 OAI21_X1 _29528_ (.A(_07062_),
    .B1(_07063_),
    .B2(_07050_),
    .ZN(_07064_));
 AOI21_X1 _29529_ (.A(_07058_),
    .B1(_07060_),
    .B2(_07064_),
    .ZN(_07065_));
 BUF_X4 _29530_ (.A(_06894_),
    .Z(_07066_));
 BUF_X4 _29531_ (.A(_07066_),
    .Z(_07067_));
 BUF_X4 _29532_ (.A(_06899_),
    .Z(_07068_));
 BUF_X4 _29533_ (.A(_07068_),
    .Z(_07069_));
 BUF_X4 _29534_ (.A(_06909_),
    .Z(_07070_));
 NOR3_X2 _29535_ (.A1(_07050_),
    .A2(_07020_),
    .A3(_07070_),
    .ZN(_07071_));
 OAI221_X2 _29536_ (.A(_07067_),
    .B1(_07069_),
    .B2(_06974_),
    .C1(_07071_),
    .C2(_06829_),
    .ZN(_07072_));
 OAI221_X2 _29537_ (.A(_07049_),
    .B1(_07056_),
    .B2(_07004_),
    .C1(_07065_),
    .C2(_07072_),
    .ZN(_07073_));
 BUF_X4 _29538_ (.A(_07001_),
    .Z(_07074_));
 OAI21_X2 _29539_ (.A(_07051_),
    .B1(_07074_),
    .B2(_07068_),
    .ZN(_07075_));
 BUF_X4 _29540_ (.A(_06731_),
    .Z(_07076_));
 BUF_X4 _29541_ (.A(_06856_),
    .Z(_07077_));
 CLKBUF_X3 _29542_ (.A(_07077_),
    .Z(_07078_));
 BUF_X4 _29543_ (.A(_06904_),
    .Z(_07079_));
 BUF_X4 _29544_ (.A(_07079_),
    .Z(_07080_));
 NOR3_X2 _29545_ (.A1(_07076_),
    .A2(_07078_),
    .A3(_07080_),
    .ZN(_07081_));
 NOR2_X4 _29546_ (.A1(_06974_),
    .A2(_06951_),
    .ZN(_07082_));
 BUF_X8 _29547_ (.A(_06989_),
    .Z(_07083_));
 AOI22_X4 _29548_ (.A1(_07075_),
    .A2(_07081_),
    .B1(_07082_),
    .B2(_07083_),
    .ZN(_07084_));
 BUF_X4 _29549_ (.A(_07076_),
    .Z(_07085_));
 BUF_X4 _29550_ (.A(_07057_),
    .Z(_07086_));
 BUF_X4 _29551_ (.A(_06885_),
    .Z(_07087_));
 AOI22_X4 _29552_ (.A1(_06799_),
    .A2(_06953_),
    .B1(_06923_),
    .B2(_06924_),
    .ZN(_07088_));
 NOR4_X2 _29553_ (.A1(_07086_),
    .A2(_07079_),
    .A3(_07087_),
    .A4(_07088_),
    .ZN(_07089_));
 BUF_X4 _29554_ (.A(_06876_),
    .Z(_07090_));
 BUF_X4 _29555_ (.A(_06902_),
    .Z(_07091_));
 CLKBUF_X3 _29556_ (.A(_07091_),
    .Z(_07092_));
 BUF_X4 _29557_ (.A(_06968_),
    .Z(_07093_));
 NOR4_X2 _29558_ (.A1(_06900_),
    .A2(_07090_),
    .A3(_07092_),
    .A4(_07093_),
    .ZN(_07094_));
 OAI21_X2 _29559_ (.A(_07085_),
    .B1(_07089_),
    .B2(_07094_),
    .ZN(_07095_));
 NOR3_X2 _29560_ (.A1(_07061_),
    .A2(_07063_),
    .A3(_07078_),
    .ZN(_07096_));
 BUF_X4 _29561_ (.A(_06914_),
    .Z(_07097_));
 BUF_X4 _29562_ (.A(_07097_),
    .Z(_07098_));
 CLKBUF_X3 _29563_ (.A(_07098_),
    .Z(_07099_));
 OAI22_X1 _29564_ (.A1(_07063_),
    .A2(_07078_),
    .B1(_07080_),
    .B2(_07099_),
    .ZN(_07100_));
 AOI21_X2 _29565_ (.A(_07096_),
    .B1(_07100_),
    .B2(_07060_),
    .ZN(_07101_));
 BUF_X4 _29566_ (.A(_06962_),
    .Z(_07102_));
 OAI211_X4 _29567_ (.A(_07084_),
    .B(_07095_),
    .C1(_07101_),
    .C2(_07102_),
    .ZN(_07103_));
 BUF_X4 _29568_ (.A(_06808_),
    .Z(_07104_));
 BUF_X4 _29569_ (.A(_07104_),
    .Z(_07105_));
 BUF_X4 _29570_ (.A(_07105_),
    .Z(_07106_));
 CLKBUF_X3 _29571_ (.A(_06885_),
    .Z(_07107_));
 BUF_X4 _29572_ (.A(_06936_),
    .Z(_07108_));
 BUF_X4 _29573_ (.A(_07108_),
    .Z(_07109_));
 AOI221_X2 _29574_ (.A(_06728_),
    .B1(_06923_),
    .B2(_06924_),
    .C1(_07109_),
    .C2(_06840_),
    .ZN(_07110_));
 OAI33_X1 _29575_ (.A1(_07076_),
    .A2(_07092_),
    .A3(_07078_),
    .B1(_07079_),
    .B2(_07107_),
    .B3(_07110_),
    .ZN(_07111_));
 BUF_X4 _29576_ (.A(_07066_),
    .Z(_07112_));
 NOR2_X1 _29577_ (.A1(_07112_),
    .A2(_07051_),
    .ZN(_07113_));
 AOI22_X2 _29578_ (.A1(_07106_),
    .A2(_07111_),
    .B1(_07113_),
    .B2(_07023_),
    .ZN(_07114_));
 NOR2_X1 _29579_ (.A1(_07069_),
    .A2(_07114_),
    .ZN(_07115_));
 NOR3_X2 _29580_ (.A1(_06993_),
    .A2(_07103_),
    .A3(_07115_),
    .ZN(_07116_));
 NOR3_X4 _29581_ (.A1(_06871_),
    .A2(_06826_),
    .A3(_06909_),
    .ZN(_07117_));
 AOI221_X2 _29582_ (.A(_07117_),
    .B1(_06985_),
    .B2(_06872_),
    .C1(_06799_),
    .C2(_06953_),
    .ZN(_07118_));
 BUF_X4 _29583_ (.A(_06872_),
    .Z(_07119_));
 BUF_X4 _29584_ (.A(_07119_),
    .Z(_07120_));
 AOI21_X1 _29585_ (.A(_07105_),
    .B1(_07120_),
    .B2(_07045_),
    .ZN(_07121_));
 AOI221_X2 _29586_ (.A(_06836_),
    .B1(_06812_),
    .B2(_06811_),
    .C1(_06813_),
    .C2(_07108_),
    .ZN(_07122_));
 OR2_X2 _29587_ (.A1(_00357_),
    .A2(_06886_),
    .ZN(_07123_));
 AOI22_X4 _29588_ (.A1(_06821_),
    .A2(_06980_),
    .B1(_06744_),
    .B2(_07123_),
    .ZN(_07124_));
 NOR2_X2 _29589_ (.A1(_06756_),
    .A2(_06886_),
    .ZN(_07125_));
 NOR4_X4 _29590_ (.A1(_06755_),
    .A2(_06816_),
    .A3(_07125_),
    .A4(_06977_),
    .ZN(_07126_));
 AOI22_X1 _29591_ (.A1(_07122_),
    .A2(_07124_),
    .B1(_07126_),
    .B2(_06880_),
    .ZN(_07127_));
 NOR4_X4 _29592_ (.A1(_06777_),
    .A2(_06774_),
    .A3(_06834_),
    .A4(_06836_),
    .ZN(_07128_));
 BUF_X4 _29593_ (.A(_06987_),
    .Z(_07129_));
 AOI221_X2 _29594_ (.A(_06755_),
    .B1(_06744_),
    .B2(_07123_),
    .C1(_07109_),
    .C2(_06823_),
    .ZN(_07130_));
 CLKBUF_X3 _29595_ (.A(_06913_),
    .Z(_07131_));
 AOI22_X1 _29596_ (.A1(_07128_),
    .A2(_07129_),
    .B1(_07130_),
    .B2(_07131_),
    .ZN(_07132_));
 MUX2_X1 _29597_ (.A(_07127_),
    .B(_07132_),
    .S(_07119_),
    .Z(_07133_));
 AOI211_X2 _29598_ (.A(_06922_),
    .B(_07118_),
    .C1(_07121_),
    .C2(_07133_),
    .ZN(_07134_));
 NOR3_X2 _29599_ (.A1(_06876_),
    .A2(_06872_),
    .A3(_06909_),
    .ZN(_07135_));
 AOI221_X2 _29600_ (.A(_07135_),
    .B1(_06827_),
    .B2(_07119_),
    .C1(_06799_),
    .C2(_06953_),
    .ZN(_07136_));
 BUF_X4 _29601_ (.A(_07104_),
    .Z(_07137_));
 BUF_X4 _29602_ (.A(_06827_),
    .Z(_07138_));
 AOI21_X1 _29603_ (.A(_07137_),
    .B1(_07060_),
    .B2(_07138_),
    .ZN(_07139_));
 BUF_X4 _29604_ (.A(_06904_),
    .Z(_07140_));
 NOR4_X2 _29605_ (.A1(_06894_),
    .A2(_06874_),
    .A3(_07097_),
    .A4(_07140_),
    .ZN(_07141_));
 OAI33_X1 _29606_ (.A1(_07035_),
    .A2(_07025_),
    .A3(_07091_),
    .B1(_07098_),
    .B2(_07104_),
    .B3(_06855_),
    .ZN(_07142_));
 AOI21_X1 _29607_ (.A(_07141_),
    .B1(_07142_),
    .B2(_07112_),
    .ZN(_07143_));
 BUF_X4 _29608_ (.A(_07120_),
    .Z(_07144_));
 OAI33_X1 _29609_ (.A1(_07004_),
    .A2(_07136_),
    .A3(_07139_),
    .B1(_07143_),
    .B2(_07058_),
    .B3(_07144_),
    .ZN(_07145_));
 BUF_X4 _29610_ (.A(_06782_),
    .Z(_07146_));
 NOR2_X4 _29611_ (.A1(_06962_),
    .A2(_06968_),
    .ZN(_07147_));
 NOR3_X2 _29612_ (.A1(_06894_),
    .A2(_06855_),
    .A3(_06856_),
    .ZN(_07148_));
 XNOR2_X1 _29613_ (.A(_06899_),
    .B(_07001_),
    .ZN(_07149_));
 AOI222_X2 _29614_ (.A1(_06947_),
    .A2(_07146_),
    .B1(_07083_),
    .B2(_07147_),
    .C1(_07148_),
    .C2(_07149_),
    .ZN(_07150_));
 NOR2_X4 _29615_ (.A1(_06943_),
    .A2(_06974_),
    .ZN(_07151_));
 NOR2_X2 _29616_ (.A1(_06944_),
    .A2(_07004_),
    .ZN(_07152_));
 NOR4_X4 _29617_ (.A1(_07090_),
    .A2(_06944_),
    .A3(_07004_),
    .A4(_07052_),
    .ZN(_07153_));
 OAI22_X2 _29618_ (.A1(_07151_),
    .A2(_07152_),
    .B1(_07153_),
    .B2(_06857_),
    .ZN(_07154_));
 BUF_X4 _29619_ (.A(_06833_),
    .Z(_07155_));
 NOR3_X4 _29620_ (.A1(_06871_),
    .A2(_06884_),
    .A3(_06908_),
    .ZN(_07156_));
 NOR3_X1 _29621_ (.A1(_07098_),
    .A2(_07079_),
    .A3(_07046_),
    .ZN(_07157_));
 OAI21_X1 _29622_ (.A(_07155_),
    .B1(_07156_),
    .B2(_07157_),
    .ZN(_07158_));
 BUF_X4 _29623_ (.A(_06819_),
    .Z(_07159_));
 AOI22_X4 _29624_ (.A1(_07045_),
    .A2(_07147_),
    .B1(_07151_),
    .B2(_07159_),
    .ZN(_07160_));
 NAND4_X2 _29625_ (.A1(_07150_),
    .A2(_07154_),
    .A3(_07158_),
    .A4(_07160_),
    .ZN(_07161_));
 NOR2_X4 _29626_ (.A1(_06731_),
    .A2(_07057_),
    .ZN(_07162_));
 NOR3_X1 _29627_ (.A1(_07080_),
    .A2(_07107_),
    .A3(_07020_),
    .ZN(_07163_));
 AOI221_X2 _29628_ (.A(_06851_),
    .B1(_06923_),
    .B2(_06924_),
    .C1(_07108_),
    .C2(_06797_),
    .ZN(_07164_));
 BUF_X4 _29629_ (.A(_07164_),
    .Z(_07165_));
 NOR3_X1 _29630_ (.A1(_07098_),
    .A2(_07079_),
    .A3(_07165_),
    .ZN(_07166_));
 OAI21_X1 _29631_ (.A(_07162_),
    .B1(_07163_),
    .B2(_07166_),
    .ZN(_07167_));
 NOR2_X4 _29632_ (.A1(_06893_),
    .A2(_06898_),
    .ZN(_07168_));
 NAND3_X1 _29633_ (.A1(_07168_),
    .A2(_07165_),
    .A3(_07055_),
    .ZN(_07169_));
 NAND2_X1 _29634_ (.A1(_07167_),
    .A2(_07169_),
    .ZN(_07170_));
 NOR4_X4 _29635_ (.A1(_07134_),
    .A2(_07145_),
    .A3(_07161_),
    .A4(_07170_),
    .ZN(_07171_));
 NOR2_X4 _29636_ (.A1(_06921_),
    .A2(_06808_),
    .ZN(_07172_));
 AND2_X1 _29637_ (.A1(_06839_),
    .A2(_07172_),
    .ZN(_07173_));
 NOR3_X1 _29638_ (.A1(_06914_),
    .A2(_06951_),
    .A3(_06909_),
    .ZN(_07174_));
 NOR4_X1 _29639_ (.A1(_06855_),
    .A2(_06928_),
    .A3(_06885_),
    .A4(_06962_),
    .ZN(_07175_));
 NOR4_X1 _29640_ (.A1(_06902_),
    .A2(_06872_),
    .A3(_06884_),
    .A4(_06943_),
    .ZN(_07176_));
 OR3_X1 _29641_ (.A1(_07174_),
    .A2(_07175_),
    .A3(_07176_),
    .ZN(_07177_));
 BUF_X4 _29642_ (.A(_06985_),
    .Z(_07178_));
 AOI221_X2 _29643_ (.A(_07173_),
    .B1(_07177_),
    .B2(_07105_),
    .C1(_06945_),
    .C2(_07178_),
    .ZN(_07179_));
 MUX2_X1 _29644_ (.A(_07092_),
    .B(_07079_),
    .S(_07066_),
    .Z(_07180_));
 NAND3_X2 _29645_ (.A1(_07068_),
    .A2(_07129_),
    .A3(_07093_),
    .ZN(_07181_));
 NOR2_X1 _29646_ (.A1(_07180_),
    .A2(_07181_),
    .ZN(_07182_));
 NOR2_X1 _29647_ (.A1(_07068_),
    .A2(_07120_),
    .ZN(_07183_));
 AOI22_X4 _29648_ (.A1(_06811_),
    .A2(_06812_),
    .B1(_06814_),
    .B2(_06767_),
    .ZN(_07184_));
 NAND4_X1 _29649_ (.A1(_07076_),
    .A2(_07137_),
    .A3(_07129_),
    .A4(_07184_),
    .ZN(_07185_));
 NAND2_X2 _29650_ (.A1(_06894_),
    .A2(_06874_),
    .ZN(_07186_));
 NAND2_X2 _29651_ (.A1(_07122_),
    .A2(_07124_),
    .ZN(_07187_));
 OAI21_X1 _29652_ (.A(_07185_),
    .B1(_07186_),
    .B2(_07187_),
    .ZN(_07188_));
 AOI21_X1 _29653_ (.A(_07182_),
    .B1(_07183_),
    .B2(_07188_),
    .ZN(_07189_));
 NOR3_X1 _29654_ (.A1(_07076_),
    .A2(_07098_),
    .A3(_07053_),
    .ZN(_07190_));
 OAI22_X2 _29655_ (.A1(_06849_),
    .A2(_06851_),
    .B1(_06816_),
    .B2(_06817_),
    .ZN(_07191_));
 NOR4_X2 _29656_ (.A1(_07066_),
    .A2(_07059_),
    .A3(_07191_),
    .A4(_06889_),
    .ZN(_07192_));
 OAI21_X1 _29657_ (.A(_07068_),
    .B1(_07190_),
    .B2(_07192_),
    .ZN(_07193_));
 NAND3_X1 _29658_ (.A1(_07062_),
    .A2(_06847_),
    .A3(_06973_),
    .ZN(_07194_));
 NOR2_X2 _29659_ (.A1(_07061_),
    .A2(_07004_),
    .ZN(_07195_));
 NOR3_X1 _29660_ (.A1(_07059_),
    .A2(_07087_),
    .A3(_07070_),
    .ZN(_07196_));
 OAI21_X2 _29661_ (.A(_07195_),
    .B1(_07196_),
    .B2(_07005_),
    .ZN(_07197_));
 AND3_X1 _29662_ (.A1(_07193_),
    .A2(_07194_),
    .A3(_07197_),
    .ZN(_07198_));
 NAND4_X1 _29663_ (.A1(_07129_),
    .A2(_07122_),
    .A3(_07088_),
    .A4(_06847_),
    .ZN(_07199_));
 AOI22_X4 _29664_ (.A1(_06787_),
    .A2(_06845_),
    .B1(_06799_),
    .B2(_06953_),
    .ZN(_07200_));
 AOI22_X4 _29665_ (.A1(_06842_),
    .A2(_06844_),
    .B1(_06923_),
    .B2(_06924_),
    .ZN(_07201_));
 NOR4_X4 _29666_ (.A1(_06712_),
    .A2(_06728_),
    .A3(_06860_),
    .A4(_06870_),
    .ZN(_07202_));
 OAI21_X2 _29667_ (.A(_07200_),
    .B1(_07201_),
    .B2(_07202_),
    .ZN(_07203_));
 NAND2_X4 _29668_ (.A1(_07126_),
    .A2(_07184_),
    .ZN(_07204_));
 OR2_X1 _29669_ (.A1(_06876_),
    .A2(_07140_),
    .ZN(_07205_));
 NAND2_X1 _29670_ (.A1(_07165_),
    .A2(_06833_),
    .ZN(_07206_));
 OAI221_X2 _29671_ (.A(_07199_),
    .B1(_07203_),
    .B2(_07204_),
    .C1(_07205_),
    .C2(_07206_),
    .ZN(_07207_));
 NAND2_X2 _29672_ (.A1(_07128_),
    .A2(_07126_),
    .ZN(_07208_));
 MUX2_X1 _29673_ (.A(_07025_),
    .B(_06891_),
    .S(_06795_),
    .Z(_07209_));
 NAND2_X1 _29674_ (.A1(_06874_),
    .A2(_06971_),
    .ZN(_07210_));
 NOR2_X1 _29675_ (.A1(_06755_),
    .A2(_06977_),
    .ZN(_07211_));
 NAND4_X1 _29676_ (.A1(_06893_),
    .A2(_07131_),
    .A3(_06872_),
    .A4(_07211_),
    .ZN(_07212_));
 OAI33_X1 _29677_ (.A1(_06922_),
    .A2(_06853_),
    .A3(_07208_),
    .B1(_07209_),
    .B2(_07210_),
    .B3(_07212_),
    .ZN(_07213_));
 NAND2_X1 _29678_ (.A1(_06880_),
    .A2(_07124_),
    .ZN(_07214_));
 AND2_X1 _29679_ (.A1(_07093_),
    .A2(_06979_),
    .ZN(_07215_));
 OAI221_X2 _29680_ (.A(_07066_),
    .B1(_07208_),
    .B2(_07051_),
    .C1(_07214_),
    .C2(_07215_),
    .ZN(_07216_));
 NAND3_X1 _29681_ (.A1(_07129_),
    .A2(_07165_),
    .A3(_07184_),
    .ZN(_07217_));
 AOI21_X1 _29682_ (.A(_06900_),
    .B1(_07217_),
    .B2(_06731_),
    .ZN(_07218_));
 AOI211_X2 _29683_ (.A(_07207_),
    .B(_07213_),
    .C1(_07216_),
    .C2(_07218_),
    .ZN(_07219_));
 AND4_X1 _29684_ (.A1(_07179_),
    .A2(_07189_),
    .A3(_07198_),
    .A4(_07219_),
    .ZN(_07220_));
 NAND3_X2 _29685_ (.A1(_07116_),
    .A2(_07171_),
    .A3(_07220_),
    .ZN(_07221_));
 NOR3_X4 _29686_ (.A1(_07044_),
    .A2(_07073_),
    .A3(_07221_),
    .ZN(_07222_));
 OR2_X2 _29687_ (.A1(_06707_),
    .A2(_07222_),
    .ZN(_07223_));
 CLKBUF_X3 _29688_ (.A(_06703_),
    .Z(_07224_));
 NAND3_X1 _29689_ (.A1(_16240_),
    .A2(_06694_),
    .A3(_16246_),
    .ZN(_07225_));
 OR2_X1 _29690_ (.A1(_16235_),
    .A2(_06691_),
    .ZN(_07226_));
 NAND2_X2 _29691_ (.A1(_07225_),
    .A2(_07226_),
    .ZN(_07227_));
 CLKBUF_X3 _29692_ (.A(_07227_),
    .Z(_07228_));
 CLKBUF_X3 _29693_ (.A(_07228_),
    .Z(_07229_));
 NAND3_X1 _29694_ (.A1(_16239_),
    .A2(_06690_),
    .A3(_16238_),
    .ZN(_07230_));
 BUF_X4 _29695_ (.A(_07230_),
    .Z(_07231_));
 BUF_X4 _29696_ (.A(_07231_),
    .Z(_07232_));
 NOR2_X1 _29697_ (.A1(\core.enc_block.block_w3_reg[0] ),
    .A2(_07232_),
    .ZN(_07233_));
 CLKBUF_X3 _29698_ (.A(\core.enc_block.block_w0_reg[24] ),
    .Z(_07234_));
 BUF_X4 _29699_ (.A(\core.enc_block.block_w0_reg[31] ),
    .Z(_07235_));
 XNOR2_X2 _29700_ (.A(_07234_),
    .B(_07235_),
    .ZN(_07236_));
 CLKBUF_X3 _29701_ (.A(\core.enc_block.block_w2_reg[8] ),
    .Z(_07237_));
 CLKBUF_X3 _29702_ (.A(\core.enc_block.block_w1_reg[16] ),
    .Z(_07238_));
 XNOR2_X1 _29703_ (.A(_07237_),
    .B(_07238_),
    .ZN(_07239_));
 XNOR2_X1 _29704_ (.A(_07236_),
    .B(_07239_),
    .ZN(_07240_));
 XNOR2_X1 _29705_ (.A(_06742_),
    .B(_07240_),
    .ZN(_07241_));
 BUF_X4 _29706_ (.A(_07231_),
    .Z(_07242_));
 BUF_X4 _29707_ (.A(_07242_),
    .Z(_07243_));
 AOI21_X2 _29708_ (.A(_07233_),
    .B1(_07241_),
    .B2(_07243_),
    .ZN(_07244_));
 NAND2_X1 _29709_ (.A1(_07229_),
    .A2(_07244_),
    .ZN(_07245_));
 NAND3_X4 _29710_ (.A1(_16235_),
    .A2(_16239_),
    .A3(_06694_),
    .ZN(_07246_));
 CLKBUF_X3 _29711_ (.A(_07246_),
    .Z(_07247_));
 BUF_X4 _29712_ (.A(_07247_),
    .Z(_07248_));
 INV_X1 _29713_ (.A(\block_reg[0][0] ),
    .ZN(_07249_));
 OAI21_X1 _29714_ (.A(_07245_),
    .B1(_07248_),
    .B2(_07249_),
    .ZN(_07250_));
 BUF_X4 _29715_ (.A(_07247_),
    .Z(_07251_));
 AND2_X1 _29716_ (.A1(_07225_),
    .A2(_07226_),
    .ZN(_07252_));
 CLKBUF_X3 _29717_ (.A(_07252_),
    .Z(_07253_));
 CLKBUF_X3 _29718_ (.A(_07253_),
    .Z(_07254_));
 OAI22_X1 _29719_ (.A1(\block_reg[0][0] ),
    .A2(_07251_),
    .B1(_07254_),
    .B2(_07244_),
    .ZN(_07255_));
 MUX2_X1 _29720_ (.A(_07250_),
    .B(_07255_),
    .S(_16550_),
    .Z(_07256_));
 NOR2_X1 _29721_ (.A1(_07224_),
    .A2(_07256_),
    .ZN(_07257_));
 AOI22_X1 _29722_ (.A1(_06689_),
    .A2(_06705_),
    .B1(_07223_),
    .B2(_07257_),
    .ZN(_00702_));
 BUF_X2 _29723_ (.A(\core.enc_block.block_w0_reg[10] ),
    .Z(_07258_));
 INV_X1 _29724_ (.A(_07258_),
    .ZN(_07259_));
 BUF_X8 _29725_ (.A(_06698_),
    .Z(_07260_));
 BUF_X4 _29726_ (.A(\core.keymem.prev_key1_reg[8] ),
    .Z(_07261_));
 INV_X4 _29727_ (.A(_07261_),
    .ZN(_07262_));
 NOR2_X4 _29728_ (.A1(_07262_),
    .A2(_06837_),
    .ZN(_07263_));
 BUF_X4 _29729_ (.A(_06738_),
    .Z(_07264_));
 AOI21_X1 _29730_ (.A(_06866_),
    .B1(_07237_),
    .B2(_07264_),
    .ZN(_07265_));
 BUF_X4 _29731_ (.A(_06750_),
    .Z(_07266_));
 CLKBUF_X3 _29732_ (.A(\core.enc_block.block_w1_reg[8] ),
    .Z(_07267_));
 INV_X1 _29733_ (.A(_07267_),
    .ZN(_07268_));
 OAI221_X2 _29734_ (.A(_07265_),
    .B1(_07266_),
    .B2(_07268_),
    .C1(_00394_),
    .C2(_16252_),
    .ZN(_07269_));
 NAND2_X2 _29735_ (.A1(_06702_),
    .A2(_00393_),
    .ZN(_07270_));
 AND4_X4 _29736_ (.A1(_06843_),
    .A2(_06757_),
    .A3(_07269_),
    .A4(_07270_),
    .ZN(_07271_));
 BUF_X4 _29737_ (.A(_00398_),
    .Z(_07272_));
 NOR2_X4 _29738_ (.A1(_07272_),
    .A2(_06820_),
    .ZN(_07273_));
 BUF_X4 _29739_ (.A(\core.enc_block.block_w2_reg[10] ),
    .Z(_07274_));
 AOI21_X1 _29740_ (.A(_06713_),
    .B1(_07274_),
    .B2(_06716_),
    .ZN(_07275_));
 CLKBUF_X3 _29741_ (.A(\core.enc_block.block_w1_reg[10] ),
    .Z(_07276_));
 INV_X1 _29742_ (.A(_07276_),
    .ZN(_07277_));
 OAI221_X2 _29743_ (.A(_07275_),
    .B1(_06720_),
    .B2(_07277_),
    .C1(_00400_),
    .C2(_16251_),
    .ZN(_07278_));
 NAND2_X1 _29744_ (.A1(_06701_),
    .A2(_00399_),
    .ZN(_07279_));
 AND4_X1 _29745_ (.A1(_06696_),
    .A2(_06835_),
    .A3(_07278_),
    .A4(_07279_),
    .ZN(_07280_));
 BUF_X4 _29746_ (.A(_07280_),
    .Z(_07281_));
 OAI22_X4 _29747_ (.A1(_07263_),
    .A2(_07271_),
    .B1(_07273_),
    .B2(_07281_),
    .ZN(_07282_));
 CLKBUF_X3 _29748_ (.A(\core.enc_block.block_w2_reg[11] ),
    .Z(_07283_));
 AOI21_X1 _29749_ (.A(_06700_),
    .B1(_07283_),
    .B2(_06716_),
    .ZN(_07284_));
 BUF_X2 _29750_ (.A(\core.enc_block.block_w1_reg[11] ),
    .Z(_07285_));
 INV_X1 _29751_ (.A(_07285_),
    .ZN(_07286_));
 OAI221_X2 _29752_ (.A(_07284_),
    .B1(_07266_),
    .B2(_07286_),
    .C1(_00403_),
    .C2(_16251_),
    .ZN(_07287_));
 NAND2_X1 _29753_ (.A1(_06866_),
    .A2(_00402_),
    .ZN(_07288_));
 NAND4_X4 _29754_ (.A1(_06843_),
    .A2(_06779_),
    .A3(_07287_),
    .A4(_07288_),
    .ZN(_07289_));
 CLKBUF_X3 _29755_ (.A(_00395_),
    .Z(_07290_));
 NOR2_X4 _29756_ (.A1(_07290_),
    .A2(_06757_),
    .ZN(_07291_));
 CLKBUF_X3 _29757_ (.A(\core.enc_block.block_w2_reg[9] ),
    .Z(_07292_));
 AOI21_X1 _29758_ (.A(_06700_),
    .B1(_07292_),
    .B2(_07264_),
    .ZN(_07293_));
 BUF_X2 _29759_ (.A(\core.enc_block.block_w1_reg[9] ),
    .Z(_07294_));
 INV_X1 _29760_ (.A(_07294_),
    .ZN(_07295_));
 BUF_X2 _29761_ (.A(_00397_),
    .Z(_07296_));
 OAI221_X2 _29762_ (.A(_07293_),
    .B1(_07266_),
    .B2(_07295_),
    .C1(_07296_),
    .C2(_16251_),
    .ZN(_07297_));
 BUF_X2 _29763_ (.A(_00396_),
    .Z(_07298_));
 NAND2_X1 _29764_ (.A1(_06866_),
    .A2(_07298_),
    .ZN(_07299_));
 AND4_X1 _29765_ (.A1(_06760_),
    .A2(_06745_),
    .A3(_07297_),
    .A4(_07299_),
    .ZN(_07300_));
 BUF_X4 _29766_ (.A(_07300_),
    .Z(_07301_));
 CLKBUF_X3 _29767_ (.A(_00401_),
    .Z(_07302_));
 OAI221_X2 _29768_ (.A(_07289_),
    .B1(_07291_),
    .B2(_07301_),
    .C1(_06934_),
    .C2(_07302_),
    .ZN(_07303_));
 BUF_X4 _29769_ (.A(_07303_),
    .Z(_07304_));
 NOR2_X4 _29770_ (.A1(_07282_),
    .A2(_07304_),
    .ZN(_07305_));
 BUF_X2 _29771_ (.A(\core.enc_block.block_w2_reg[13] ),
    .Z(_07306_));
 AOI21_X1 _29772_ (.A(_06700_),
    .B1(_07306_),
    .B2(_06716_),
    .ZN(_07307_));
 BUF_X2 _29773_ (.A(\core.enc_block.block_w1_reg[13] ),
    .Z(_07308_));
 INV_X1 _29774_ (.A(_07308_),
    .ZN(_07309_));
 OAI221_X2 _29775_ (.A(_07307_),
    .B1(_07266_),
    .B2(_07309_),
    .C1(_00386_),
    .C2(_16251_),
    .ZN(_07310_));
 NAND2_X2 _29776_ (.A1(_06866_),
    .A2(_00385_),
    .ZN(_07311_));
 NAND4_X4 _29777_ (.A1(_06843_),
    .A2(_06779_),
    .A3(_07310_),
    .A4(_07311_),
    .ZN(_07312_));
 BUF_X4 _29778_ (.A(\core.keymem.prev_key1_reg[12] ),
    .Z(_07313_));
 INV_X1 _29779_ (.A(_07313_),
    .ZN(_07314_));
 BUF_X8 _29780_ (.A(_06745_),
    .Z(_07315_));
 NOR2_X4 _29781_ (.A1(_07314_),
    .A2(_07315_),
    .ZN(_07316_));
 BUF_X2 _29782_ (.A(\core.enc_block.block_w2_reg[12] ),
    .Z(_07317_));
 AOI21_X1 _29783_ (.A(_06700_),
    .B1(_07317_),
    .B2(_06716_),
    .ZN(_07318_));
 CLKBUF_X2 _29784_ (.A(\core.enc_block.block_w1_reg[12] ),
    .Z(_07319_));
 INV_X1 _29785_ (.A(_07319_),
    .ZN(_07320_));
 BUF_X2 _29786_ (.A(_00383_),
    .Z(_07321_));
 OAI221_X2 _29787_ (.A(_07318_),
    .B1(_06720_),
    .B2(_07320_),
    .C1(_07321_),
    .C2(_16251_),
    .ZN(_07322_));
 CLKBUF_X2 _29788_ (.A(_00382_),
    .Z(_07323_));
 NAND2_X1 _29789_ (.A1(_06866_),
    .A2(_07323_),
    .ZN(_07324_));
 AND4_X1 _29790_ (.A1(_06696_),
    .A2(_06835_),
    .A3(_07322_),
    .A4(_07324_),
    .ZN(_07325_));
 BUF_X4 _29791_ (.A(_07325_),
    .Z(_07326_));
 OAI221_X2 _29792_ (.A(_07312_),
    .B1(_07316_),
    .B2(_07326_),
    .C1(_06919_),
    .C2(_00384_),
    .ZN(_07327_));
 BUF_X4 _29793_ (.A(_07327_),
    .Z(_07328_));
 BUF_X4 _29794_ (.A(\core.enc_block.block_w2_reg[14] ),
    .Z(_07329_));
 AOI21_X1 _29795_ (.A(_06713_),
    .B1(_07329_),
    .B2(_06716_),
    .ZN(_07330_));
 BUF_X2 _29796_ (.A(\core.enc_block.block_w1_reg[14] ),
    .Z(_07331_));
 INV_X1 _29797_ (.A(_07331_),
    .ZN(_07332_));
 OAI221_X2 _29798_ (.A(_07330_),
    .B1(_06720_),
    .B2(_07332_),
    .C1(_00389_),
    .C2(_16251_),
    .ZN(_07333_));
 NAND2_X1 _29799_ (.A1(_06701_),
    .A2(_00388_),
    .ZN(_07334_));
 AND4_X1 _29800_ (.A1(_06696_),
    .A2(_06835_),
    .A3(_07333_),
    .A4(_07334_),
    .ZN(_07335_));
 BUF_X4 _29801_ (.A(_07335_),
    .Z(_07336_));
 NOR2_X4 _29802_ (.A1(_00387_),
    .A2(_06779_),
    .ZN(_07337_));
 BUF_X4 _29803_ (.A(\core.enc_block.block_w2_reg[15] ),
    .Z(_07338_));
 AOI21_X1 _29804_ (.A(_06725_),
    .B1(_07338_),
    .B2(_07264_),
    .ZN(_07339_));
 BUF_X4 _29805_ (.A(\core.enc_block.block_w1_reg[15] ),
    .Z(_07340_));
 INV_X1 _29806_ (.A(_07340_),
    .ZN(_07341_));
 OAI221_X2 _29807_ (.A(_07339_),
    .B1(_07266_),
    .B2(_07341_),
    .C1(_00392_),
    .C2(_16252_),
    .ZN(_07342_));
 NAND2_X2 _29808_ (.A1(_06702_),
    .A2(_00391_),
    .ZN(_07343_));
 AND4_X4 _29809_ (.A1(_06733_),
    .A2(_06711_),
    .A3(_07342_),
    .A4(_07343_),
    .ZN(_07344_));
 NOR2_X4 _29810_ (.A1(_00390_),
    .A2(_06820_),
    .ZN(_07345_));
 OAI22_X4 _29811_ (.A1(_07336_),
    .A2(_07337_),
    .B1(_07344_),
    .B2(_07345_),
    .ZN(_07346_));
 NOR2_X4 _29812_ (.A1(_07328_),
    .A2(_07346_),
    .ZN(_07347_));
 NAND4_X4 _29813_ (.A1(_06843_),
    .A2(_07315_),
    .A3(_07333_),
    .A4(_07334_),
    .ZN(_07348_));
 BUF_X4 _29814_ (.A(\core.keymem.prev_key1_reg[14] ),
    .Z(_07349_));
 NAND2_X4 _29815_ (.A1(_07349_),
    .A2(_06938_),
    .ZN(_07350_));
 NOR2_X4 _29816_ (.A1(_00384_),
    .A2(_06735_),
    .ZN(_07351_));
 AND4_X4 _29817_ (.A1(_06760_),
    .A2(_06735_),
    .A3(_07310_),
    .A4(_07311_),
    .ZN(_07352_));
 OAI211_X4 _29818_ (.A(_07348_),
    .B(_07350_),
    .C1(_07351_),
    .C2(_07352_),
    .ZN(_07353_));
 NAND2_X4 _29819_ (.A1(_07313_),
    .A2(_06841_),
    .ZN(_07354_));
 NAND4_X4 _29820_ (.A1(_06697_),
    .A2(_07315_),
    .A3(_07322_),
    .A4(_07324_),
    .ZN(_07355_));
 NAND4_X4 _29821_ (.A1(_06697_),
    .A2(_07315_),
    .A3(_07342_),
    .A4(_07343_),
    .ZN(_07356_));
 BUF_X4 _29822_ (.A(\core.keymem.prev_key1_reg[15] ),
    .Z(_07357_));
 NAND2_X2 _29823_ (.A1(_07357_),
    .A2(_06841_),
    .ZN(_07358_));
 NAND4_X4 _29824_ (.A1(_07354_),
    .A2(_07355_),
    .A3(_07356_),
    .A4(_07358_),
    .ZN(_07359_));
 BUF_X4 _29825_ (.A(_07359_),
    .Z(_07360_));
 NOR2_X1 _29826_ (.A1(_07353_),
    .A2(_07360_),
    .ZN(_07361_));
 CLKBUF_X3 _29827_ (.A(_07361_),
    .Z(_07362_));
 OAI21_X1 _29828_ (.A(_07305_),
    .B1(_07347_),
    .B2(_07362_),
    .ZN(_07363_));
 INV_X1 _29829_ (.A(_07357_),
    .ZN(_07364_));
 OAI221_X2 _29830_ (.A(_07356_),
    .B1(_07337_),
    .B2(_07336_),
    .C1(_07364_),
    .C2(_06822_),
    .ZN(_07365_));
 BUF_X8 _29831_ (.A(_07365_),
    .Z(_07366_));
 OAI22_X4 _29832_ (.A1(_07351_),
    .A2(_07352_),
    .B1(_07316_),
    .B2(_07326_),
    .ZN(_07367_));
 NOR2_X4 _29833_ (.A1(_07366_),
    .A2(_07367_),
    .ZN(_07368_));
 BUF_X4 _29834_ (.A(_07368_),
    .Z(_07369_));
 INV_X4 _29835_ (.A(_07290_),
    .ZN(_07370_));
 NAND2_X4 _29836_ (.A1(_07370_),
    .A2(_06841_),
    .ZN(_07371_));
 NAND4_X4 _29837_ (.A1(_06697_),
    .A2(_07315_),
    .A3(_07297_),
    .A4(_07299_),
    .ZN(_07372_));
 NAND2_X4 _29838_ (.A1(_07371_),
    .A2(_07372_),
    .ZN(_07373_));
 BUF_X4 _29839_ (.A(_07373_),
    .Z(_07374_));
 NOR2_X4 _29840_ (.A1(_07302_),
    .A2(_06779_),
    .ZN(_07375_));
 AND4_X1 _29841_ (.A1(_06760_),
    .A2(_06745_),
    .A3(_07287_),
    .A4(_07288_),
    .ZN(_07376_));
 BUF_X8 _29842_ (.A(_07376_),
    .Z(_07377_));
 OAI22_X4 _29843_ (.A1(_07375_),
    .A2(_07377_),
    .B1(_07273_),
    .B2(_07281_),
    .ZN(_07378_));
 NOR2_X4 _29844_ (.A1(_07374_),
    .A2(_07378_),
    .ZN(_07379_));
 NOR2_X4 _29845_ (.A1(_07291_),
    .A2(_07301_),
    .ZN(_07380_));
 BUF_X4 _29846_ (.A(_07380_),
    .Z(_07381_));
 INV_X4 _29847_ (.A(_07302_),
    .ZN(_07382_));
 NAND2_X4 _29848_ (.A1(_07382_),
    .A2(_06938_),
    .ZN(_07383_));
 INV_X1 _29849_ (.A(_07272_),
    .ZN(_07384_));
 NAND2_X4 _29850_ (.A1(_07384_),
    .A2(_06841_),
    .ZN(_07385_));
 NAND4_X4 _29851_ (.A1(_06843_),
    .A2(_06757_),
    .A3(_07278_),
    .A4(_07279_),
    .ZN(_07386_));
 NAND4_X4 _29852_ (.A1(_07383_),
    .A2(_07289_),
    .A3(_07385_),
    .A4(_07386_),
    .ZN(_07387_));
 BUF_X4 _29853_ (.A(_07387_),
    .Z(_07388_));
 NOR2_X1 _29854_ (.A1(_07381_),
    .A2(_07388_),
    .ZN(_07389_));
 BUF_X4 _29855_ (.A(_07389_),
    .Z(_07390_));
 NOR2_X4 _29856_ (.A1(_07316_),
    .A2(_07326_),
    .ZN(_07391_));
 BUF_X4 _29857_ (.A(_07366_),
    .Z(_07392_));
 BUF_X4 _29858_ (.A(_07392_),
    .Z(_07393_));
 NOR2_X1 _29859_ (.A1(_07391_),
    .A2(_07393_),
    .ZN(_07394_));
 AOI22_X2 _29860_ (.A1(_07369_),
    .A2(_07379_),
    .B1(_07390_),
    .B2(_07394_),
    .ZN(_07395_));
 NOR2_X4 _29861_ (.A1(_07263_),
    .A2(_07271_),
    .ZN(_07396_));
 BUF_X4 _29862_ (.A(_07396_),
    .Z(_07397_));
 BUF_X4 _29863_ (.A(_07397_),
    .Z(_07398_));
 BUF_X4 _29864_ (.A(_07398_),
    .Z(_07399_));
 BUF_X4 _29865_ (.A(_07399_),
    .Z(_07400_));
 OAI21_X2 _29866_ (.A(_07363_),
    .B1(_07395_),
    .B2(_07400_),
    .ZN(_07401_));
 BUF_X4 _29867_ (.A(_07346_),
    .Z(_07402_));
 BUF_X4 _29868_ (.A(_07367_),
    .Z(_07403_));
 NOR2_X4 _29869_ (.A1(_07402_),
    .A2(_07403_),
    .ZN(_07404_));
 NAND2_X4 _29870_ (.A1(_07261_),
    .A2(_06841_),
    .ZN(_07405_));
 NAND4_X4 _29871_ (.A1(_06843_),
    .A2(_06757_),
    .A3(_07269_),
    .A4(_07270_),
    .ZN(_07406_));
 NAND2_X4 _29872_ (.A1(_07405_),
    .A2(_07406_),
    .ZN(_07407_));
 BUF_X4 _29873_ (.A(_07407_),
    .Z(_07408_));
 NAND2_X4 _29874_ (.A1(_07385_),
    .A2(_07386_),
    .ZN(_07409_));
 BUF_X4 _29875_ (.A(_07409_),
    .Z(_07410_));
 BUF_X4 _29876_ (.A(_07410_),
    .Z(_07411_));
 NOR2_X2 _29877_ (.A1(_07408_),
    .A2(_07411_),
    .ZN(_07412_));
 NAND2_X1 _29878_ (.A1(_07404_),
    .A2(_07412_),
    .ZN(_07413_));
 NOR2_X4 _29879_ (.A1(_07273_),
    .A2(_07281_),
    .ZN(_07414_));
 BUF_X4 _29880_ (.A(_07414_),
    .Z(_07415_));
 BUF_X4 _29881_ (.A(_07415_),
    .Z(_07416_));
 BUF_X4 _29882_ (.A(_07416_),
    .Z(_07417_));
 CLKBUF_X3 _29883_ (.A(_07393_),
    .Z(_07418_));
 BUF_X8 _29884_ (.A(_07315_),
    .Z(_07419_));
 OAI221_X2 _29885_ (.A(_07355_),
    .B1(_07352_),
    .B2(_07351_),
    .C1(_07314_),
    .C2(_07419_),
    .ZN(_07420_));
 BUF_X4 _29886_ (.A(_07420_),
    .Z(_07421_));
 BUF_X4 _29887_ (.A(_07421_),
    .Z(_07422_));
 NOR3_X2 _29888_ (.A1(_07417_),
    .A2(_07418_),
    .A3(_07422_),
    .ZN(_07423_));
 OR2_X4 _29889_ (.A1(_00384_),
    .A2(_06837_),
    .ZN(_07424_));
 NAND4_X4 _29890_ (.A1(_07424_),
    .A2(_07312_),
    .A3(_07348_),
    .A4(_07350_),
    .ZN(_07425_));
 NOR2_X4 _29891_ (.A1(_07425_),
    .A2(_07360_),
    .ZN(_07426_));
 BUF_X4 _29892_ (.A(_07416_),
    .Z(_07427_));
 BUF_X4 _29893_ (.A(_07427_),
    .Z(_07428_));
 AOI21_X1 _29894_ (.A(_07423_),
    .B1(_07426_),
    .B2(_07428_),
    .ZN(_07429_));
 OAI21_X2 _29895_ (.A(_07413_),
    .B1(_07429_),
    .B2(_07400_),
    .ZN(_07430_));
 NAND2_X4 _29896_ (.A1(_07383_),
    .A2(_07289_),
    .ZN(_07431_));
 BUF_X4 _29897_ (.A(_07431_),
    .Z(_07432_));
 NOR2_X4 _29898_ (.A1(_07432_),
    .A2(_07374_),
    .ZN(_07433_));
 AOI21_X4 _29899_ (.A(_07401_),
    .B1(_07430_),
    .B2(_07433_),
    .ZN(_07434_));
 NOR2_X4 _29900_ (.A1(_07375_),
    .A2(_07377_),
    .ZN(_07435_));
 BUF_X4 _29901_ (.A(_07435_),
    .Z(_07436_));
 BUF_X4 _29902_ (.A(_07436_),
    .Z(_07437_));
 BUF_X4 _29903_ (.A(_07437_),
    .Z(_07438_));
 BUF_X4 _29904_ (.A(_07438_),
    .Z(_07439_));
 AOI22_X4 _29905_ (.A1(_07405_),
    .A2(_07406_),
    .B1(_07385_),
    .B2(_07386_),
    .ZN(_07440_));
 BUF_X4 _29906_ (.A(_07328_),
    .Z(_07441_));
 NOR2_X1 _29907_ (.A1(_07441_),
    .A2(_07392_),
    .ZN(_07442_));
 BUF_X4 _29908_ (.A(_07442_),
    .Z(_07443_));
 NOR2_X4 _29909_ (.A1(_07407_),
    .A2(_07373_),
    .ZN(_07444_));
 NOR3_X4 _29910_ (.A1(_07409_),
    .A2(_07366_),
    .A3(_07420_),
    .ZN(_07445_));
 AOI22_X2 _29911_ (.A1(_07440_),
    .A2(_07443_),
    .B1(_07444_),
    .B2(_07445_),
    .ZN(_07446_));
 BUF_X4 _29912_ (.A(_07411_),
    .Z(_07447_));
 BUF_X4 _29913_ (.A(_07432_),
    .Z(_07448_));
 BUF_X4 _29914_ (.A(_07448_),
    .Z(_07449_));
 BUF_X4 _29915_ (.A(_07381_),
    .Z(_07450_));
 BUF_X4 _29916_ (.A(_07402_),
    .Z(_07451_));
 CLKBUF_X3 _29917_ (.A(_07451_),
    .Z(_07452_));
 NAND4_X4 _29918_ (.A1(_07424_),
    .A2(_07312_),
    .A3(_07354_),
    .A4(_07355_),
    .ZN(_07453_));
 BUF_X4 _29919_ (.A(_07453_),
    .Z(_07454_));
 CLKBUF_X3 _29920_ (.A(_07454_),
    .Z(_07455_));
 NOR4_X1 _29921_ (.A1(_07449_),
    .A2(_07450_),
    .A3(_07452_),
    .A4(_07455_),
    .ZN(_07456_));
 BUF_X4 _29922_ (.A(_07374_),
    .Z(_07457_));
 BUF_X4 _29923_ (.A(_07403_),
    .Z(_07458_));
 CLKBUF_X3 _29924_ (.A(_07458_),
    .Z(_07459_));
 NOR4_X1 _29925_ (.A1(_07438_),
    .A2(_07418_),
    .A3(_07457_),
    .A4(_07459_),
    .ZN(_07460_));
 NOR3_X1 _29926_ (.A1(_07447_),
    .A2(_07456_),
    .A3(_07460_),
    .ZN(_07461_));
 AOI221_X2 _29927_ (.A(_07301_),
    .B1(_07289_),
    .B2(_07383_),
    .C1(_07370_),
    .C2(_07109_),
    .ZN(_07462_));
 CLKBUF_X3 _29928_ (.A(_07462_),
    .Z(_07463_));
 NOR3_X2 _29929_ (.A1(_07397_),
    .A2(_07392_),
    .A3(_07422_),
    .ZN(_07464_));
 OAI22_X4 _29930_ (.A1(_07263_),
    .A2(_07271_),
    .B1(_07291_),
    .B2(_07301_),
    .ZN(_07465_));
 INV_X2 _29931_ (.A(_07349_),
    .ZN(_07466_));
 OAI221_X2 _29932_ (.A(_07348_),
    .B1(_07344_),
    .B2(_07345_),
    .C1(_06822_),
    .C2(_07466_),
    .ZN(_07467_));
 BUF_X4 _29933_ (.A(_07467_),
    .Z(_07468_));
 NOR3_X4 _29934_ (.A1(_07431_),
    .A2(_07403_),
    .A3(_07468_),
    .ZN(_07469_));
 AOI221_X2 _29935_ (.A(_07427_),
    .B1(_07463_),
    .B2(_07464_),
    .C1(_07465_),
    .C2(_07469_),
    .ZN(_07470_));
 OAI22_X2 _29936_ (.A1(_07439_),
    .A2(_07446_),
    .B1(_07461_),
    .B2(_07470_),
    .ZN(_07471_));
 NOR2_X4 _29937_ (.A1(_07366_),
    .A2(_07421_),
    .ZN(_07472_));
 AOI221_X2 _29938_ (.A(_07271_),
    .B1(_07371_),
    .B2(_07372_),
    .C1(_06936_),
    .C2(_07261_),
    .ZN(_07473_));
 BUF_X4 _29939_ (.A(_07473_),
    .Z(_07474_));
 BUF_X4 _29940_ (.A(_07468_),
    .Z(_07475_));
 BUF_X4 _29941_ (.A(_07475_),
    .Z(_07476_));
 OAI221_X2 _29942_ (.A(_07386_),
    .B1(_07377_),
    .B2(_07375_),
    .C1(_07272_),
    .C2(_06887_),
    .ZN(_07477_));
 OAI33_X1 _29943_ (.A1(_07436_),
    .A2(_07422_),
    .A3(_07476_),
    .B1(_07477_),
    .B2(_07392_),
    .B3(_07441_),
    .ZN(_07478_));
 OAI221_X2 _29944_ (.A(_07356_),
    .B1(_07326_),
    .B2(_07316_),
    .C1(_07364_),
    .C2(_06886_),
    .ZN(_07479_));
 BUF_X4 _29945_ (.A(_07479_),
    .Z(_07480_));
 NOR2_X2 _29946_ (.A1(_07425_),
    .A2(_07480_),
    .ZN(_07481_));
 BUF_X4 _29947_ (.A(_07481_),
    .Z(_07482_));
 AOI222_X2 _29948_ (.A1(_07472_),
    .A2(_07305_),
    .B1(_07474_),
    .B2(_07478_),
    .C1(_07482_),
    .C2(_07379_),
    .ZN(_07483_));
 BUF_X4 _29949_ (.A(_07441_),
    .Z(_07484_));
 BUF_X8 _29950_ (.A(_07372_),
    .Z(_07485_));
 BUF_X4 _29951_ (.A(_06919_),
    .Z(_07486_));
 OAI221_X2 _29952_ (.A(_07485_),
    .B1(_07281_),
    .B2(_07273_),
    .C1(_07290_),
    .C2(_07486_),
    .ZN(_07487_));
 OAI221_X2 _29953_ (.A(_07386_),
    .B1(_07291_),
    .B2(_07301_),
    .C1(_06887_),
    .C2(_07272_),
    .ZN(_07488_));
 CLKBUF_X3 _29954_ (.A(_07422_),
    .Z(_07489_));
 OAI22_X1 _29955_ (.A1(_07484_),
    .A2(_07487_),
    .B1(_07488_),
    .B2(_07489_),
    .ZN(_07490_));
 BUF_X4 _29956_ (.A(_07408_),
    .Z(_07491_));
 NOR3_X1 _29957_ (.A1(_07438_),
    .A2(_07491_),
    .A3(_07452_),
    .ZN(_07492_));
 NOR2_X4 _29958_ (.A1(_07328_),
    .A2(_07468_),
    .ZN(_07493_));
 BUF_X4 _29959_ (.A(_07493_),
    .Z(_07494_));
 NOR3_X4 _29960_ (.A1(_07435_),
    .A2(_07409_),
    .A3(_07373_),
    .ZN(_07495_));
 NAND4_X4 _29961_ (.A1(_07383_),
    .A2(_07289_),
    .A3(_07371_),
    .A4(_07485_),
    .ZN(_07496_));
 BUF_X4 _29962_ (.A(_07496_),
    .Z(_07497_));
 OAI221_X1 _29963_ (.A(_07386_),
    .B1(_07271_),
    .B2(_07263_),
    .C1(_07272_),
    .C2(_07486_),
    .ZN(_07498_));
 CLKBUF_X3 _29964_ (.A(_07498_),
    .Z(_07499_));
 NOR2_X2 _29965_ (.A1(_07497_),
    .A2(_07499_),
    .ZN(_07500_));
 AOI222_X2 _29966_ (.A1(_07490_),
    .A2(_07492_),
    .B1(_07494_),
    .B2(_07495_),
    .C1(_07500_),
    .C2(_07347_),
    .ZN(_07501_));
 NAND2_X1 _29967_ (.A1(_07483_),
    .A2(_07501_),
    .ZN(_07502_));
 OAI221_X2 _29968_ (.A(_07406_),
    .B1(_07273_),
    .B2(_07281_),
    .C1(_06919_),
    .C2(_07262_),
    .ZN(_07503_));
 BUF_X4 _29969_ (.A(_07503_),
    .Z(_07504_));
 OAI22_X4 _29970_ (.A1(_07375_),
    .A2(_07377_),
    .B1(_07291_),
    .B2(_07301_),
    .ZN(_07505_));
 NOR4_X4 _29971_ (.A1(_07366_),
    .A2(_07420_),
    .A3(_07504_),
    .A4(_07505_),
    .ZN(_07506_));
 NOR2_X4 _29972_ (.A1(_07421_),
    .A2(_07475_),
    .ZN(_07507_));
 AOI21_X1 _29973_ (.A(_07506_),
    .B1(_07507_),
    .B2(_07305_),
    .ZN(_07508_));
 BUF_X4 _29974_ (.A(_07346_),
    .Z(_07509_));
 NOR3_X2 _29975_ (.A1(_07436_),
    .A2(_07509_),
    .A3(_07454_),
    .ZN(_07510_));
 AOI221_X2 _29976_ (.A(_07301_),
    .B1(_07406_),
    .B2(_07405_),
    .C1(_07370_),
    .C2(_06936_),
    .ZN(_07511_));
 BUF_X4 _29977_ (.A(_07511_),
    .Z(_07512_));
 AOI221_X2 _29978_ (.A(_07281_),
    .B1(_07371_),
    .B2(_07485_),
    .C1(_06936_),
    .C2(_07384_),
    .ZN(_07513_));
 OAI21_X1 _29979_ (.A(_07510_),
    .B1(_07512_),
    .B2(_07513_),
    .ZN(_07514_));
 AOI22_X4 _29980_ (.A1(_07405_),
    .A2(_07406_),
    .B1(_07371_),
    .B2(_07485_),
    .ZN(_07515_));
 OAI221_X2 _29981_ (.A(_07289_),
    .B1(_07273_),
    .B2(_07281_),
    .C1(_06934_),
    .C2(_07302_),
    .ZN(_07516_));
 BUF_X4 _29982_ (.A(_07516_),
    .Z(_07517_));
 NOR2_X1 _29983_ (.A1(_07515_),
    .A2(_07517_),
    .ZN(_07518_));
 NOR3_X1 _29984_ (.A1(_07398_),
    .A2(_07484_),
    .A3(_07393_),
    .ZN(_07519_));
 OAI21_X1 _29985_ (.A(_07518_),
    .B1(_07519_),
    .B2(_07362_),
    .ZN(_07520_));
 NAND3_X2 _29986_ (.A1(_07508_),
    .A2(_07514_),
    .A3(_07520_),
    .ZN(_07521_));
 BUF_X4 _29987_ (.A(_07457_),
    .Z(_07522_));
 NAND2_X4 _29988_ (.A1(_07356_),
    .A2(_07358_),
    .ZN(_07523_));
 BUF_X4 _29989_ (.A(_07523_),
    .Z(_07524_));
 NAND2_X2 _29990_ (.A1(_07348_),
    .A2(_07350_),
    .ZN(_07525_));
 BUF_X4 _29991_ (.A(_07525_),
    .Z(_07526_));
 NOR2_X1 _29992_ (.A1(_07524_),
    .A2(_07526_),
    .ZN(_07527_));
 NAND2_X1 _29993_ (.A1(_07522_),
    .A2(_07527_),
    .ZN(_07528_));
 NOR2_X2 _29994_ (.A1(_07351_),
    .A2(_07352_),
    .ZN(_07529_));
 CLKBUF_X3 _29995_ (.A(_07529_),
    .Z(_07530_));
 NAND2_X4 _29996_ (.A1(_07354_),
    .A2(_07355_),
    .ZN(_07531_));
 CLKBUF_X3 _29997_ (.A(_07531_),
    .Z(_07532_));
 NOR2_X1 _29998_ (.A1(_07437_),
    .A2(_07499_),
    .ZN(_07533_));
 NAND3_X1 _29999_ (.A1(_07530_),
    .A2(_07532_),
    .A3(_07533_),
    .ZN(_07534_));
 NAND2_X4 _30000_ (.A1(_07424_),
    .A2(_07312_),
    .ZN(_07535_));
 BUF_X4 _30001_ (.A(_07535_),
    .Z(_07536_));
 OAI221_X2 _30002_ (.A(_07289_),
    .B1(_07316_),
    .B2(_07326_),
    .C1(_06888_),
    .C2(_07302_),
    .ZN(_07537_));
 NOR3_X1 _30003_ (.A1(_07427_),
    .A2(_07536_),
    .A3(_07537_),
    .ZN(_07538_));
 NOR3_X1 _30004_ (.A1(_07438_),
    .A2(_07447_),
    .A3(_07489_),
    .ZN(_07539_));
 OAI21_X1 _30005_ (.A(_07400_),
    .B1(_07538_),
    .B2(_07539_),
    .ZN(_07540_));
 AOI21_X2 _30006_ (.A(_07528_),
    .B1(_07534_),
    .B2(_07540_),
    .ZN(_07541_));
 NOR4_X2 _30007_ (.A1(_07471_),
    .A2(_07502_),
    .A3(_07521_),
    .A4(_07541_),
    .ZN(_07542_));
 BUF_X4 _30008_ (.A(_07450_),
    .Z(_07543_));
 NOR2_X4 _30009_ (.A1(_07353_),
    .A2(_07480_),
    .ZN(_07544_));
 CLKBUF_X3 _30010_ (.A(_07544_),
    .Z(_07545_));
 NAND2_X1 _30011_ (.A1(_07428_),
    .A2(_07545_),
    .ZN(_07546_));
 BUF_X4 _30012_ (.A(_07408_),
    .Z(_07547_));
 OAI21_X1 _30013_ (.A(_07547_),
    .B1(_07445_),
    .B2(_07545_),
    .ZN(_07548_));
 AOI21_X1 _30014_ (.A(_07449_),
    .B1(_07546_),
    .B2(_07548_),
    .ZN(_07549_));
 BUF_X4 _30015_ (.A(_07477_),
    .Z(_07550_));
 NOR2_X4 _30016_ (.A1(_07367_),
    .A2(_07468_),
    .ZN(_07551_));
 BUF_X4 _30017_ (.A(_07551_),
    .Z(_07552_));
 NAND2_X1 _30018_ (.A1(_07484_),
    .A2(_07489_),
    .ZN(_07553_));
 AOI21_X1 _30019_ (.A(_07552_),
    .B1(_07527_),
    .B2(_07553_),
    .ZN(_07554_));
 NOR2_X1 _30020_ (.A1(_07550_),
    .A2(_07554_),
    .ZN(_07555_));
 OAI21_X2 _30021_ (.A(_07543_),
    .B1(_07549_),
    .B2(_07555_),
    .ZN(_07556_));
 AOI22_X4 _30022_ (.A1(_07385_),
    .A2(_07386_),
    .B1(_07371_),
    .B2(_07485_),
    .ZN(_07557_));
 NOR3_X1 _30023_ (.A1(_07454_),
    .A2(_07475_),
    .A3(_07557_),
    .ZN(_07558_));
 AOI221_X2 _30024_ (.A(_07377_),
    .B1(_07371_),
    .B2(_07485_),
    .C1(_07108_),
    .C2(_07382_),
    .ZN(_07559_));
 AOI211_X2 _30025_ (.A(_07453_),
    .B(_07468_),
    .C1(_07559_),
    .C2(_07396_),
    .ZN(_07560_));
 NOR2_X4 _30026_ (.A1(_07402_),
    .A2(_07454_),
    .ZN(_07561_));
 NOR2_X4 _30027_ (.A1(_07453_),
    .A2(_07468_),
    .ZN(_07562_));
 OAI222_X2 _30028_ (.A1(_07437_),
    .A2(_07558_),
    .B1(_07560_),
    .B2(_07410_),
    .C1(_07561_),
    .C2(_07562_),
    .ZN(_07563_));
 NOR2_X2 _30029_ (.A1(_07381_),
    .A2(_07378_),
    .ZN(_07564_));
 OR2_X2 _30030_ (.A1(_00387_),
    .A2(_06934_),
    .ZN(_07565_));
 OAI22_X4 _30031_ (.A1(_07316_),
    .A2(_07326_),
    .B1(_07344_),
    .B2(_07345_),
    .ZN(_07566_));
 AOI221_X2 _30032_ (.A(_07535_),
    .B1(_07348_),
    .B2(_07565_),
    .C1(_07566_),
    .C2(_07360_),
    .ZN(_07567_));
 NAND2_X1 _30033_ (.A1(_07564_),
    .A2(_07567_),
    .ZN(_07568_));
 NOR2_X4 _30034_ (.A1(_07432_),
    .A2(_07415_),
    .ZN(_07569_));
 NOR2_X1 _30035_ (.A1(_07530_),
    .A2(_07509_),
    .ZN(_07570_));
 BUF_X4 _30036_ (.A(_07374_),
    .Z(_07571_));
 XNOR2_X1 _30037_ (.A(_07391_),
    .B(_07571_),
    .ZN(_07572_));
 NAND3_X2 _30038_ (.A1(_07569_),
    .A2(_07570_),
    .A3(_07572_),
    .ZN(_07573_));
 NAND3_X2 _30039_ (.A1(_07563_),
    .A2(_07568_),
    .A3(_07573_),
    .ZN(_07574_));
 NOR3_X1 _30040_ (.A1(_07532_),
    .A2(_07378_),
    .A3(_07474_),
    .ZN(_07575_));
 NOR3_X1 _30041_ (.A1(_07536_),
    .A2(_07524_),
    .A3(_07526_),
    .ZN(_07576_));
 OAI21_X2 _30042_ (.A(_07575_),
    .B1(_07576_),
    .B2(_07570_),
    .ZN(_07577_));
 BUF_X4 _30043_ (.A(_07360_),
    .Z(_07578_));
 NOR3_X2 _30044_ (.A1(_07336_),
    .A2(_07337_),
    .A3(_07350_),
    .ZN(_07579_));
 OAI22_X4 _30045_ (.A1(_07391_),
    .A2(_07451_),
    .B1(_07578_),
    .B2(_07579_),
    .ZN(_07580_));
 OAI221_X2 _30046_ (.A(_07406_),
    .B1(_07291_),
    .B2(_07301_),
    .C1(_06886_),
    .C2(_07262_),
    .ZN(_07581_));
 BUF_X4 _30047_ (.A(_07581_),
    .Z(_07582_));
 NOR3_X2 _30048_ (.A1(_07535_),
    .A2(_07582_),
    .A3(_07477_),
    .ZN(_07583_));
 AOI22_X4 _30049_ (.A1(_07390_),
    .A2(_07494_),
    .B1(_07580_),
    .B2(_07583_),
    .ZN(_07584_));
 CLKBUF_X3 _30050_ (.A(_07476_),
    .Z(_07585_));
 CLKBUF_X3 _30051_ (.A(_07425_),
    .Z(_07586_));
 OAI33_X1 _30052_ (.A1(_07439_),
    .A2(_07459_),
    .A3(_07585_),
    .B1(_07586_),
    .B2(_07578_),
    .B3(_07388_),
    .ZN(_07587_));
 NAND2_X1 _30053_ (.A1(_07474_),
    .A2(_07587_),
    .ZN(_07588_));
 NAND3_X2 _30054_ (.A1(_07577_),
    .A2(_07584_),
    .A3(_07588_),
    .ZN(_07589_));
 NOR4_X4 _30055_ (.A1(_07447_),
    .A2(_07524_),
    .A3(_07526_),
    .A4(_07474_),
    .ZN(_07590_));
 OAI21_X2 _30056_ (.A(_07489_),
    .B1(_07450_),
    .B2(_07484_),
    .ZN(_07591_));
 NOR2_X2 _30057_ (.A1(_07417_),
    .A2(_07582_),
    .ZN(_07592_));
 AOI22_X4 _30058_ (.A1(_07590_),
    .A2(_07591_),
    .B1(_07592_),
    .B2(_07507_),
    .ZN(_07593_));
 NOR2_X4 _30059_ (.A1(_07366_),
    .A2(_07453_),
    .ZN(_07594_));
 BUF_X4 _30060_ (.A(_07282_),
    .Z(_07595_));
 NOR2_X2 _30061_ (.A1(_07595_),
    .A2(_07457_),
    .ZN(_07596_));
 NOR2_X1 _30062_ (.A1(_07447_),
    .A2(_07582_),
    .ZN(_07597_));
 OAI21_X2 _30063_ (.A(_07594_),
    .B1(_07596_),
    .B2(_07597_),
    .ZN(_07598_));
 AOI21_X4 _30064_ (.A(_07449_),
    .B1(_07593_),
    .B2(_07598_),
    .ZN(_07599_));
 NOR3_X1 _30065_ (.A1(_07489_),
    .A2(_07585_),
    .A3(_07487_),
    .ZN(_07600_));
 NOR4_X1 _30066_ (.A1(_07418_),
    .A2(_07450_),
    .A3(_07489_),
    .A4(_07550_),
    .ZN(_07601_));
 OAI21_X1 _30067_ (.A(_07547_),
    .B1(_07600_),
    .B2(_07601_),
    .ZN(_07602_));
 NOR3_X4 _30068_ (.A1(_07436_),
    .A2(_07509_),
    .A3(_07458_),
    .ZN(_07603_));
 NOR3_X4 _30069_ (.A1(_07448_),
    .A2(_07484_),
    .A3(_07451_),
    .ZN(_07604_));
 OAI21_X1 _30070_ (.A(_07513_),
    .B1(_07603_),
    .B2(_07604_),
    .ZN(_07605_));
 NAND2_X1 _30071_ (.A1(_07379_),
    .A2(_07494_),
    .ZN(_07606_));
 NOR2_X4 _30072_ (.A1(_07304_),
    .A2(_07504_),
    .ZN(_07607_));
 NOR3_X1 _30073_ (.A1(_07530_),
    .A2(_07524_),
    .A3(_07526_),
    .ZN(_07608_));
 NOR2_X1 _30074_ (.A1(_07535_),
    .A2(_07451_),
    .ZN(_07609_));
 OAI221_X2 _30075_ (.A(_07607_),
    .B1(_07608_),
    .B2(_07609_),
    .C1(_07316_),
    .C2(_07326_),
    .ZN(_07610_));
 NAND4_X2 _30076_ (.A1(_07602_),
    .A2(_07605_),
    .A3(_07606_),
    .A4(_07610_),
    .ZN(_07611_));
 NOR4_X4 _30077_ (.A1(_07574_),
    .A2(_07589_),
    .A3(_07599_),
    .A4(_07611_),
    .ZN(_07612_));
 NAND4_X4 _30078_ (.A1(_07434_),
    .A2(_07542_),
    .A3(_07556_),
    .A4(_07612_),
    .ZN(_07613_));
 AOI221_X2 _30079_ (.A(_07326_),
    .B1(_07312_),
    .B2(_07424_),
    .C1(_07313_),
    .C2(_07109_),
    .ZN(_07614_));
 OR2_X2 _30080_ (.A1(_00390_),
    .A2(_06934_),
    .ZN(_07615_));
 AOI22_X4 _30081_ (.A1(_07348_),
    .A2(_07565_),
    .B1(_07356_),
    .B2(_07615_),
    .ZN(_07616_));
 NAND3_X1 _30082_ (.A1(_07543_),
    .A2(_07614_),
    .A3(_07616_),
    .ZN(_07617_));
 AOI21_X1 _30083_ (.A(_07439_),
    .B1(_07428_),
    .B2(_07617_),
    .ZN(_07618_));
 OAI22_X4 _30084_ (.A1(_07375_),
    .A2(_07377_),
    .B1(_07316_),
    .B2(_07326_),
    .ZN(_07619_));
 NOR2_X2 _30085_ (.A1(_07344_),
    .A2(_07345_),
    .ZN(_07620_));
 BUF_X4 _30086_ (.A(_07620_),
    .Z(_07621_));
 OAI33_X1 _30087_ (.A1(_07449_),
    .A2(_07452_),
    .A3(_07459_),
    .B1(_07586_),
    .B2(_07619_),
    .B3(_07621_),
    .ZN(_07622_));
 NOR3_X4 _30088_ (.A1(_07436_),
    .A2(_07441_),
    .A3(_07402_),
    .ZN(_07623_));
 MUX2_X1 _30089_ (.A(_07622_),
    .B(_07623_),
    .S(_07543_),
    .Z(_07624_));
 OAI21_X1 _30090_ (.A(_07428_),
    .B1(_07618_),
    .B2(_07624_),
    .ZN(_07625_));
 OAI21_X1 _30091_ (.A(_07618_),
    .B1(_07545_),
    .B2(_07404_),
    .ZN(_07626_));
 AOI21_X2 _30092_ (.A(_07400_),
    .B1(_07625_),
    .B2(_07626_),
    .ZN(_07627_));
 NOR3_X4 _30093_ (.A1(_07416_),
    .A2(_07535_),
    .A3(_07304_),
    .ZN(_07628_));
 NOR2_X4 _30094_ (.A1(_07526_),
    .A2(_07360_),
    .ZN(_07629_));
 AOI22_X4 _30095_ (.A1(_07552_),
    .A2(_07390_),
    .B1(_07628_),
    .B2(_07629_),
    .ZN(_07630_));
 NOR4_X2 _30096_ (.A1(_07415_),
    .A2(_07380_),
    .A3(_07525_),
    .A4(_07359_),
    .ZN(_07631_));
 NOR2_X1 _30097_ (.A1(_07435_),
    .A2(_07529_),
    .ZN(_07632_));
 NOR3_X4 _30098_ (.A1(_07415_),
    .A2(_07366_),
    .A3(_07403_),
    .ZN(_07633_));
 AOI221_X2 _30099_ (.A(_07397_),
    .B1(_07631_),
    .B2(_07632_),
    .C1(_07633_),
    .C2(_07436_),
    .ZN(_07634_));
 OAI221_X2 _30100_ (.A(_07485_),
    .B1(_07377_),
    .B2(_07375_),
    .C1(_07290_),
    .C2(_06919_),
    .ZN(_07635_));
 OAI33_X1 _30101_ (.A1(_07431_),
    .A2(_07403_),
    .A3(_07468_),
    .B1(_07353_),
    .B2(_07480_),
    .B3(_07635_),
    .ZN(_07636_));
 NOR3_X1 _30102_ (.A1(_07374_),
    .A2(_07403_),
    .A3(_07475_),
    .ZN(_07637_));
 NOR2_X4 _30103_ (.A1(_07435_),
    .A2(_07414_),
    .ZN(_07638_));
 AOI221_X2 _30104_ (.A(_07407_),
    .B1(_07415_),
    .B2(_07636_),
    .C1(_07637_),
    .C2(_07638_),
    .ZN(_07639_));
 OAI21_X2 _30105_ (.A(_07630_),
    .B1(_07634_),
    .B2(_07639_),
    .ZN(_07640_));
 OR2_X4 _30106_ (.A1(_07627_),
    .A2(_07640_),
    .ZN(_07641_));
 OAI21_X2 _30107_ (.A(_07260_),
    .B1(_07613_),
    .B2(_07641_),
    .ZN(_07642_));
 CLKBUF_X3 _30108_ (.A(\core.enc_block.block_w0_reg[26] ),
    .Z(_07643_));
 BUF_X4 _30109_ (.A(\core.enc_block.block_w1_reg[18] ),
    .Z(_07644_));
 BUF_X2 _30110_ (.A(\core.enc_block.block_w3_reg[1] ),
    .Z(_07645_));
 XNOR2_X1 _30111_ (.A(_07644_),
    .B(_07645_),
    .ZN(_07646_));
 XNOR2_X2 _30112_ (.A(_07643_),
    .B(_07646_),
    .ZN(_07647_));
 BUF_X2 _30113_ (.A(\core.enc_block.block_w3_reg[2] ),
    .Z(_07648_));
 XOR2_X1 _30114_ (.A(_00312_),
    .B(_07648_),
    .Z(_07649_));
 XNOR2_X1 _30115_ (.A(_07647_),
    .B(_07649_),
    .ZN(_07650_));
 BUF_X4 _30116_ (.A(_07231_),
    .Z(_07651_));
 MUX2_X2 _30117_ (.A(_07274_),
    .B(_07650_),
    .S(_07651_),
    .Z(_07652_));
 NAND2_X1 _30118_ (.A1(_07229_),
    .A2(_07652_),
    .ZN(_07653_));
 INV_X1 _30119_ (.A(\block_reg[0][10] ),
    .ZN(_07654_));
 OAI21_X1 _30120_ (.A(_07653_),
    .B1(_07248_),
    .B2(_07654_),
    .ZN(_07655_));
 OAI22_X1 _30121_ (.A1(\block_reg[0][10] ),
    .A2(_07251_),
    .B1(_07254_),
    .B2(_07652_),
    .ZN(_07656_));
 MUX2_X2 _30122_ (.A(_07655_),
    .B(_07656_),
    .S(_17739_),
    .Z(_07657_));
 NOR2_X1 _30123_ (.A1(_07224_),
    .A2(_07657_),
    .ZN(_07658_));
 AOI22_X1 _30124_ (.A1(_07259_),
    .A2(_06705_),
    .B1(_07642_),
    .B2(_07658_),
    .ZN(_00703_));
 CLKBUF_X3 _30125_ (.A(\core.enc_block.block_w0_reg[11] ),
    .Z(_07659_));
 INV_X1 _30126_ (.A(_07659_),
    .ZN(_07660_));
 BUF_X4 _30127_ (.A(_06704_),
    .Z(_07661_));
 BUF_X8 _30128_ (.A(_07260_),
    .Z(_07662_));
 BUF_X4 _30129_ (.A(_07505_),
    .Z(_07663_));
 NOR4_X1 _30130_ (.A1(_07427_),
    .A2(_07489_),
    .A3(_07585_),
    .A4(_07663_),
    .ZN(_07664_));
 NOR2_X2 _30131_ (.A1(_07410_),
    .A2(_07374_),
    .ZN(_07665_));
 AOI21_X1 _30132_ (.A(_07664_),
    .B1(_07665_),
    .B2(_07469_),
    .ZN(_07666_));
 NOR3_X4 _30133_ (.A1(_07571_),
    .A2(_07454_),
    .A3(_07475_),
    .ZN(_07667_));
 AOI22_X2 _30134_ (.A1(_07439_),
    .A2(_07445_),
    .B1(_07638_),
    .B2(_07667_),
    .ZN(_07668_));
 AOI21_X2 _30135_ (.A(_07400_),
    .B1(_07666_),
    .B2(_07668_),
    .ZN(_07669_));
 BUF_X4 _30136_ (.A(_07504_),
    .Z(_07670_));
 NOR4_X2 _30137_ (.A1(_07422_),
    .A2(_07451_),
    .A3(_07304_),
    .A4(_07670_),
    .ZN(_07671_));
 AOI221_X2 _30138_ (.A(_07397_),
    .B1(_07487_),
    .B2(_07488_),
    .C1(_07289_),
    .C2(_07383_),
    .ZN(_07672_));
 AOI221_X2 _30139_ (.A(_07671_),
    .B1(_07672_),
    .B2(_07552_),
    .C1(_07390_),
    .C2(_07507_),
    .ZN(_07673_));
 NOR2_X1 _30140_ (.A1(_07457_),
    .A2(_07499_),
    .ZN(_07674_));
 AOI21_X1 _30141_ (.A(_07455_),
    .B1(_07585_),
    .B2(_07418_),
    .ZN(_07675_));
 AOI22_X2 _30142_ (.A1(_07594_),
    .A2(_07674_),
    .B1(_07675_),
    .B2(_07592_),
    .ZN(_07676_));
 OAI21_X2 _30143_ (.A(_07673_),
    .B1(_07676_),
    .B2(_07439_),
    .ZN(_07677_));
 NOR2_X2 _30144_ (.A1(_07473_),
    .A2(_07512_),
    .ZN(_07678_));
 MUX2_X1 _30145_ (.A(_07369_),
    .B(_07545_),
    .S(_07678_),
    .Z(_07679_));
 AND2_X1 _30146_ (.A1(_07569_),
    .A2(_07679_),
    .ZN(_07680_));
 NOR2_X4 _30147_ (.A1(_07436_),
    .A2(_07410_),
    .ZN(_07681_));
 BUF_X4 _30148_ (.A(_07480_),
    .Z(_07682_));
 NOR4_X4 _30149_ (.A1(_07425_),
    .A2(_07682_),
    .A3(_07473_),
    .A4(_07512_),
    .ZN(_07683_));
 NAND2_X1 _30150_ (.A1(_07681_),
    .A2(_07683_),
    .ZN(_07684_));
 NOR3_X1 _30151_ (.A1(_07450_),
    .A2(_07451_),
    .A3(_07459_),
    .ZN(_07685_));
 OAI22_X1 _30152_ (.A1(_07418_),
    .A2(_07489_),
    .B1(_07452_),
    .B2(_07459_),
    .ZN(_07686_));
 AOI21_X1 _30153_ (.A(_07685_),
    .B1(_07686_),
    .B2(_07491_),
    .ZN(_07687_));
 NOR2_X4 _30154_ (.A1(_07397_),
    .A2(_07497_),
    .ZN(_07688_));
 AOI22_X4 _30155_ (.A1(_07474_),
    .A2(_07603_),
    .B1(_07629_),
    .B2(_07688_),
    .ZN(_07689_));
 OAI221_X2 _30156_ (.A(_07684_),
    .B1(_07687_),
    .B2(_07550_),
    .C1(_07689_),
    .C2(_07428_),
    .ZN(_07690_));
 NOR4_X4 _30157_ (.A1(_07669_),
    .A2(_07677_),
    .A3(_07680_),
    .A4(_07690_),
    .ZN(_07691_));
 AOI221_X2 _30158_ (.A(_07417_),
    .B1(_07433_),
    .B2(_07482_),
    .C1(_07561_),
    .C2(_07449_),
    .ZN(_07692_));
 NOR4_X1 _30159_ (.A1(_07438_),
    .A2(_07457_),
    .A3(_07489_),
    .A4(_07452_),
    .ZN(_07693_));
 BUF_X4 _30160_ (.A(_07453_),
    .Z(_07694_));
 NOR3_X2 _30161_ (.A1(_07397_),
    .A2(_07509_),
    .A3(_07694_),
    .ZN(_07695_));
 AOI21_X2 _30162_ (.A(_07693_),
    .B1(_07695_),
    .B2(_07522_),
    .ZN(_07696_));
 AOI21_X2 _30163_ (.A(_07692_),
    .B1(_07696_),
    .B2(_07428_),
    .ZN(_07697_));
 OAI21_X1 _30164_ (.A(_07494_),
    .B1(_07390_),
    .B2(_07638_),
    .ZN(_07698_));
 NOR2_X2 _30165_ (.A1(_07635_),
    .A2(_07670_),
    .ZN(_07699_));
 NOR2_X4 _30166_ (.A1(_07421_),
    .A2(_07346_),
    .ZN(_07700_));
 OAI21_X1 _30167_ (.A(_07699_),
    .B1(_07700_),
    .B2(_07594_),
    .ZN(_07701_));
 NAND2_X1 _30168_ (.A1(_07472_),
    .A2(_07390_),
    .ZN(_07702_));
 NOR2_X2 _30169_ (.A1(_07497_),
    .A2(_07504_),
    .ZN(_07703_));
 NOR3_X4 _30170_ (.A1(_07407_),
    .A2(_07409_),
    .A3(_07496_),
    .ZN(_07704_));
 AOI22_X2 _30171_ (.A1(_07552_),
    .A2(_07703_),
    .B1(_07704_),
    .B2(_07594_),
    .ZN(_07705_));
 NAND4_X2 _30172_ (.A1(_07698_),
    .A2(_07701_),
    .A3(_07702_),
    .A4(_07705_),
    .ZN(_07706_));
 NOR2_X1 _30173_ (.A1(_07491_),
    .A2(_07550_),
    .ZN(_07707_));
 NOR3_X4 _30174_ (.A1(_07381_),
    .A2(_07421_),
    .A3(_07475_),
    .ZN(_07708_));
 OAI21_X1 _30175_ (.A(_07707_),
    .B1(_07708_),
    .B2(_07369_),
    .ZN(_07709_));
 NOR3_X2 _30176_ (.A1(_07416_),
    .A2(_07441_),
    .A3(_07475_),
    .ZN(_07710_));
 AOI21_X1 _30177_ (.A(_07710_),
    .B1(_07513_),
    .B2(_07426_),
    .ZN(_07711_));
 NAND2_X2 _30178_ (.A1(_07438_),
    .A2(_07491_),
    .ZN(_07712_));
 OAI21_X2 _30179_ (.A(_07709_),
    .B1(_07711_),
    .B2(_07712_),
    .ZN(_07713_));
 NOR4_X2 _30180_ (.A1(_07586_),
    .A2(_07578_),
    .A3(_07670_),
    .A4(_07663_),
    .ZN(_07714_));
 BUF_X4 _30181_ (.A(_07353_),
    .Z(_07715_));
 NOR4_X2 _30182_ (.A1(_07595_),
    .A2(_07635_),
    .A3(_07715_),
    .A4(_07360_),
    .ZN(_07716_));
 NOR4_X2 _30183_ (.A1(_07422_),
    .A2(_07451_),
    .A3(_07388_),
    .A4(_07582_),
    .ZN(_07717_));
 NOR4_X2 _30184_ (.A1(_07484_),
    .A2(_07509_),
    .A3(_07499_),
    .A4(_07663_),
    .ZN(_07718_));
 NOR4_X2 _30185_ (.A1(_07714_),
    .A2(_07716_),
    .A3(_07717_),
    .A4(_07718_),
    .ZN(_07719_));
 NOR2_X1 _30186_ (.A1(_07466_),
    .A2(_06934_),
    .ZN(_07720_));
 NOR2_X2 _30187_ (.A1(_07336_),
    .A2(_07720_),
    .ZN(_07721_));
 OAI22_X2 _30188_ (.A1(_07621_),
    .A2(_07459_),
    .B1(_07578_),
    .B2(_07536_),
    .ZN(_07722_));
 NAND3_X1 _30189_ (.A1(_07721_),
    .A2(_07607_),
    .A3(_07722_),
    .ZN(_07723_));
 NAND2_X1 _30190_ (.A1(_07719_),
    .A2(_07723_),
    .ZN(_07724_));
 NOR4_X4 _30191_ (.A1(_07697_),
    .A2(_07706_),
    .A3(_07713_),
    .A4(_07724_),
    .ZN(_07725_));
 NOR2_X1 _30192_ (.A1(_07582_),
    .A2(_07477_),
    .ZN(_07726_));
 AOI22_X1 _30193_ (.A1(_07494_),
    .A2(_07726_),
    .B1(_07699_),
    .B2(_07426_),
    .ZN(_07727_));
 NOR2_X2 _30194_ (.A1(_07398_),
    .A2(_07411_),
    .ZN(_07728_));
 NAND3_X1 _30195_ (.A1(_07463_),
    .A2(_07494_),
    .A3(_07728_),
    .ZN(_07729_));
 NAND2_X1 _30196_ (.A1(_07727_),
    .A2(_07729_),
    .ZN(_07730_));
 NAND3_X1 _30197_ (.A1(_07463_),
    .A2(_07552_),
    .A3(_07412_),
    .ZN(_07731_));
 AOI22_X1 _30198_ (.A1(_07472_),
    .A2(_07463_),
    .B1(_07552_),
    .B2(_07559_),
    .ZN(_07732_));
 OAI21_X1 _30199_ (.A(_07731_),
    .B1(_07732_),
    .B2(_07595_),
    .ZN(_07733_));
 NOR2_X2 _30200_ (.A1(_07730_),
    .A2(_07733_),
    .ZN(_07734_));
 NOR2_X1 _30201_ (.A1(_07452_),
    .A2(_07497_),
    .ZN(_07735_));
 NAND2_X1 _30202_ (.A1(_07398_),
    .A2(_07455_),
    .ZN(_07736_));
 NOR2_X2 _30203_ (.A1(_07415_),
    .A2(_07458_),
    .ZN(_07737_));
 AND2_X1 _30204_ (.A1(_07416_),
    .A2(_07458_),
    .ZN(_07738_));
 OAI221_X2 _30205_ (.A(_07735_),
    .B1(_07736_),
    .B2(_07737_),
    .C1(_07399_),
    .C2(_07738_),
    .ZN(_07739_));
 NOR3_X1 _30206_ (.A1(_07536_),
    .A2(_07621_),
    .A3(_07663_),
    .ZN(_07740_));
 NOR3_X1 _30207_ (.A1(_07411_),
    .A2(_07532_),
    .A3(_07526_),
    .ZN(_07741_));
 NOR2_X4 _30208_ (.A1(_07336_),
    .A2(_07337_),
    .ZN(_07742_));
 NOR3_X1 _30209_ (.A1(_07417_),
    .A2(_07391_),
    .A3(_07742_),
    .ZN(_07743_));
 OAI21_X2 _30210_ (.A(_07740_),
    .B1(_07741_),
    .B2(_07743_),
    .ZN(_07744_));
 NAND2_X2 _30211_ (.A1(_07482_),
    .A2(_07699_),
    .ZN(_07745_));
 NAND3_X4 _30212_ (.A1(_07739_),
    .A2(_07744_),
    .A3(_07745_),
    .ZN(_07746_));
 NAND2_X1 _30213_ (.A1(_07433_),
    .A2(_07562_),
    .ZN(_07747_));
 NOR3_X2 _30214_ (.A1(_07448_),
    .A2(_07694_),
    .A3(_07476_),
    .ZN(_07748_));
 AOI22_X4 _30215_ (.A1(_07383_),
    .A2(_07289_),
    .B1(_07371_),
    .B2(_07485_),
    .ZN(_07749_));
 AOI21_X1 _30216_ (.A(_07748_),
    .B1(_07749_),
    .B2(_07426_),
    .ZN(_07750_));
 OAI21_X1 _30217_ (.A(_07747_),
    .B1(_07750_),
    .B2(_07400_),
    .ZN(_07751_));
 AOI21_X2 _30218_ (.A(_07746_),
    .B1(_07751_),
    .B2(_07428_),
    .ZN(_07752_));
 NAND4_X4 _30219_ (.A1(_07691_),
    .A2(_07725_),
    .A3(_07734_),
    .A4(_07752_),
    .ZN(_07753_));
 NOR3_X1 _30220_ (.A1(_07436_),
    .A2(_07441_),
    .A3(_07392_),
    .ZN(_07754_));
 NOR4_X4 _30221_ (.A1(_07366_),
    .A2(_07453_),
    .A3(_07515_),
    .A4(_07517_),
    .ZN(_07755_));
 NOR4_X2 _30222_ (.A1(_07380_),
    .A2(_07402_),
    .A3(_07403_),
    .A4(_07388_),
    .ZN(_07756_));
 NOR4_X2 _30223_ (.A1(_07506_),
    .A2(_07754_),
    .A3(_07755_),
    .A4(_07756_),
    .ZN(_07757_));
 AOI221_X2 _30224_ (.A(_07344_),
    .B1(_07565_),
    .B2(_07348_),
    .C1(_07357_),
    .C2(_07109_),
    .ZN(_07758_));
 AOI21_X1 _30225_ (.A(_07616_),
    .B1(_07758_),
    .B2(_07408_),
    .ZN(_07759_));
 NAND2_X1 _30226_ (.A1(_07614_),
    .A2(_07564_),
    .ZN(_07760_));
 NOR2_X1 _30227_ (.A1(_07531_),
    .A2(_07620_),
    .ZN(_07761_));
 OAI22_X4 _30228_ (.A1(_07375_),
    .A2(_07377_),
    .B1(_07336_),
    .B2(_07337_),
    .ZN(_07762_));
 NOR3_X1 _30229_ (.A1(_07409_),
    .A2(_07535_),
    .A3(_07762_),
    .ZN(_07763_));
 NOR2_X1 _30230_ (.A1(_07431_),
    .A2(_07504_),
    .ZN(_07764_));
 AOI221_X2 _30231_ (.A(_07374_),
    .B1(_07761_),
    .B2(_07763_),
    .C1(_07764_),
    .C2(_07347_),
    .ZN(_07765_));
 NOR3_X4 _30232_ (.A1(_07431_),
    .A2(_07366_),
    .A3(_07453_),
    .ZN(_07766_));
 AOI221_X2 _30233_ (.A(_07380_),
    .B1(_07551_),
    .B2(_07638_),
    .C1(_07766_),
    .C2(_07415_),
    .ZN(_07767_));
 OAI221_X2 _30234_ (.A(_07757_),
    .B1(_07759_),
    .B2(_07760_),
    .C1(_07765_),
    .C2(_07767_),
    .ZN(_07768_));
 OAI22_X4 _30235_ (.A1(_07351_),
    .A2(_07352_),
    .B1(_07336_),
    .B2(_07337_),
    .ZN(_07769_));
 OAI21_X1 _30236_ (.A(_07769_),
    .B1(_07586_),
    .B2(_07408_),
    .ZN(_07770_));
 NAND3_X1 _30237_ (.A1(_07543_),
    .A2(_07761_),
    .A3(_07770_),
    .ZN(_07771_));
 OAI21_X1 _30238_ (.A(_07491_),
    .B1(_07443_),
    .B2(_07685_),
    .ZN(_07772_));
 AOI21_X2 _30239_ (.A(_07517_),
    .B1(_07771_),
    .B2(_07772_),
    .ZN(_07773_));
 NOR4_X1 _30240_ (.A1(_07530_),
    .A2(_07381_),
    .A3(_07621_),
    .A4(_07499_),
    .ZN(_07774_));
 OAI22_X1 _30241_ (.A1(_07526_),
    .A2(_07537_),
    .B1(_07762_),
    .B2(_07532_),
    .ZN(_07775_));
 NAND2_X1 _30242_ (.A1(_07774_),
    .A2(_07775_),
    .ZN(_07776_));
 NOR2_X4 _30243_ (.A1(_07432_),
    .A2(_07410_),
    .ZN(_07777_));
 NOR2_X2 _30244_ (.A1(_07473_),
    .A2(_07517_),
    .ZN(_07778_));
 AOI22_X2 _30245_ (.A1(_07777_),
    .A2(_07482_),
    .B1(_07507_),
    .B2(_07778_),
    .ZN(_07779_));
 NOR4_X1 _30246_ (.A1(_07448_),
    .A2(_07715_),
    .A3(_07360_),
    .A4(_07499_),
    .ZN(_07780_));
 NOR2_X1 _30247_ (.A1(_07437_),
    .A2(_07670_),
    .ZN(_07781_));
 AOI21_X1 _30248_ (.A(_07780_),
    .B1(_07781_),
    .B2(_07545_),
    .ZN(_07782_));
 OAI221_X2 _30249_ (.A(_07776_),
    .B1(_07779_),
    .B2(_07512_),
    .C1(_07522_),
    .C2(_07782_),
    .ZN(_07783_));
 NOR3_X1 _30250_ (.A1(_07768_),
    .A2(_07773_),
    .A3(_07783_),
    .ZN(_07784_));
 NAND2_X2 _30251_ (.A1(_07434_),
    .A2(_07784_),
    .ZN(_07785_));
 OAI21_X4 _30252_ (.A(_07662_),
    .B1(_07753_),
    .B2(_07785_),
    .ZN(_07786_));
 CLKBUF_X3 _30253_ (.A(_07247_),
    .Z(_07787_));
 BUF_X4 _30254_ (.A(_07253_),
    .Z(_07788_));
 BUF_X4 _30255_ (.A(_07651_),
    .Z(_07789_));
 BUF_X2 _30256_ (.A(\core.enc_block.block_w3_reg[3] ),
    .Z(_07790_));
 CLKBUF_X3 _30257_ (.A(\core.enc_block.block_w3_reg[7] ),
    .Z(_07791_));
 XNOR2_X1 _30258_ (.A(_07338_),
    .B(_07791_),
    .ZN(_07792_));
 XNOR2_X1 _30259_ (.A(_07790_),
    .B(_07792_),
    .ZN(_07793_));
 CLKBUF_X3 _30260_ (.A(\core.enc_block.block_w1_reg[19] ),
    .Z(_07794_));
 CLKBUF_X3 _30261_ (.A(\core.enc_block.block_w0_reg[27] ),
    .Z(_07795_));
 XNOR2_X2 _30262_ (.A(_07794_),
    .B(_07795_),
    .ZN(_07796_));
 XNOR2_X1 _30263_ (.A(_07274_),
    .B(_07648_),
    .ZN(_07797_));
 XNOR2_X1 _30264_ (.A(_07796_),
    .B(_07797_),
    .ZN(_07798_));
 XNOR2_X1 _30265_ (.A(_07793_),
    .B(_07798_),
    .ZN(_07799_));
 NAND2_X1 _30266_ (.A1(_07789_),
    .A2(_07799_),
    .ZN(_07800_));
 BUF_X4 _30267_ (.A(_07232_),
    .Z(_07801_));
 OAI21_X2 _30268_ (.A(_07800_),
    .B1(_07801_),
    .B2(_00313_),
    .ZN(_07802_));
 OAI22_X1 _30269_ (.A1(\block_reg[0][11] ),
    .A2(_07787_),
    .B1(_07788_),
    .B2(_07802_),
    .ZN(_07803_));
 OR2_X1 _30270_ (.A1(_18063_),
    .A2(_07803_),
    .ZN(_07804_));
 NOR3_X4 _30271_ (.A1(_16234_),
    .A2(_16240_),
    .A3(_06690_),
    .ZN(_07805_));
 CLKBUF_X3 _30272_ (.A(_07805_),
    .Z(_07806_));
 BUF_X4 _30273_ (.A(_07806_),
    .Z(_07807_));
 BUF_X4 _30274_ (.A(_07228_),
    .Z(_07808_));
 CLKBUF_X3 _30275_ (.A(_07808_),
    .Z(_07809_));
 AOI22_X1 _30276_ (.A1(\block_reg[0][11] ),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_07802_),
    .ZN(_07810_));
 NAND2_X1 _30277_ (.A1(_18063_),
    .A2(_07810_),
    .ZN(_07811_));
 AOI21_X2 _30278_ (.A(_06704_),
    .B1(_07804_),
    .B2(_07811_),
    .ZN(_07812_));
 AOI22_X1 _30279_ (.A1(_07660_),
    .A2(_07661_),
    .B1(_07786_),
    .B2(_07812_),
    .ZN(_00704_));
 BUF_X2 _30280_ (.A(\core.enc_block.block_w0_reg[12] ),
    .Z(_07813_));
 INV_X1 _30281_ (.A(_07813_),
    .ZN(_07814_));
 OAI221_X2 _30282_ (.A(_07485_),
    .B1(_07271_),
    .B2(_07263_),
    .C1(_07290_),
    .C2(_06887_),
    .ZN(_07815_));
 OAI21_X1 _30283_ (.A(_07815_),
    .B1(_07474_),
    .B2(_07417_),
    .ZN(_07816_));
 NAND3_X1 _30284_ (.A1(_07449_),
    .A2(_07507_),
    .A3(_07816_),
    .ZN(_07817_));
 NOR2_X4 _30285_ (.A1(_07387_),
    .A2(_07581_),
    .ZN(_07818_));
 NOR2_X1 _30286_ (.A1(_07595_),
    .A2(_07663_),
    .ZN(_07819_));
 AOI22_X2 _30287_ (.A1(_07562_),
    .A2(_07818_),
    .B1(_07819_),
    .B2(_07544_),
    .ZN(_07820_));
 NAND2_X2 _30288_ (.A1(_07817_),
    .A2(_07820_),
    .ZN(_07821_));
 NOR3_X1 _30289_ (.A1(_07484_),
    .A2(_07393_),
    .A3(_07381_),
    .ZN(_07822_));
 OAI21_X2 _30290_ (.A(_07437_),
    .B1(_07667_),
    .B2(_07822_),
    .ZN(_07823_));
 NOR4_X2 _30291_ (.A1(_07435_),
    .A2(_07396_),
    .A3(_07420_),
    .A4(_07346_),
    .ZN(_07824_));
 NAND2_X1 _30292_ (.A1(_07397_),
    .A2(_07505_),
    .ZN(_07825_));
 AOI221_X2 _30293_ (.A(_07824_),
    .B1(_07825_),
    .B2(_07562_),
    .C1(_07444_),
    .C2(_07766_),
    .ZN(_07826_));
 AOI21_X4 _30294_ (.A(_07427_),
    .B1(_07823_),
    .B2(_07826_),
    .ZN(_07827_));
 OR2_X4 _30295_ (.A1(_07821_),
    .A2(_07827_),
    .ZN(_07828_));
 NOR2_X4 _30296_ (.A1(_07504_),
    .A2(_07663_),
    .ZN(_07829_));
 AOI222_X2 _30297_ (.A1(_07482_),
    .A2(_07829_),
    .B1(_07594_),
    .B2(_07607_),
    .C1(_07704_),
    .C2(_07368_),
    .ZN(_07830_));
 NOR4_X4 _30298_ (.A1(_07435_),
    .A2(_07414_),
    .A3(_07328_),
    .A4(_07468_),
    .ZN(_07831_));
 AOI21_X1 _30299_ (.A(_07831_),
    .B1(_07533_),
    .B2(_07482_),
    .ZN(_07832_));
 NOR2_X1 _30300_ (.A1(_07415_),
    .A2(_07497_),
    .ZN(_07833_));
 AOI221_X2 _30301_ (.A(_07831_),
    .B1(_07833_),
    .B2(_07551_),
    .C1(_07390_),
    .C2(_07472_),
    .ZN(_07834_));
 OAI221_X2 _30302_ (.A(_07830_),
    .B1(_07832_),
    .B2(_07522_),
    .C1(_07834_),
    .C2(_07399_),
    .ZN(_07835_));
 INV_X1 _30303_ (.A(_07835_),
    .ZN(_07836_));
 NOR3_X2 _30304_ (.A1(_07432_),
    .A2(_07441_),
    .A3(_07475_),
    .ZN(_07837_));
 NAND3_X1 _30305_ (.A1(_07457_),
    .A2(_07728_),
    .A3(_07837_),
    .ZN(_07838_));
 AOI22_X2 _30306_ (.A1(_07417_),
    .A2(_07603_),
    .B1(_07700_),
    .B2(_07569_),
    .ZN(_07839_));
 AOI22_X2 _30307_ (.A1(_07369_),
    .A2(_07681_),
    .B1(_07837_),
    .B2(_07411_),
    .ZN(_07840_));
 OAI221_X2 _30308_ (.A(_07838_),
    .B1(_07839_),
    .B2(_07815_),
    .C1(_07582_),
    .C2(_07840_),
    .ZN(_07841_));
 NOR2_X1 _30309_ (.A1(_07438_),
    .A2(_07426_),
    .ZN(_07842_));
 NOR3_X1 _30310_ (.A1(_07448_),
    .A2(_07472_),
    .A3(_07347_),
    .ZN(_07843_));
 OAI33_X1 _30311_ (.A1(_07586_),
    .A2(_07578_),
    .A3(_07712_),
    .B1(_07842_),
    .B2(_07843_),
    .B3(_07491_),
    .ZN(_07844_));
 AOI21_X2 _30312_ (.A(_07841_),
    .B1(_07844_),
    .B2(_07665_),
    .ZN(_07845_));
 NAND2_X2 _30313_ (.A1(_07609_),
    .A2(_07607_),
    .ZN(_07846_));
 OR2_X1 _30314_ (.A1(_07388_),
    .A2(_07678_),
    .ZN(_07847_));
 AOI221_X2 _30315_ (.A(_07336_),
    .B1(_07356_),
    .B2(_07615_),
    .C1(_07109_),
    .C2(_07349_),
    .ZN(_07848_));
 NAND2_X1 _30316_ (.A1(_07614_),
    .A2(_07848_),
    .ZN(_07849_));
 XNOR2_X1 _30317_ (.A(_07530_),
    .B(_07571_),
    .ZN(_07850_));
 AOI21_X1 _30318_ (.A(_07464_),
    .B1(_07394_),
    .B2(_07850_),
    .ZN(_07851_));
 OAI221_X2 _30319_ (.A(_07846_),
    .B1(_07847_),
    .B2(_07849_),
    .C1(_07550_),
    .C2(_07851_),
    .ZN(_07852_));
 NOR3_X4 _30320_ (.A1(_07328_),
    .A2(_07380_),
    .A3(_07346_),
    .ZN(_07853_));
 OAI221_X2 _30321_ (.A(_07777_),
    .B1(_07361_),
    .B2(_07853_),
    .C1(_07381_),
    .C2(_07397_),
    .ZN(_07854_));
 AOI21_X1 _30322_ (.A(_07633_),
    .B1(_07726_),
    .B2(_07552_),
    .ZN(_07855_));
 NOR2_X4 _30323_ (.A1(_07374_),
    .A2(_07388_),
    .ZN(_07856_));
 OAI21_X1 _30324_ (.A(_07443_),
    .B1(_07829_),
    .B2(_07856_),
    .ZN(_07857_));
 NAND3_X1 _30325_ (.A1(_07854_),
    .A2(_07855_),
    .A3(_07857_),
    .ZN(_07858_));
 NOR2_X1 _30326_ (.A1(_07398_),
    .A2(_07635_),
    .ZN(_07859_));
 NOR3_X1 _30327_ (.A1(_07417_),
    .A2(_07458_),
    .A3(_07476_),
    .ZN(_07860_));
 NOR3_X2 _30328_ (.A1(_07410_),
    .A2(_07715_),
    .A3(_07682_),
    .ZN(_07861_));
 OAI21_X1 _30329_ (.A(_07859_),
    .B1(_07860_),
    .B2(_07861_),
    .ZN(_07862_));
 NOR4_X4 _30330_ (.A1(_07535_),
    .A2(_07525_),
    .A3(_07359_),
    .A4(_07378_),
    .ZN(_07863_));
 NOR3_X1 _30331_ (.A1(_07586_),
    .A2(_07682_),
    .A3(_07517_),
    .ZN(_07864_));
 OAI21_X1 _30332_ (.A(_07582_),
    .B1(_07863_),
    .B2(_07864_),
    .ZN(_07865_));
 NOR3_X1 _30333_ (.A1(_07398_),
    .A2(_07586_),
    .A3(_07682_),
    .ZN(_07866_));
 OAI21_X1 _30334_ (.A(_07390_),
    .B1(_07866_),
    .B2(_07426_),
    .ZN(_07867_));
 NOR2_X1 _30335_ (.A1(_07304_),
    .A2(_07499_),
    .ZN(_07868_));
 OAI22_X2 _30336_ (.A1(_07407_),
    .A2(_07304_),
    .B1(_07815_),
    .B2(_07435_),
    .ZN(_07869_));
 NOR3_X2 _30337_ (.A1(_07409_),
    .A2(_07403_),
    .A3(_07475_),
    .ZN(_07870_));
 AOI222_X2 _30338_ (.A1(_07829_),
    .A2(_07544_),
    .B1(_07594_),
    .B2(_07868_),
    .C1(_07869_),
    .C2(_07870_),
    .ZN(_07871_));
 NAND4_X1 _30339_ (.A1(_07862_),
    .A2(_07865_),
    .A3(_07867_),
    .A4(_07871_),
    .ZN(_07872_));
 NOR4_X2 _30340_ (.A1(_07521_),
    .A2(_07852_),
    .A3(_07858_),
    .A4(_07872_),
    .ZN(_07873_));
 NOR3_X1 _30341_ (.A1(_07450_),
    .A2(_07715_),
    .A3(_07578_),
    .ZN(_07874_));
 OAI21_X1 _30342_ (.A(_07491_),
    .B1(_07347_),
    .B2(_07874_),
    .ZN(_07875_));
 AOI21_X1 _30343_ (.A(_07853_),
    .B1(_07362_),
    .B2(_07444_),
    .ZN(_07876_));
 AOI21_X2 _30344_ (.A(_07550_),
    .B1(_07875_),
    .B2(_07876_),
    .ZN(_07877_));
 AOI222_X2 _30345_ (.A1(_07472_),
    .A2(_07379_),
    .B1(_07389_),
    .B2(_07700_),
    .C1(_07778_),
    .C2(_07544_),
    .ZN(_07878_));
 AOI21_X1 _30346_ (.A(_07594_),
    .B1(_07493_),
    .B2(_07571_),
    .ZN(_07879_));
 NOR3_X1 _30347_ (.A1(_07416_),
    .A2(_07404_),
    .A3(_07362_),
    .ZN(_07880_));
 NOR3_X1 _30348_ (.A1(_07571_),
    .A2(_07421_),
    .A3(_07402_),
    .ZN(_07881_));
 OAI21_X1 _30349_ (.A(_07432_),
    .B1(_07410_),
    .B2(_07881_),
    .ZN(_07882_));
 OAI221_X2 _30350_ (.A(_07878_),
    .B1(_07879_),
    .B2(_07550_),
    .C1(_07880_),
    .C2(_07882_),
    .ZN(_07883_));
 NOR3_X1 _30351_ (.A1(_07381_),
    .A2(_07422_),
    .A3(_07509_),
    .ZN(_07884_));
 NOR2_X1 _30352_ (.A1(_07399_),
    .A2(_07884_),
    .ZN(_07885_));
 NOR3_X1 _30353_ (.A1(_07392_),
    .A2(_07381_),
    .A3(_07421_),
    .ZN(_07886_));
 NOR3_X1 _30354_ (.A1(_07571_),
    .A2(_07425_),
    .A3(_07360_),
    .ZN(_07887_));
 NOR3_X1 _30355_ (.A1(_07408_),
    .A2(_07886_),
    .A3(_07887_),
    .ZN(_07888_));
 NOR3_X2 _30356_ (.A1(_07517_),
    .A2(_07885_),
    .A3(_07888_),
    .ZN(_07889_));
 NOR4_X4 _30357_ (.A1(_07746_),
    .A2(_07877_),
    .A3(_07883_),
    .A4(_07889_),
    .ZN(_07890_));
 NAND4_X4 _30358_ (.A1(_07836_),
    .A2(_07845_),
    .A3(_07873_),
    .A4(_07890_),
    .ZN(_07891_));
 OAI21_X2 _30359_ (.A(_07260_),
    .B1(_07828_),
    .B2(_07891_),
    .ZN(_07892_));
 BUF_X4 _30360_ (.A(_07788_),
    .Z(_07893_));
 OR2_X1 _30361_ (.A1(_00314_),
    .A2(_07651_),
    .ZN(_07894_));
 CLKBUF_X3 _30362_ (.A(\core.enc_block.block_w1_reg[20] ),
    .Z(_07895_));
 XOR2_X2 _30363_ (.A(_07895_),
    .B(\core.enc_block.block_w0_reg[28] ),
    .Z(_07896_));
 BUF_X2 _30364_ (.A(\core.enc_block.block_w3_reg[4] ),
    .Z(_07897_));
 XNOR2_X1 _30365_ (.A(_07283_),
    .B(_07897_),
    .ZN(_07898_));
 XNOR2_X1 _30366_ (.A(_07896_),
    .B(_07898_),
    .ZN(_07899_));
 XNOR2_X1 _30367_ (.A(_07793_),
    .B(_07899_),
    .ZN(_07900_));
 NOR3_X2 _30368_ (.A1(_16240_),
    .A2(_06694_),
    .A3(_16246_),
    .ZN(_07901_));
 BUF_X4 _30369_ (.A(_07901_),
    .Z(_07902_));
 OAI21_X2 _30370_ (.A(_07894_),
    .B1(_07900_),
    .B2(_07902_),
    .ZN(_07903_));
 CLKBUF_X3 _30371_ (.A(_07246_),
    .Z(_07904_));
 CLKBUF_X3 _30372_ (.A(_07904_),
    .Z(_07905_));
 BUF_X4 _30373_ (.A(_07905_),
    .Z(_07906_));
 OAI221_X2 _30374_ (.A(_18325_),
    .B1(_07893_),
    .B2(_07903_),
    .C1(_07906_),
    .C2(\block_reg[0][12] ),
    .ZN(_07907_));
 CLKBUF_X3 _30375_ (.A(_07228_),
    .Z(_07908_));
 NAND2_X1 _30376_ (.A1(_07908_),
    .A2(_07903_),
    .ZN(_07909_));
 OAI21_X1 _30377_ (.A(_07909_),
    .B1(_07787_),
    .B2(_06160_),
    .ZN(_07910_));
 OR2_X1 _30378_ (.A1(_18325_),
    .A2(_07910_),
    .ZN(_07911_));
 AOI21_X4 _30379_ (.A(_06704_),
    .B1(_07907_),
    .B2(_07911_),
    .ZN(_07912_));
 AOI22_X1 _30380_ (.A1(_07814_),
    .A2(_07661_),
    .B1(_07892_),
    .B2(_07912_),
    .ZN(_00705_));
 BUF_X2 _30381_ (.A(\core.enc_block.block_w0_reg[13] ),
    .Z(_07913_));
 INV_X1 _30382_ (.A(_07913_),
    .ZN(_07914_));
 AOI22_X2 _30383_ (.A1(_07544_),
    .A2(_07607_),
    .B1(_07856_),
    .B2(_07594_),
    .ZN(_07915_));
 NOR2_X1 _30384_ (.A1(_07742_),
    .A2(_07421_),
    .ZN(_07916_));
 OAI21_X1 _30385_ (.A(_07523_),
    .B1(_07374_),
    .B2(_07621_),
    .ZN(_07917_));
 AOI22_X2 _30386_ (.A1(_07347_),
    .A2(_07512_),
    .B1(_07916_),
    .B2(_07917_),
    .ZN(_07918_));
 AOI22_X1 _30387_ (.A1(_07531_),
    .A2(_07616_),
    .B1(_07426_),
    .B2(_07512_),
    .ZN(_07919_));
 OAI221_X2 _30388_ (.A(_07915_),
    .B1(_07918_),
    .B2(_07517_),
    .C1(_07919_),
    .C2(_07550_),
    .ZN(_07920_));
 OR2_X1 _30389_ (.A1(_07586_),
    .A2(_07682_),
    .ZN(_07921_));
 NOR4_X1 _30390_ (.A1(_07415_),
    .A2(_07374_),
    .A3(_07421_),
    .A4(_07402_),
    .ZN(_07922_));
 AOI21_X1 _30391_ (.A(_07922_),
    .B1(_07886_),
    .B2(_07416_),
    .ZN(_07923_));
 AOI21_X1 _30392_ (.A(_07437_),
    .B1(_07921_),
    .B2(_07923_),
    .ZN(_07924_));
 OAI21_X1 _30393_ (.A(_07305_),
    .B1(_07362_),
    .B2(_07567_),
    .ZN(_07925_));
 NOR4_X2 _30394_ (.A1(_07328_),
    .A2(_07346_),
    .A3(_07304_),
    .A4(_07504_),
    .ZN(_07926_));
 NOR4_X2 _30395_ (.A1(_07380_),
    .A2(_07353_),
    .A3(_07359_),
    .A4(_07388_),
    .ZN(_07927_));
 NOR4_X4 _30396_ (.A1(_07831_),
    .A2(_07863_),
    .A3(_07926_),
    .A4(_07927_),
    .ZN(_07928_));
 NOR3_X2 _30397_ (.A1(_07410_),
    .A2(_07425_),
    .A3(_07480_),
    .ZN(_07929_));
 NOR3_X1 _30398_ (.A1(_07454_),
    .A2(_07475_),
    .A3(_07378_),
    .ZN(_07930_));
 OAI21_X1 _30399_ (.A(_07571_),
    .B1(_07929_),
    .B2(_07930_),
    .ZN(_07931_));
 NAND3_X1 _30400_ (.A1(_07925_),
    .A2(_07928_),
    .A3(_07931_),
    .ZN(_07932_));
 NOR4_X1 _30401_ (.A1(_07883_),
    .A2(_07920_),
    .A3(_07924_),
    .A4(_07932_),
    .ZN(_07933_));
 NOR4_X1 _30402_ (.A1(_07432_),
    .A2(_07409_),
    .A3(_07535_),
    .A4(_07402_),
    .ZN(_07934_));
 AOI21_X1 _30403_ (.A(_07934_),
    .B1(_07708_),
    .B2(_07448_),
    .ZN(_07935_));
 NOR3_X1 _30404_ (.A1(_07402_),
    .A2(_07403_),
    .A3(_07465_),
    .ZN(_07936_));
 AOI21_X1 _30405_ (.A(_07936_),
    .B1(_07362_),
    .B2(_07465_),
    .ZN(_07937_));
 NOR2_X1 _30406_ (.A1(_07410_),
    .A2(_07531_),
    .ZN(_07938_));
 NAND2_X1 _30407_ (.A1(_07530_),
    .A2(_07512_),
    .ZN(_07939_));
 AOI21_X1 _30408_ (.A(_07737_),
    .B1(_07938_),
    .B2(_07939_),
    .ZN(_07940_));
 NAND2_X1 _30409_ (.A1(_07448_),
    .A2(_07527_),
    .ZN(_07941_));
 OAI221_X2 _30410_ (.A(_07935_),
    .B1(_07937_),
    .B2(_07517_),
    .C1(_07940_),
    .C2(_07941_),
    .ZN(_07942_));
 OAI21_X1 _30411_ (.A(_07621_),
    .B1(_07571_),
    .B2(_07524_),
    .ZN(_07943_));
 NOR2_X1 _30412_ (.A1(_07694_),
    .A2(_07762_),
    .ZN(_07944_));
 NAND3_X1 _30413_ (.A1(_07411_),
    .A2(_07943_),
    .A3(_07944_),
    .ZN(_07945_));
 NOR3_X1 _30414_ (.A1(_07531_),
    .A2(_07509_),
    .A3(_07663_),
    .ZN(_07946_));
 AOI21_X1 _30415_ (.A(_07946_),
    .B1(_07362_),
    .B2(_07433_),
    .ZN(_07947_));
 OAI21_X1 _30416_ (.A(_07945_),
    .B1(_07947_),
    .B2(_07411_),
    .ZN(_07948_));
 NOR3_X1 _30417_ (.A1(_07574_),
    .A2(_07942_),
    .A3(_07948_),
    .ZN(_07949_));
 NOR3_X1 _30418_ (.A1(_07509_),
    .A2(_07458_),
    .A3(_07582_),
    .ZN(_07950_));
 OAI21_X1 _30419_ (.A(_07569_),
    .B1(_07950_),
    .B2(_07481_),
    .ZN(_07951_));
 NOR4_X2 _30420_ (.A1(_07435_),
    .A2(_07403_),
    .A3(_07468_),
    .A4(_07557_),
    .ZN(_07952_));
 NAND3_X1 _30421_ (.A1(_07396_),
    .A2(_07415_),
    .A3(_07380_),
    .ZN(_07953_));
 NOR3_X1 _30422_ (.A1(_07431_),
    .A2(_07425_),
    .A3(_07359_),
    .ZN(_07954_));
 AOI221_X2 _30423_ (.A(_07952_),
    .B1(_07953_),
    .B2(_07954_),
    .C1(_07493_),
    .C2(_07495_),
    .ZN(_07955_));
 NAND2_X1 _30424_ (.A1(_07951_),
    .A2(_07955_),
    .ZN(_07956_));
 OAI21_X1 _30425_ (.A(_07497_),
    .B1(_07749_),
    .B2(_07529_),
    .ZN(_07957_));
 NAND4_X1 _30426_ (.A1(_07416_),
    .A2(_07531_),
    .A3(_07721_),
    .A4(_07957_),
    .ZN(_07958_));
 NOR2_X1 _30427_ (.A1(_07391_),
    .A2(_07742_),
    .ZN(_07959_));
 NAND3_X1 _30428_ (.A1(_07436_),
    .A2(_07530_),
    .A3(_07959_),
    .ZN(_07960_));
 AOI21_X1 _30429_ (.A(_07524_),
    .B1(_07958_),
    .B2(_07960_),
    .ZN(_07961_));
 NOR4_X2 _30430_ (.A1(_07373_),
    .A2(_07566_),
    .A3(_07387_),
    .A4(_07769_),
    .ZN(_07962_));
 OAI33_X1 _30431_ (.A1(_07414_),
    .A2(_07328_),
    .A3(_07742_),
    .B1(_07420_),
    .B2(_07720_),
    .B3(_07336_),
    .ZN(_07963_));
 NOR2_X1 _30432_ (.A1(_07620_),
    .A2(_07635_),
    .ZN(_07964_));
 NOR3_X4 _30433_ (.A1(_07523_),
    .A2(_07353_),
    .A3(_07619_),
    .ZN(_07965_));
 AOI221_X2 _30434_ (.A(_07962_),
    .B1(_07963_),
    .B2(_07964_),
    .C1(_07965_),
    .C2(_07513_),
    .ZN(_07966_));
 OAI21_X1 _30435_ (.A(_07523_),
    .B1(_07620_),
    .B2(_07431_),
    .ZN(_07967_));
 NOR4_X2 _30436_ (.A1(_07409_),
    .A2(_07742_),
    .A3(_07373_),
    .A4(_07420_),
    .ZN(_07968_));
 AOI221_X2 _30437_ (.A(_07368_),
    .B1(_07562_),
    .B2(_07818_),
    .C1(_07967_),
    .C2(_07968_),
    .ZN(_07969_));
 AOI21_X1 _30438_ (.A(_07445_),
    .B1(_07694_),
    .B2(_07848_),
    .ZN(_07970_));
 OAI211_X2 _30439_ (.A(_07966_),
    .B(_07969_),
    .C1(_07970_),
    .C2(_07448_),
    .ZN(_07971_));
 NOR4_X1 _30440_ (.A1(_07768_),
    .A2(_07956_),
    .A3(_07961_),
    .A4(_07971_),
    .ZN(_07972_));
 AND3_X1 _30441_ (.A1(_07933_),
    .A2(_07949_),
    .A3(_07972_),
    .ZN(_07973_));
 BUF_X4 _30442_ (.A(_07973_),
    .Z(_07974_));
 NOR3_X2 _30443_ (.A1(_07536_),
    .A2(_07578_),
    .A3(_07762_),
    .ZN(_07975_));
 NAND3_X1 _30444_ (.A1(_07447_),
    .A2(_07543_),
    .A3(_07975_),
    .ZN(_07976_));
 OAI21_X2 _30445_ (.A(_07715_),
    .B1(_07742_),
    .B2(_07536_),
    .ZN(_07977_));
 NOR3_X1 _30446_ (.A1(_07437_),
    .A2(_07532_),
    .A3(_07524_),
    .ZN(_07978_));
 AOI22_X2 _30447_ (.A1(_07369_),
    .A2(_07749_),
    .B1(_07977_),
    .B2(_07978_),
    .ZN(_07979_));
 AOI21_X1 _30448_ (.A(_07437_),
    .B1(_07487_),
    .B2(_07488_),
    .ZN(_07980_));
 AOI22_X1 _30449_ (.A1(_07369_),
    .A2(_07980_),
    .B1(_07975_),
    .B2(_07427_),
    .ZN(_07981_));
 OAI221_X2 _30450_ (.A(_07976_),
    .B1(_07979_),
    .B2(_07670_),
    .C1(_07981_),
    .C2(_07400_),
    .ZN(_07982_));
 NOR3_X2 _30451_ (.A1(_07432_),
    .A2(_07392_),
    .A3(_07422_),
    .ZN(_07983_));
 NAND4_X4 _30452_ (.A1(_07405_),
    .A2(_07406_),
    .A3(_07371_),
    .A4(_07485_),
    .ZN(_07984_));
 AND2_X1 _30453_ (.A1(_07595_),
    .A2(_07984_),
    .ZN(_07985_));
 AOI22_X2 _30454_ (.A1(_07426_),
    .A2(_07518_),
    .B1(_07983_),
    .B2(_07985_),
    .ZN(_07986_));
 NOR3_X2 _30455_ (.A1(_07381_),
    .A2(_07425_),
    .A3(_07682_),
    .ZN(_07987_));
 NOR4_X2 _30456_ (.A1(_07398_),
    .A2(_07457_),
    .A3(_07694_),
    .A4(_07476_),
    .ZN(_07988_));
 OAI221_X2 _30457_ (.A(_07595_),
    .B1(_07987_),
    .B2(_07988_),
    .C1(_07377_),
    .C2(_07375_),
    .ZN(_07989_));
 NOR3_X2 _30458_ (.A1(_07416_),
    .A2(_07694_),
    .A3(_07476_),
    .ZN(_07990_));
 OAI221_X2 _30459_ (.A(_07749_),
    .B1(_07861_),
    .B2(_07990_),
    .C1(_07271_),
    .C2(_07263_),
    .ZN(_07991_));
 OAI21_X2 _30460_ (.A(_07833_),
    .B1(_07494_),
    .B2(_07404_),
    .ZN(_07992_));
 NAND4_X4 _30461_ (.A1(_07986_),
    .A2(_07989_),
    .A3(_07991_),
    .A4(_07992_),
    .ZN(_07993_));
 NOR3_X2 _30462_ (.A1(_07491_),
    .A2(_07929_),
    .A3(_07990_),
    .ZN(_07994_));
 NOR3_X1 _30463_ (.A1(_07427_),
    .A2(_07586_),
    .A3(_07682_),
    .ZN(_07995_));
 OAI21_X1 _30464_ (.A(_07463_),
    .B1(_07995_),
    .B2(_07399_),
    .ZN(_07996_));
 NOR4_X2 _30465_ (.A1(_07416_),
    .A2(_07441_),
    .A3(_07392_),
    .A4(_07497_),
    .ZN(_07997_));
 AOI221_X2 _30466_ (.A(_07997_),
    .B1(_07495_),
    .B2(_07442_),
    .C1(_07417_),
    .C2(_07510_),
    .ZN(_07998_));
 OAI22_X2 _30467_ (.A1(_07994_),
    .A2(_07996_),
    .B1(_07998_),
    .B2(_07547_),
    .ZN(_07999_));
 NOR4_X4 _30468_ (.A1(_07599_),
    .A2(_07942_),
    .A3(_07993_),
    .A4(_07999_),
    .ZN(_08000_));
 OAI33_X1 _30469_ (.A1(_07484_),
    .A2(_07585_),
    .A3(_07497_),
    .B1(_07663_),
    .B2(_07459_),
    .B3(_07452_),
    .ZN(_08001_));
 INV_X1 _30470_ (.A(_07863_),
    .ZN(_08002_));
 NAND3_X1 _30471_ (.A1(_07399_),
    .A2(_07777_),
    .A3(_07545_),
    .ZN(_08003_));
 NAND2_X1 _30472_ (.A1(_08002_),
    .A2(_08003_),
    .ZN(_08004_));
 AOI221_X2 _30473_ (.A(_07852_),
    .B1(_08001_),
    .B2(_07412_),
    .C1(_08004_),
    .C2(_07522_),
    .ZN(_08005_));
 AOI211_X2 _30474_ (.A(_07441_),
    .B(_07393_),
    .C1(_07582_),
    .C2(_07815_),
    .ZN(_08006_));
 OAI21_X2 _30475_ (.A(_07569_),
    .B1(_07683_),
    .B2(_08006_),
    .ZN(_08007_));
 NOR3_X1 _30476_ (.A1(_07595_),
    .A2(_07418_),
    .A3(_07422_),
    .ZN(_08008_));
 NOR3_X1 _30477_ (.A1(_07440_),
    .A2(_07459_),
    .A3(_07585_),
    .ZN(_08009_));
 OAI21_X2 _30478_ (.A(_07749_),
    .B1(_08008_),
    .B2(_08009_),
    .ZN(_08010_));
 NOR4_X4 _30479_ (.A1(_07437_),
    .A2(_07451_),
    .A3(_07458_),
    .A4(_07670_),
    .ZN(_08011_));
 NOR4_X2 _30480_ (.A1(_07484_),
    .A2(_07393_),
    .A3(_07465_),
    .A4(_07388_),
    .ZN(_08012_));
 NOR4_X2 _30481_ (.A1(_07595_),
    .A2(_07509_),
    .A3(_07454_),
    .A4(_07497_),
    .ZN(_08013_));
 NOR4_X2 _30482_ (.A1(_07595_),
    .A2(_07393_),
    .A3(_07454_),
    .A4(_07304_),
    .ZN(_08014_));
 NOR4_X4 _30483_ (.A1(_08011_),
    .A2(_08012_),
    .A3(_08013_),
    .A4(_08014_),
    .ZN(_08015_));
 NAND3_X2 _30484_ (.A1(_08007_),
    .A2(_08010_),
    .A3(_08015_),
    .ZN(_08016_));
 NAND3_X1 _30485_ (.A1(_07428_),
    .A2(_07522_),
    .A3(_07562_),
    .ZN(_08017_));
 NAND4_X1 _30486_ (.A1(_07547_),
    .A2(_07447_),
    .A3(_07543_),
    .A4(_07561_),
    .ZN(_08018_));
 AOI21_X2 _30487_ (.A(_07439_),
    .B1(_08017_),
    .B2(_08018_),
    .ZN(_08019_));
 NOR2_X1 _30488_ (.A1(_07526_),
    .A2(_07388_),
    .ZN(_08020_));
 NOR3_X1 _30489_ (.A1(_07491_),
    .A2(_07530_),
    .A3(_07566_),
    .ZN(_08021_));
 NOR3_X1 _30490_ (.A1(_07399_),
    .A2(_07536_),
    .A3(_07578_),
    .ZN(_08022_));
 OAI21_X1 _30491_ (.A(_08020_),
    .B1(_08021_),
    .B2(_08022_),
    .ZN(_08023_));
 OAI33_X1 _30492_ (.A1(_07399_),
    .A2(_07450_),
    .A3(_07550_),
    .B1(_07670_),
    .B2(_07463_),
    .B3(_07559_),
    .ZN(_08024_));
 NAND2_X1 _30493_ (.A1(_07700_),
    .A2(_08024_),
    .ZN(_08025_));
 NAND3_X1 _30494_ (.A1(_07721_),
    .A2(_07390_),
    .A3(_07722_),
    .ZN(_08026_));
 NAND3_X2 _30495_ (.A1(_08023_),
    .A2(_08025_),
    .A3(_08026_),
    .ZN(_08027_));
 AOI222_X2 _30496_ (.A1(_07369_),
    .A2(_07305_),
    .B1(_07700_),
    .B2(_07856_),
    .C1(_07704_),
    .C2(_07507_),
    .ZN(_08028_));
 OAI221_X2 _30497_ (.A(_07728_),
    .B1(_07623_),
    .B2(_07748_),
    .C1(_07301_),
    .C2(_07291_),
    .ZN(_08029_));
 NOR3_X1 _30498_ (.A1(_07449_),
    .A2(_07418_),
    .A3(_07459_),
    .ZN(_08030_));
 OAI21_X1 _30499_ (.A(_08030_),
    .B1(_07674_),
    .B2(_07592_),
    .ZN(_08031_));
 AOI222_X2 _30500_ (.A1(_07552_),
    .A2(_07379_),
    .B1(_07347_),
    .B2(_07495_),
    .C1(_07500_),
    .C2(_07404_),
    .ZN(_08032_));
 NAND4_X2 _30501_ (.A1(_08028_),
    .A2(_08029_),
    .A3(_08031_),
    .A4(_08032_),
    .ZN(_08033_));
 NOR4_X4 _30502_ (.A1(_08016_),
    .A2(_08019_),
    .A3(_08027_),
    .A4(_08033_),
    .ZN(_08034_));
 NAND4_X4 _30503_ (.A1(_07734_),
    .A2(_08000_),
    .A3(_08005_),
    .A4(_08034_),
    .ZN(_08035_));
 OR3_X2 _30504_ (.A1(_07974_),
    .A2(_07982_),
    .A3(_08035_),
    .ZN(_08036_));
 NAND2_X2 _30505_ (.A1(_07662_),
    .A2(_08036_),
    .ZN(_08037_));
 BUF_X4 _30506_ (.A(_07231_),
    .Z(_08038_));
 BUF_X4 _30507_ (.A(_08038_),
    .Z(_08039_));
 CLKBUF_X3 _30508_ (.A(\core.enc_block.block_w1_reg[21] ),
    .Z(_08040_));
 CLKBUF_X3 _30509_ (.A(\core.enc_block.block_w0_reg[29] ),
    .Z(_08041_));
 XOR2_X2 _30510_ (.A(_08041_),
    .B(_07897_),
    .Z(_08042_));
 BUF_X2 _30511_ (.A(\core.enc_block.block_w3_reg[5] ),
    .Z(_08043_));
 XNOR2_X1 _30512_ (.A(_00314_),
    .B(_08043_),
    .ZN(_08044_));
 XNOR2_X1 _30513_ (.A(_08042_),
    .B(_08044_),
    .ZN(_08045_));
 XNOR2_X1 _30514_ (.A(_08040_),
    .B(_08045_),
    .ZN(_08046_));
 NAND2_X1 _30515_ (.A1(_08039_),
    .A2(_08046_),
    .ZN(_08047_));
 BUF_X4 _30516_ (.A(_07242_),
    .Z(_08048_));
 OAI21_X2 _30517_ (.A(_08047_),
    .B1(_08048_),
    .B2(_00316_),
    .ZN(_08049_));
 NAND2_X1 _30518_ (.A1(_07229_),
    .A2(_08049_),
    .ZN(_08050_));
 INV_X1 _30519_ (.A(\block_reg[0][13] ),
    .ZN(_08051_));
 OAI21_X1 _30520_ (.A(_08050_),
    .B1(_07248_),
    .B2(_08051_),
    .ZN(_08052_));
 OAI22_X1 _30521_ (.A1(\block_reg[0][13] ),
    .A2(_07251_),
    .B1(_07254_),
    .B2(_08049_),
    .ZN(_08053_));
 MUX2_X2 _30522_ (.A(_08052_),
    .B(_08053_),
    .S(_18409_),
    .Z(_08054_));
 NOR2_X1 _30523_ (.A1(_07224_),
    .A2(_08054_),
    .ZN(_08055_));
 AOI22_X1 _30524_ (.A1(_07914_),
    .A2(_07661_),
    .B1(_08037_),
    .B2(_08055_),
    .ZN(_00706_));
 BUF_X2 _30525_ (.A(\core.enc_block.block_w0_reg[14] ),
    .Z(_08056_));
 INV_X1 _30526_ (.A(_08056_),
    .ZN(_08057_));
 AOI22_X1 _30527_ (.A1(_07488_),
    .A2(_07604_),
    .B1(_07980_),
    .B2(_07561_),
    .ZN(_08058_));
 NOR2_X1 _30528_ (.A1(_07547_),
    .A2(_08058_),
    .ZN(_08059_));
 NAND2_X1 _30529_ (.A1(_07427_),
    .A2(_07853_),
    .ZN(_08060_));
 NAND3_X1 _30530_ (.A1(_07561_),
    .A2(_07487_),
    .A3(_07488_),
    .ZN(_08061_));
 AOI21_X2 _30531_ (.A(_07712_),
    .B1(_08060_),
    .B2(_08061_),
    .ZN(_08062_));
 NOR3_X1 _30532_ (.A1(_07398_),
    .A2(_07715_),
    .A3(_07682_),
    .ZN(_08063_));
 NOR3_X1 _30533_ (.A1(_07411_),
    .A2(_07715_),
    .A3(_07578_),
    .ZN(_08064_));
 OAI21_X1 _30534_ (.A(_07749_),
    .B1(_08063_),
    .B2(_08064_),
    .ZN(_08065_));
 NOR2_X1 _30535_ (.A1(_07443_),
    .A2(_07708_),
    .ZN(_08066_));
 OAI33_X1 _30536_ (.A1(_07398_),
    .A2(_07694_),
    .A3(_07476_),
    .B1(_07715_),
    .B2(_07360_),
    .B3(_07571_),
    .ZN(_08067_));
 AOI22_X2 _30537_ (.A1(_07444_),
    .A2(_07562_),
    .B1(_08067_),
    .B2(_07411_),
    .ZN(_08068_));
 OAI221_X2 _30538_ (.A(_08065_),
    .B1(_08066_),
    .B2(_07378_),
    .C1(_07438_),
    .C2(_08068_),
    .ZN(_08069_));
 NOR4_X4 _30539_ (.A1(_07835_),
    .A2(_08059_),
    .A3(_08062_),
    .A4(_08069_),
    .ZN(_08070_));
 MUX2_X1 _30540_ (.A(_07328_),
    .B(_07421_),
    .S(_07431_),
    .Z(_08071_));
 OR4_X2 _30541_ (.A1(_07410_),
    .A2(_07392_),
    .A3(_07474_),
    .A4(_08071_),
    .ZN(_08072_));
 AOI22_X2 _30542_ (.A1(_07562_),
    .A2(_07607_),
    .B1(_07818_),
    .B2(_07369_),
    .ZN(_08073_));
 NAND3_X1 _30543_ (.A1(_07463_),
    .A2(_07404_),
    .A3(_07412_),
    .ZN(_08074_));
 AOI22_X2 _30544_ (.A1(_07472_),
    .A2(_07856_),
    .B1(_07704_),
    .B2(_07494_),
    .ZN(_08075_));
 NAND4_X2 _30545_ (.A1(_08072_),
    .A2(_08073_),
    .A3(_08074_),
    .A4(_08075_),
    .ZN(_08076_));
 NAND4_X2 _30546_ (.A1(_07577_),
    .A2(_07584_),
    .A3(_07951_),
    .A4(_07955_),
    .ZN(_08077_));
 NOR4_X4 _30547_ (.A1(_07773_),
    .A2(_07783_),
    .A3(_08076_),
    .A4(_08077_),
    .ZN(_08078_));
 NAND2_X1 _30548_ (.A1(_07552_),
    .A2(_07607_),
    .ZN(_08079_));
 AOI21_X1 _30549_ (.A(_07450_),
    .B1(_07507_),
    .B2(_07491_),
    .ZN(_08080_));
 OAI21_X1 _30550_ (.A(_07681_),
    .B1(_07507_),
    .B2(_07443_),
    .ZN(_08081_));
 OAI33_X1 _30551_ (.A1(_07742_),
    .A2(_07524_),
    .A3(_07459_),
    .B1(_07585_),
    .B2(_07694_),
    .B3(_07411_),
    .ZN(_08082_));
 AOI22_X1 _30552_ (.A1(_07547_),
    .A2(_07633_),
    .B1(_08082_),
    .B2(_07474_),
    .ZN(_08083_));
 OAI221_X2 _30553_ (.A(_08079_),
    .B1(_08080_),
    .B2(_08081_),
    .C1(_08083_),
    .C2(_07439_),
    .ZN(_08084_));
 INV_X1 _30554_ (.A(_08084_),
    .ZN(_08085_));
 AOI211_X2 _30555_ (.A(_07454_),
    .B(_07476_),
    .C1(_07465_),
    .C2(_07984_),
    .ZN(_08086_));
 OAI21_X1 _30556_ (.A(_07777_),
    .B1(_08063_),
    .B2(_08086_),
    .ZN(_08087_));
 NOR4_X1 _30557_ (.A1(_07399_),
    .A2(_07393_),
    .A3(_07455_),
    .A4(_07635_),
    .ZN(_08088_));
 NOR3_X1 _30558_ (.A1(_07715_),
    .A2(_07578_),
    .A3(_07304_),
    .ZN(_08089_));
 OAI21_X1 _30559_ (.A(_07447_),
    .B1(_08088_),
    .B2(_08089_),
    .ZN(_08090_));
 NOR4_X2 _30560_ (.A1(_07282_),
    .A2(_07425_),
    .A3(_07480_),
    .A4(_07663_),
    .ZN(_08091_));
 AOI221_X2 _30561_ (.A(_08091_),
    .B1(_07665_),
    .B2(_07469_),
    .C1(_07561_),
    .C2(_07495_),
    .ZN(_08092_));
 NAND4_X2 _30562_ (.A1(_08028_),
    .A2(_08087_),
    .A3(_08090_),
    .A4(_08092_),
    .ZN(_08093_));
 AOI21_X2 _30563_ (.A(_07423_),
    .B1(_07681_),
    .B2(_07567_),
    .ZN(_08094_));
 AOI211_X2 _30564_ (.A(_07391_),
    .B(_07402_),
    .C1(_07435_),
    .C2(_07529_),
    .ZN(_08095_));
 NOR2_X1 _30565_ (.A1(_07448_),
    .A2(_07398_),
    .ZN(_08096_));
 AOI221_X2 _30566_ (.A(_07983_),
    .B1(_08095_),
    .B2(_07408_),
    .C1(_08096_),
    .C2(_07594_),
    .ZN(_08097_));
 OAI22_X4 _30567_ (.A1(_07547_),
    .A2(_08094_),
    .B1(_08097_),
    .B2(_07428_),
    .ZN(_08098_));
 AOI21_X4 _30568_ (.A(_08093_),
    .B1(_08098_),
    .B2(_07543_),
    .ZN(_08099_));
 NAND4_X4 _30569_ (.A1(_08070_),
    .A2(_08078_),
    .A3(_08085_),
    .A4(_08099_),
    .ZN(_08100_));
 OR2_X2 _30570_ (.A1(_07974_),
    .A2(_08100_),
    .ZN(_08101_));
 NAND2_X2 _30571_ (.A1(_07662_),
    .A2(_08101_),
    .ZN(_08102_));
 INV_X1 _30572_ (.A(\block_reg[0][14] ),
    .ZN(_08103_));
 CLKBUF_X3 _30573_ (.A(_07246_),
    .Z(_08104_));
 CLKBUF_X3 _30574_ (.A(_07253_),
    .Z(_08105_));
 CLKBUF_X3 _30575_ (.A(\core.enc_block.block_w1_reg[22] ),
    .Z(_08106_));
 CLKBUF_X3 _30576_ (.A(\core.enc_block.block_w0_reg[30] ),
    .Z(_08107_));
 XNOR2_X2 _30577_ (.A(_08106_),
    .B(_08107_),
    .ZN(_08108_));
 XNOR2_X2 _30578_ (.A(_08043_),
    .B(_08108_),
    .ZN(_08109_));
 BUF_X2 _30579_ (.A(\core.enc_block.block_w3_reg[6] ),
    .Z(_08110_));
 XNOR2_X1 _30580_ (.A(_08110_),
    .B(_00316_),
    .ZN(_08111_));
 XNOR2_X1 _30581_ (.A(_08109_),
    .B(_08111_),
    .ZN(_08112_));
 MUX2_X1 _30582_ (.A(_00317_),
    .B(_08112_),
    .S(_07232_),
    .Z(_08113_));
 OAI22_X1 _30583_ (.A1(_08103_),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_08113_),
    .ZN(_08114_));
 NOR2_X1 _30584_ (.A1(_18477_),
    .A2(_08114_),
    .ZN(_08115_));
 BUF_X4 _30585_ (.A(_07806_),
    .Z(_08116_));
 BUF_X4 _30586_ (.A(_07808_),
    .Z(_08117_));
 AOI22_X1 _30587_ (.A1(_08103_),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_08113_),
    .ZN(_08118_));
 AOI21_X2 _30588_ (.A(_08115_),
    .B1(_08118_),
    .B2(_18477_),
    .ZN(_08119_));
 NOR2_X1 _30589_ (.A1(_07224_),
    .A2(_08119_),
    .ZN(_08120_));
 AOI22_X1 _30590_ (.A1(_08057_),
    .A2(_07661_),
    .B1(_08102_),
    .B2(_08120_),
    .ZN(_00707_));
 BUF_X4 _30591_ (.A(\core.enc_block.block_w0_reg[15] ),
    .Z(_08121_));
 INV_X1 _30592_ (.A(_08121_),
    .ZN(_08122_));
 AND4_X1 _30593_ (.A1(_08028_),
    .A2(_08087_),
    .A3(_08090_),
    .A4(_08092_),
    .ZN(_08123_));
 NAND2_X1 _30594_ (.A1(_07984_),
    .A2(_07633_),
    .ZN(_08124_));
 NOR3_X1 _30595_ (.A1(_07418_),
    .A2(_07450_),
    .A3(_07455_),
    .ZN(_08125_));
 OAI21_X1 _30596_ (.A(_07428_),
    .B1(_07482_),
    .B2(_08125_),
    .ZN(_08126_));
 AOI21_X2 _30597_ (.A(_07439_),
    .B1(_08124_),
    .B2(_08126_),
    .ZN(_08127_));
 AOI221_X2 _30598_ (.A(_07506_),
    .B1(_07778_),
    .B2(_07551_),
    .C1(_07493_),
    .C2(_07500_),
    .ZN(_08128_));
 OAI21_X2 _30599_ (.A(_07681_),
    .B1(_07700_),
    .B2(_07362_),
    .ZN(_08129_));
 NOR3_X1 _30600_ (.A1(_07408_),
    .A2(_07422_),
    .A3(_07509_),
    .ZN(_08130_));
 NOR3_X1 _30601_ (.A1(_07397_),
    .A2(_07353_),
    .A3(_07360_),
    .ZN(_08131_));
 NOR3_X2 _30602_ (.A1(_07457_),
    .A2(_08130_),
    .A3(_08131_),
    .ZN(_08132_));
 OAI211_X4 _30603_ (.A(_07854_),
    .B(_08128_),
    .C1(_08129_),
    .C2(_08132_),
    .ZN(_08133_));
 AOI211_X2 _30604_ (.A(_07393_),
    .B(_07458_),
    .C1(_07477_),
    .C2(_07517_),
    .ZN(_08134_));
 NOR3_X1 _30605_ (.A1(_07455_),
    .A2(_07585_),
    .A3(_07550_),
    .ZN(_08135_));
 OAI21_X1 _30606_ (.A(_07543_),
    .B1(_08134_),
    .B2(_08135_),
    .ZN(_08136_));
 NAND4_X2 _30607_ (.A1(_08007_),
    .A2(_08010_),
    .A3(_08015_),
    .A4(_08136_),
    .ZN(_08137_));
 NOR4_X4 _30608_ (.A1(_07841_),
    .A2(_08127_),
    .A3(_08133_),
    .A4(_08137_),
    .ZN(_08138_));
 OAI22_X1 _30609_ (.A1(_07536_),
    .A2(_07418_),
    .B1(_07452_),
    .B2(_07455_),
    .ZN(_08139_));
 AOI21_X1 _30610_ (.A(_07494_),
    .B1(_08139_),
    .B2(_07984_),
    .ZN(_08140_));
 OAI21_X1 _30611_ (.A(_07638_),
    .B1(_07678_),
    .B2(_07561_),
    .ZN(_08141_));
 OAI211_X2 _30612_ (.A(_07483_),
    .B(_07966_),
    .C1(_08140_),
    .C2(_08141_),
    .ZN(_08142_));
 AOI21_X1 _30613_ (.A(_07667_),
    .B1(_07494_),
    .B2(_07522_),
    .ZN(_08143_));
 NAND2_X1 _30614_ (.A1(_07438_),
    .A2(_07440_),
    .ZN(_08144_));
 AOI22_X2 _30615_ (.A1(_07443_),
    .A2(_07495_),
    .B1(_07628_),
    .B2(_07629_),
    .ZN(_08145_));
 OAI221_X2 _30616_ (.A(_07719_),
    .B1(_08143_),
    .B2(_08144_),
    .C1(_08145_),
    .C2(_07400_),
    .ZN(_08146_));
 OAI21_X1 _30617_ (.A(_07818_),
    .B1(_07482_),
    .B2(_07404_),
    .ZN(_08147_));
 OAI21_X1 _30618_ (.A(_07445_),
    .B1(_07512_),
    .B2(_07438_),
    .ZN(_08148_));
 NAND4_X2 _30619_ (.A1(_07573_),
    .A2(_07846_),
    .A3(_08147_),
    .A4(_08148_),
    .ZN(_08149_));
 AOI21_X2 _30620_ (.A(_07863_),
    .B1(_07777_),
    .B2(_07443_),
    .ZN(_08150_));
 AOI21_X2 _30621_ (.A(_07965_),
    .B1(_07426_),
    .B2(_07433_),
    .ZN(_08151_));
 OAI22_X4 _30622_ (.A1(_07815_),
    .A2(_08150_),
    .B1(_08151_),
    .B2(_07670_),
    .ZN(_08152_));
 NOR4_X4 _30623_ (.A1(_08142_),
    .A2(_08146_),
    .A3(_08149_),
    .A4(_08152_),
    .ZN(_08153_));
 NOR3_X1 _30624_ (.A1(_07450_),
    .A2(_07452_),
    .A3(_07455_),
    .ZN(_08154_));
 OAI21_X1 _30625_ (.A(_07440_),
    .B1(_08154_),
    .B2(_07545_),
    .ZN(_08155_));
 NAND3_X1 _30626_ (.A1(_07400_),
    .A2(_07561_),
    .A3(_07665_),
    .ZN(_08156_));
 AOI21_X2 _30627_ (.A(_07449_),
    .B1(_08155_),
    .B2(_08156_),
    .ZN(_08157_));
 AOI22_X2 _30628_ (.A1(_07482_),
    .A2(_07856_),
    .B1(_07819_),
    .B2(_07347_),
    .ZN(_08158_));
 AOI22_X2 _30629_ (.A1(_07728_),
    .A2(_07766_),
    .B1(_07781_),
    .B2(_07700_),
    .ZN(_08159_));
 AOI22_X1 _30630_ (.A1(_07369_),
    .A2(_07777_),
    .B1(_07564_),
    .B2(_07700_),
    .ZN(_08160_));
 OAI221_X2 _30631_ (.A(_08158_),
    .B1(_08159_),
    .B2(_07522_),
    .C1(_08160_),
    .C2(_07400_),
    .ZN(_08161_));
 NOR3_X2 _30632_ (.A1(_07730_),
    .A2(_08157_),
    .A3(_08161_),
    .ZN(_08162_));
 NAND4_X4 _30633_ (.A1(_08123_),
    .A2(_08138_),
    .A3(_08153_),
    .A4(_08162_),
    .ZN(_08163_));
 NAND2_X2 _30634_ (.A1(_07260_),
    .A2(_08163_),
    .ZN(_08164_));
 BUF_X4 _30635_ (.A(\core.enc_block.block_w1_reg[23] ),
    .Z(_08165_));
 XNOR2_X2 _30636_ (.A(_08165_),
    .B(_07235_),
    .ZN(_08166_));
 XNOR2_X1 _30637_ (.A(_08110_),
    .B(_08166_),
    .ZN(_08167_));
 XOR2_X1 _30638_ (.A(_07791_),
    .B(_00317_),
    .Z(_08168_));
 XNOR2_X1 _30639_ (.A(_08167_),
    .B(_08168_),
    .ZN(_08169_));
 NOR2_X1 _30640_ (.A1(_07902_),
    .A2(_08169_),
    .ZN(_08170_));
 AOI21_X2 _30641_ (.A(_08170_),
    .B1(_07902_),
    .B2(_00315_),
    .ZN(_08171_));
 OAI221_X2 _30642_ (.A(_18549_),
    .B1(_07893_),
    .B2(_08171_),
    .C1(_07906_),
    .C2(\block_reg[0][15] ),
    .ZN(_08172_));
 MUX2_X2 _30643_ (.A(_00198_),
    .B(_18548_),
    .S(_16489_),
    .Z(_08173_));
 AOI22_X1 _30644_ (.A1(\block_reg[0][15] ),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_08171_),
    .ZN(_08174_));
 NAND2_X1 _30645_ (.A1(_08173_),
    .A2(_08174_),
    .ZN(_08175_));
 AOI21_X2 _30646_ (.A(_06704_),
    .B1(_08172_),
    .B2(_08175_),
    .ZN(_08176_));
 AOI22_X1 _30647_ (.A1(_08122_),
    .A2(_07661_),
    .B1(_08164_),
    .B2(_08176_),
    .ZN(_00708_));
 BUF_X4 _30648_ (.A(_06703_),
    .Z(_08177_));
 BUF_X4 _30649_ (.A(\core.enc_block.block_w2_reg[16] ),
    .Z(_08178_));
 AOI21_X1 _30650_ (.A(_06713_),
    .B1(_08178_),
    .B2(_06716_),
    .ZN(_08179_));
 INV_X1 _30651_ (.A(_07238_),
    .ZN(_08180_));
 OAI221_X2 _30652_ (.A(_08179_),
    .B1(_06720_),
    .B2(_08180_),
    .C1(_00424_),
    .C2(_06723_),
    .ZN(_08181_));
 NAND2_X2 _30653_ (.A1(_06701_),
    .A2(_00423_),
    .ZN(_08182_));
 AND4_X1 _30654_ (.A1(_06696_),
    .A2(_06835_),
    .A3(_08181_),
    .A4(_08182_),
    .ZN(_08183_));
 BUF_X4 _30655_ (.A(_08183_),
    .Z(_08184_));
 BUF_X4 _30656_ (.A(\core.enc_block.block_w2_reg[17] ),
    .Z(_08185_));
 AOI21_X1 _30657_ (.A(_06699_),
    .B1(_08185_),
    .B2(_06738_),
    .ZN(_08186_));
 CLKBUF_X3 _30658_ (.A(\core.enc_block.block_w1_reg[17] ),
    .Z(_08187_));
 INV_X1 _30659_ (.A(_08187_),
    .ZN(_08188_));
 OAI221_X2 _30660_ (.A(_08186_),
    .B1(_06750_),
    .B2(_08188_),
    .C1(_00427_),
    .C2(_06723_),
    .ZN(_08189_));
 NAND2_X1 _30661_ (.A1(_06725_),
    .A2(_00426_),
    .ZN(_08190_));
 NAND4_X4 _30662_ (.A1(_06733_),
    .A2(_06711_),
    .A3(_08189_),
    .A4(_08190_),
    .ZN(_08191_));
 BUF_X4 _30663_ (.A(_00425_),
    .Z(_08192_));
 INV_X2 _30664_ (.A(_08192_),
    .ZN(_08193_));
 NAND2_X4 _30665_ (.A1(_08193_),
    .A2(_06786_),
    .ZN(_08194_));
 BUF_X4 _30666_ (.A(\core.keymem.prev_key1_reg[16] ),
    .Z(_08195_));
 AOI221_X2 _30667_ (.A(_08184_),
    .B1(_08191_),
    .B2(_08194_),
    .C1(_08195_),
    .C2(_06938_),
    .ZN(_08196_));
 BUF_X4 _30668_ (.A(_08196_),
    .Z(_08197_));
 BUF_X4 _30669_ (.A(_08197_),
    .Z(_08198_));
 BUF_X4 _30670_ (.A(\core.enc_block.block_w2_reg[18] ),
    .Z(_08199_));
 AOI21_X1 _30671_ (.A(_06699_),
    .B1(_08199_),
    .B2(_06738_),
    .ZN(_08200_));
 INV_X1 _30672_ (.A(_07644_),
    .ZN(_08201_));
 OAI221_X2 _30673_ (.A(_08200_),
    .B1(_06750_),
    .B2(_08201_),
    .C1(_00430_),
    .C2(_06723_),
    .ZN(_08202_));
 NAND2_X1 _30674_ (.A1(_06725_),
    .A2(_00429_),
    .ZN(_08203_));
 NAND4_X4 _30675_ (.A1(_06733_),
    .A2(_06735_),
    .A3(_08202_),
    .A4(_08203_),
    .ZN(_08204_));
 BUF_X4 _30676_ (.A(_00431_),
    .Z(_08205_));
 NOR2_X4 _30677_ (.A1(_08205_),
    .A2(_06711_),
    .ZN(_08206_));
 BUF_X4 _30678_ (.A(\core.enc_block.block_w2_reg[19] ),
    .Z(_08207_));
 AOI21_X1 _30679_ (.A(_06713_),
    .B1(_08207_),
    .B2(_06738_),
    .ZN(_08208_));
 INV_X1 _30680_ (.A(_07794_),
    .ZN(_08209_));
 OAI221_X2 _30681_ (.A(_08208_),
    .B1(_06750_),
    .B2(_08209_),
    .C1(_00433_),
    .C2(_06723_),
    .ZN(_08210_));
 NAND2_X1 _30682_ (.A1(_06725_),
    .A2(_00432_),
    .ZN(_08211_));
 AND4_X1 _30683_ (.A1(_06732_),
    .A2(_06710_),
    .A3(_08210_),
    .A4(_08211_),
    .ZN(_08212_));
 BUF_X8 _30684_ (.A(_08212_),
    .Z(_08213_));
 CLKBUF_X3 _30685_ (.A(_00428_),
    .Z(_08214_));
 OAI221_X2 _30686_ (.A(_08204_),
    .B1(_08206_),
    .B2(_08213_),
    .C1(_07419_),
    .C2(_08214_),
    .ZN(_08215_));
 BUF_X4 _30687_ (.A(_08215_),
    .Z(_08216_));
 BUF_X4 _30688_ (.A(_08216_),
    .Z(_08217_));
 BUF_X4 _30689_ (.A(\core.enc_block.block_w2_reg[20] ),
    .Z(_08218_));
 AOI21_X1 _30690_ (.A(_06699_),
    .B1(_08218_),
    .B2(_06738_),
    .ZN(_08219_));
 INV_X1 _30691_ (.A(_07895_),
    .ZN(_08220_));
 OAI221_X2 _30692_ (.A(_08219_),
    .B1(_06750_),
    .B2(_08220_),
    .C1(_00413_),
    .C2(_16250_),
    .ZN(_08221_));
 NAND2_X1 _30693_ (.A1(_06700_),
    .A2(_00412_),
    .ZN(_08222_));
 AND4_X1 _30694_ (.A1(_06732_),
    .A2(_06734_),
    .A3(_08221_),
    .A4(_08222_),
    .ZN(_08223_));
 BUF_X4 _30695_ (.A(_08223_),
    .Z(_08224_));
 BUF_X4 _30696_ (.A(\core.enc_block.block_w2_reg[21] ),
    .Z(_08225_));
 AOI21_X1 _30697_ (.A(_06699_),
    .B1(_08225_),
    .B2(_06715_),
    .ZN(_08226_));
 INV_X1 _30698_ (.A(_08040_),
    .ZN(_08227_));
 OAI221_X2 _30699_ (.A(_08226_),
    .B1(_06750_),
    .B2(_08227_),
    .C1(_00416_),
    .C2(_16250_),
    .ZN(_08228_));
 NAND2_X2 _30700_ (.A1(_06700_),
    .A2(_00415_),
    .ZN(_08229_));
 NAND4_X4 _30701_ (.A1(_06760_),
    .A2(_06745_),
    .A3(_08228_),
    .A4(_08229_),
    .ZN(_08230_));
 INV_X2 _30702_ (.A(_00414_),
    .ZN(_08231_));
 NAND2_X4 _30703_ (.A1(_08231_),
    .A2(_06786_),
    .ZN(_08232_));
 CLKBUF_X3 _30704_ (.A(\core.keymem.prev_key1_reg[20] ),
    .Z(_08233_));
 AOI221_X2 _30705_ (.A(_08224_),
    .B1(_08230_),
    .B2(_08232_),
    .C1(_08233_),
    .C2(_06841_),
    .ZN(_08234_));
 BUF_X4 _30706_ (.A(_08234_),
    .Z(_08235_));
 BUF_X4 _30707_ (.A(\core.enc_block.block_w2_reg[23] ),
    .Z(_08236_));
 AOI21_X1 _30708_ (.A(_06699_),
    .B1(_08236_),
    .B2(_06738_),
    .ZN(_08237_));
 INV_X1 _30709_ (.A(_08165_),
    .ZN(_08238_));
 OAI221_X2 _30710_ (.A(_08237_),
    .B1(_06750_),
    .B2(_08238_),
    .C1(_00422_),
    .C2(_06723_),
    .ZN(_08239_));
 NAND2_X2 _30711_ (.A1(_06725_),
    .A2(_00421_),
    .ZN(_08240_));
 AND4_X1 _30712_ (.A1(_06732_),
    .A2(_06734_),
    .A3(_08239_),
    .A4(_08240_),
    .ZN(_08241_));
 BUF_X4 _30713_ (.A(_08241_),
    .Z(_08242_));
 CLKBUF_X3 _30714_ (.A(\core.enc_block.block_w2_reg[22] ),
    .Z(_08243_));
 AOI21_X1 _30715_ (.A(_06699_),
    .B1(_08243_),
    .B2(_06715_),
    .ZN(_08244_));
 INV_X1 _30716_ (.A(_08106_),
    .ZN(_08245_));
 OAI221_X2 _30717_ (.A(_08244_),
    .B1(_06750_),
    .B2(_08245_),
    .C1(_00419_),
    .C2(_16250_),
    .ZN(_08246_));
 NAND2_X1 _30718_ (.A1(_06713_),
    .A2(_00418_),
    .ZN(_08247_));
 NAND4_X4 _30719_ (.A1(_06760_),
    .A2(_06835_),
    .A3(_08246_),
    .A4(_08247_),
    .ZN(_08248_));
 OR2_X2 _30720_ (.A1(_00417_),
    .A2(_06835_),
    .ZN(_08249_));
 AOI221_X2 _30721_ (.A(_08242_),
    .B1(_08248_),
    .B2(_08249_),
    .C1(_06810_),
    .C2(\core.keymem.prev_key1_reg[23] ),
    .ZN(_08250_));
 BUF_X4 _30722_ (.A(_08250_),
    .Z(_08251_));
 NAND2_X4 _30723_ (.A1(_08235_),
    .A2(_08251_),
    .ZN(_08252_));
 INV_X4 _30724_ (.A(_08195_),
    .ZN(_08253_));
 NOR2_X4 _30725_ (.A1(_08253_),
    .A2(_07315_),
    .ZN(_08254_));
 OAI221_X2 _30726_ (.A(_08191_),
    .B1(_08254_),
    .B2(_08184_),
    .C1(_06886_),
    .C2(_08192_),
    .ZN(_08255_));
 BUF_X4 _30727_ (.A(_08255_),
    .Z(_08256_));
 BUF_X4 _30728_ (.A(_08256_),
    .Z(_08257_));
 NAND4_X4 _30729_ (.A1(_06733_),
    .A2(_06711_),
    .A3(_08239_),
    .A4(_08240_),
    .ZN(_08258_));
 OR2_X4 _30730_ (.A1(_00420_),
    .A2(_06711_),
    .ZN(_08259_));
 AOI22_X4 _30731_ (.A1(_08258_),
    .A2(_08259_),
    .B1(_08248_),
    .B2(_08249_),
    .ZN(_08260_));
 BUF_X4 _30732_ (.A(_08260_),
    .Z(_08261_));
 AND4_X1 _30733_ (.A1(_06732_),
    .A2(_06734_),
    .A3(_08228_),
    .A4(_08229_),
    .ZN(_08262_));
 BUF_X4 _30734_ (.A(_08262_),
    .Z(_08263_));
 NAND2_X4 _30735_ (.A1(_08233_),
    .A2(_06786_),
    .ZN(_08264_));
 NAND4_X4 _30736_ (.A1(_06696_),
    .A2(_06710_),
    .A3(_08221_),
    .A4(_08222_),
    .ZN(_08265_));
 AOI221_X2 _30737_ (.A(_08263_),
    .B1(_08264_),
    .B2(_08265_),
    .C1(_06810_),
    .C2(_08231_),
    .ZN(_08266_));
 BUF_X4 _30738_ (.A(_08266_),
    .Z(_08267_));
 BUF_X4 _30739_ (.A(_08267_),
    .Z(_08268_));
 NAND2_X4 _30740_ (.A1(_08261_),
    .A2(_08268_),
    .ZN(_08269_));
 NOR2_X4 _30741_ (.A1(_08214_),
    .A2(_06711_),
    .ZN(_08270_));
 AND4_X1 _30742_ (.A1(_06732_),
    .A2(_06710_),
    .A3(_08202_),
    .A4(_08203_),
    .ZN(_08271_));
 BUF_X8 _30743_ (.A(_08271_),
    .Z(_08272_));
 OAI22_X4 _30744_ (.A1(_08270_),
    .A2(_08272_),
    .B1(_08206_),
    .B2(_08213_),
    .ZN(_08273_));
 BUF_X4 _30745_ (.A(_08273_),
    .Z(_08274_));
 OAI33_X1 _30746_ (.A1(_08198_),
    .A2(_08217_),
    .A3(_08252_),
    .B1(_08257_),
    .B2(_08269_),
    .B3(_08274_),
    .ZN(_08275_));
 NAND2_X2 _30747_ (.A1(_08251_),
    .A2(_08268_),
    .ZN(_08276_));
 NOR2_X4 _30748_ (.A1(_08192_),
    .A2(_06779_),
    .ZN(_08277_));
 AND4_X1 _30749_ (.A1(_06732_),
    .A2(_06734_),
    .A3(_08189_),
    .A4(_08190_),
    .ZN(_08278_));
 BUF_X4 _30750_ (.A(_08278_),
    .Z(_08279_));
 NOR2_X4 _30751_ (.A1(_08277_),
    .A2(_08279_),
    .ZN(_08280_));
 BUF_X4 _30752_ (.A(_08280_),
    .Z(_08281_));
 BUF_X4 _30753_ (.A(_08281_),
    .Z(_08282_));
 BUF_X4 _30754_ (.A(_08282_),
    .Z(_08283_));
 OAI21_X1 _30755_ (.A(_08276_),
    .B1(_08252_),
    .B2(_08283_),
    .ZN(_08284_));
 INV_X1 _30756_ (.A(_08214_),
    .ZN(_08285_));
 NAND2_X4 _30757_ (.A1(_08285_),
    .A2(_06786_),
    .ZN(_08286_));
 INV_X1 _30758_ (.A(_08205_),
    .ZN(_08287_));
 NAND2_X4 _30759_ (.A1(_08287_),
    .A2(_06786_),
    .ZN(_08288_));
 NAND4_X4 _30760_ (.A1(_06760_),
    .A2(_06835_),
    .A3(_08210_),
    .A4(_08211_),
    .ZN(_08289_));
 NAND4_X4 _30761_ (.A1(_08286_),
    .A2(_08204_),
    .A3(_08288_),
    .A4(_08289_),
    .ZN(_08290_));
 BUF_X4 _30762_ (.A(_08290_),
    .Z(_08291_));
 NOR2_X1 _30763_ (.A1(_08197_),
    .A2(_08291_),
    .ZN(_08292_));
 INV_X2 _30764_ (.A(\core.keymem.prev_key1_reg[23] ),
    .ZN(_08293_));
 NOR2_X2 _30765_ (.A1(_08293_),
    .A2(_06822_),
    .ZN(_08294_));
 NOR2_X4 _30766_ (.A1(_08242_),
    .A2(_08294_),
    .ZN(_08295_));
 AND4_X1 _30767_ (.A1(_06695_),
    .A2(_06734_),
    .A3(_08246_),
    .A4(_08247_),
    .ZN(_08296_));
 BUF_X4 _30768_ (.A(_08296_),
    .Z(_08297_));
 CLKBUF_X3 _30769_ (.A(\core.keymem.prev_key1_reg[22] ),
    .Z(_08298_));
 INV_X2 _30770_ (.A(_08298_),
    .ZN(_08299_));
 NOR2_X1 _30771_ (.A1(_08299_),
    .A2(_06835_),
    .ZN(_08300_));
 NOR2_X1 _30772_ (.A1(_08297_),
    .A2(_08300_),
    .ZN(_08301_));
 BUF_X4 _30773_ (.A(_08301_),
    .Z(_08302_));
 NAND3_X4 _30774_ (.A1(_08234_),
    .A2(_08295_),
    .A3(_08302_),
    .ZN(_08303_));
 AOI22_X4 _30775_ (.A1(_08232_),
    .A2(_08230_),
    .B1(_08264_),
    .B2(_08265_),
    .ZN(_08304_));
 NAND2_X2 _30776_ (.A1(_08251_),
    .A2(_08304_),
    .ZN(_08305_));
 BUF_X4 _30777_ (.A(_08291_),
    .Z(_08306_));
 OAI22_X1 _30778_ (.A1(_08274_),
    .A2(_08303_),
    .B1(_08305_),
    .B2(_08306_),
    .ZN(_08307_));
 NAND2_X2 _30779_ (.A1(_08194_),
    .A2(_08191_),
    .ZN(_08308_));
 BUF_X4 _30780_ (.A(_08308_),
    .Z(_08309_));
 NAND2_X4 _30781_ (.A1(_08195_),
    .A2(_06786_),
    .ZN(_08310_));
 NAND4_X4 _30782_ (.A1(_06760_),
    .A2(_06745_),
    .A3(_08181_),
    .A4(_08182_),
    .ZN(_08311_));
 NAND2_X4 _30783_ (.A1(_08310_),
    .A2(_08311_),
    .ZN(_08312_));
 NOR2_X4 _30784_ (.A1(_08309_),
    .A2(_08312_),
    .ZN(_08313_));
 AOI221_X2 _30785_ (.A(_08275_),
    .B1(_08284_),
    .B2(_08292_),
    .C1(_08307_),
    .C2(_08313_),
    .ZN(_08314_));
 AOI22_X4 _30786_ (.A1(_08286_),
    .A2(_08204_),
    .B1(_08288_),
    .B2(_08289_),
    .ZN(_08315_));
 NAND4_X1 _30787_ (.A1(_08280_),
    .A2(_08261_),
    .A3(_08267_),
    .A4(_08315_),
    .ZN(_08316_));
 NOR2_X4 _30788_ (.A1(_00414_),
    .A2(_06711_),
    .ZN(_08317_));
 INV_X2 _30789_ (.A(_08233_),
    .ZN(_08318_));
 NOR2_X4 _30790_ (.A1(_08318_),
    .A2(_06735_),
    .ZN(_08319_));
 NOR4_X4 _30791_ (.A1(_08317_),
    .A2(_08263_),
    .A3(_08319_),
    .A4(_08224_),
    .ZN(_08320_));
 AOI221_X2 _30792_ (.A(_08213_),
    .B1(_08204_),
    .B2(_08286_),
    .C1(_08287_),
    .C2(_06938_),
    .ZN(_08321_));
 BUF_X4 _30793_ (.A(_08321_),
    .Z(_08322_));
 NAND4_X1 _30794_ (.A1(_08261_),
    .A2(_08320_),
    .A3(_08322_),
    .A4(_08197_),
    .ZN(_08323_));
 NOR4_X4 _30795_ (.A1(_08277_),
    .A2(_08279_),
    .A3(_08206_),
    .A4(_08213_),
    .ZN(_08324_));
 NAND3_X1 _30796_ (.A1(_08261_),
    .A2(_08324_),
    .A3(_08304_),
    .ZN(_08325_));
 AOI221_X1 _30797_ (.A(_08272_),
    .B1(_08288_),
    .B2(_08289_),
    .C1(_06841_),
    .C2(_08285_),
    .ZN(_08326_));
 CLKBUF_X3 _30798_ (.A(_08326_),
    .Z(_08327_));
 NAND4_X1 _30799_ (.A1(_08295_),
    .A2(_08267_),
    .A3(_08302_),
    .A4(_08327_),
    .ZN(_08328_));
 NAND4_X1 _30800_ (.A1(_08316_),
    .A2(_08323_),
    .A3(_08325_),
    .A4(_08328_),
    .ZN(_08329_));
 OAI221_X2 _30801_ (.A(_08265_),
    .B1(_08263_),
    .B2(_08317_),
    .C1(_08318_),
    .C2(_06822_),
    .ZN(_08330_));
 BUF_X4 _30802_ (.A(_08330_),
    .Z(_08331_));
 NOR2_X4 _30803_ (.A1(_00417_),
    .A2(_06745_),
    .ZN(_08332_));
 OAI221_X2 _30804_ (.A(_08258_),
    .B1(_08297_),
    .B2(_08332_),
    .C1(_06837_),
    .C2(_08293_),
    .ZN(_08333_));
 BUF_X4 _30805_ (.A(_08333_),
    .Z(_08334_));
 NOR2_X4 _30806_ (.A1(_08331_),
    .A2(_08334_),
    .ZN(_08335_));
 AOI221_X1 _30807_ (.A(_08279_),
    .B1(_08310_),
    .B2(_08311_),
    .C1(_06841_),
    .C2(_08193_),
    .ZN(_08336_));
 CLKBUF_X3 _30808_ (.A(_08336_),
    .Z(_08337_));
 NAND2_X2 _30809_ (.A1(_08327_),
    .A2(_08337_),
    .ZN(_08338_));
 NAND2_X2 _30810_ (.A1(_08308_),
    .A2(_08315_),
    .ZN(_08339_));
 NAND3_X1 _30811_ (.A1(_08290_),
    .A2(_08338_),
    .A3(_08339_),
    .ZN(_08340_));
 NAND2_X2 _30812_ (.A1(_08234_),
    .A2(_08260_),
    .ZN(_08341_));
 BUF_X4 _30813_ (.A(_08341_),
    .Z(_08342_));
 NAND2_X4 _30814_ (.A1(_08320_),
    .A2(_08251_),
    .ZN(_08343_));
 NAND2_X1 _30815_ (.A1(_08342_),
    .A2(_08343_),
    .ZN(_08344_));
 NOR2_X4 _30816_ (.A1(_08254_),
    .A2(_08184_),
    .ZN(_08345_));
 OAI221_X2 _30817_ (.A(_08289_),
    .B1(_08272_),
    .B2(_08270_),
    .C1(_08205_),
    .C2(_06822_),
    .ZN(_08346_));
 BUF_X8 _30818_ (.A(_08346_),
    .Z(_08347_));
 OAI221_X2 _30819_ (.A(_08311_),
    .B1(_08272_),
    .B2(_08270_),
    .C1(_08253_),
    .C2(_06887_),
    .ZN(_08348_));
 OAI221_X2 _30820_ (.A(_08289_),
    .B1(_08279_),
    .B2(_08277_),
    .C1(_08205_),
    .C2(_06919_),
    .ZN(_08349_));
 OAI221_X2 _30821_ (.A(_08191_),
    .B1(_08206_),
    .B2(_08213_),
    .C1(_06822_),
    .C2(_08192_),
    .ZN(_08350_));
 AND2_X1 _30822_ (.A1(_08349_),
    .A2(_08350_),
    .ZN(_08351_));
 OAI33_X1 _30823_ (.A1(_08281_),
    .A2(_08345_),
    .A3(_08347_),
    .B1(_08348_),
    .B2(_08351_),
    .B3(_08341_),
    .ZN(_08352_));
 AOI221_X2 _30824_ (.A(_08329_),
    .B1(_08335_),
    .B2(_08340_),
    .C1(_08344_),
    .C2(_08352_),
    .ZN(_08353_));
 NAND2_X2 _30825_ (.A1(_08288_),
    .A2(_08289_),
    .ZN(_08354_));
 BUF_X4 _30826_ (.A(_08354_),
    .Z(_08355_));
 BUF_X4 _30827_ (.A(_08355_),
    .Z(_08356_));
 NOR2_X4 _30828_ (.A1(_08317_),
    .A2(_08263_),
    .ZN(_08357_));
 NAND2_X4 _30829_ (.A1(_08264_),
    .A2(_08265_),
    .ZN(_08358_));
 CLKBUF_X3 _30830_ (.A(_08261_),
    .Z(_08359_));
 NAND2_X1 _30831_ (.A1(_08358_),
    .A2(_08359_),
    .ZN(_08360_));
 NOR2_X4 _30832_ (.A1(_08319_),
    .A2(_08224_),
    .ZN(_08361_));
 BUF_X4 _30833_ (.A(_08295_),
    .Z(_08362_));
 BUF_X4 _30834_ (.A(_08302_),
    .Z(_08363_));
 NAND3_X1 _30835_ (.A1(_08361_),
    .A2(_08362_),
    .A3(_08363_),
    .ZN(_08364_));
 AOI21_X1 _30836_ (.A(_08357_),
    .B1(_08360_),
    .B2(_08364_),
    .ZN(_08365_));
 NAND2_X4 _30837_ (.A1(_08286_),
    .A2(_08204_),
    .ZN(_08366_));
 BUF_X4 _30838_ (.A(_08366_),
    .Z(_08367_));
 NAND2_X4 _30839_ (.A1(_08261_),
    .A2(_08320_),
    .ZN(_08368_));
 NAND2_X1 _30840_ (.A1(_08367_),
    .A2(_08368_),
    .ZN(_08369_));
 OAI22_X4 _30841_ (.A1(_08317_),
    .A2(_08263_),
    .B1(_08319_),
    .B2(_08224_),
    .ZN(_08370_));
 NOR2_X4 _30842_ (.A1(_00420_),
    .A2(_06711_),
    .ZN(_08371_));
 OAI221_X2 _30843_ (.A(_08248_),
    .B1(_08371_),
    .B2(_08242_),
    .C1(_08299_),
    .C2(_07419_),
    .ZN(_08372_));
 NOR2_X2 _30844_ (.A1(_08370_),
    .A2(_08372_),
    .ZN(_08373_));
 BUF_X4 _30845_ (.A(_08373_),
    .Z(_08374_));
 BUF_X4 _30846_ (.A(_08367_),
    .Z(_08375_));
 OAI221_X2 _30847_ (.A(_08356_),
    .B1(_08365_),
    .B2(_08369_),
    .C1(_08374_),
    .C2(_08375_),
    .ZN(_08376_));
 BUF_X4 _30848_ (.A(_08320_),
    .Z(_08377_));
 NAND4_X2 _30849_ (.A1(_08377_),
    .A2(_08362_),
    .A3(_08315_),
    .A4(_08363_),
    .ZN(_08378_));
 NOR4_X4 _30850_ (.A1(_08270_),
    .A2(_08272_),
    .A3(_08206_),
    .A4(_08213_),
    .ZN(_08379_));
 NAND2_X2 _30851_ (.A1(_08309_),
    .A2(_08379_),
    .ZN(_08380_));
 BUF_X4 _30852_ (.A(_08309_),
    .Z(_08381_));
 NAND2_X1 _30853_ (.A1(_08381_),
    .A2(_08327_),
    .ZN(_08382_));
 OAI221_X2 _30854_ (.A(_08378_),
    .B1(_08380_),
    .B2(_08303_),
    .C1(_08252_),
    .C2(_08382_),
    .ZN(_08383_));
 BUF_X4 _30855_ (.A(_08304_),
    .Z(_08384_));
 AOI221_X2 _30856_ (.A(_08297_),
    .B1(_08259_),
    .B2(_08258_),
    .C1(_08298_),
    .C2(_06938_),
    .ZN(_08385_));
 BUF_X4 _30857_ (.A(_08385_),
    .Z(_08386_));
 AOI21_X2 _30858_ (.A(_08355_),
    .B1(_08384_),
    .B2(_08386_),
    .ZN(_08387_));
 NAND2_X2 _30859_ (.A1(_08248_),
    .A2(_08249_),
    .ZN(_08388_));
 NAND2_X1 _30860_ (.A1(_08381_),
    .A2(_08388_),
    .ZN(_08389_));
 NOR4_X4 _30861_ (.A1(_08270_),
    .A2(_08272_),
    .A3(_08242_),
    .A4(_08294_),
    .ZN(_08390_));
 AOI22_X4 _30862_ (.A1(_08286_),
    .A2(_08204_),
    .B1(_08258_),
    .B2(_08259_),
    .ZN(_08391_));
 AOI22_X2 _30863_ (.A1(_08377_),
    .A2(_08390_),
    .B1(_08391_),
    .B2(_08304_),
    .ZN(_08392_));
 NAND2_X2 _30864_ (.A1(_08234_),
    .A2(_08386_),
    .ZN(_08393_));
 BUF_X4 _30865_ (.A(_08312_),
    .Z(_08394_));
 AOI221_X2 _30866_ (.A(_08279_),
    .B1(_08204_),
    .B2(_08286_),
    .C1(_08193_),
    .C2(_07108_),
    .ZN(_08395_));
 NAND2_X1 _30867_ (.A1(_08394_),
    .A2(_08395_),
    .ZN(_08396_));
 OAI221_X2 _30868_ (.A(_08387_),
    .B1(_08389_),
    .B2(_08392_),
    .C1(_08393_),
    .C2(_08396_),
    .ZN(_08397_));
 NAND2_X2 _30869_ (.A1(_08366_),
    .A2(_08309_),
    .ZN(_08398_));
 BUF_X4 _30870_ (.A(_08372_),
    .Z(_08399_));
 BUF_X4 _30871_ (.A(_08399_),
    .Z(_08400_));
 BUF_X4 _30872_ (.A(_08331_),
    .Z(_08401_));
 BUF_X4 _30873_ (.A(_08401_),
    .Z(_08402_));
 OAI221_X2 _30874_ (.A(_08355_),
    .B1(_08398_),
    .B2(_08269_),
    .C1(_08400_),
    .C2(_08402_),
    .ZN(_08403_));
 AOI21_X4 _30875_ (.A(_08383_),
    .B1(_08397_),
    .B2(_08403_),
    .ZN(_08404_));
 NAND4_X4 _30876_ (.A1(_08194_),
    .A2(_08191_),
    .A3(_08310_),
    .A4(_08311_),
    .ZN(_08405_));
 NOR4_X1 _30877_ (.A1(_08401_),
    .A2(_08334_),
    .A3(_08216_),
    .A4(_08405_),
    .ZN(_08406_));
 OR2_X1 _30878_ (.A1(_08297_),
    .A2(_08300_),
    .ZN(_08407_));
 BUF_X4 _30879_ (.A(_08407_),
    .Z(_08408_));
 CLKBUF_X3 _30880_ (.A(_08408_),
    .Z(_08409_));
 NOR3_X1 _30881_ (.A1(_08358_),
    .A2(_08347_),
    .A3(_08409_),
    .ZN(_08410_));
 NAND2_X2 _30882_ (.A1(\core.keymem.prev_key1_reg[23] ),
    .A2(_06810_),
    .ZN(_08411_));
 NAND2_X4 _30883_ (.A1(_08258_),
    .A2(_08411_),
    .ZN(_08412_));
 AOI221_X2 _30884_ (.A(_08279_),
    .B1(_08232_),
    .B2(_08230_),
    .C1(_07108_),
    .C2(_08193_),
    .ZN(_08413_));
 NOR2_X2 _30885_ (.A1(_08242_),
    .A2(_08371_),
    .ZN(_08414_));
 OAI22_X1 _30886_ (.A1(_08357_),
    .A2(_08412_),
    .B1(_08413_),
    .B2(_08414_),
    .ZN(_08415_));
 AOI21_X1 _30887_ (.A(_08406_),
    .B1(_08410_),
    .B2(_08415_),
    .ZN(_08416_));
 OAI22_X2 _30888_ (.A1(_08242_),
    .A2(_08371_),
    .B1(_08297_),
    .B2(_08332_),
    .ZN(_08417_));
 BUF_X4 _30889_ (.A(_08417_),
    .Z(_08418_));
 NAND4_X4 _30890_ (.A1(_08232_),
    .A2(_08230_),
    .A3(_08264_),
    .A4(_08265_),
    .ZN(_08419_));
 NOR3_X1 _30891_ (.A1(_08418_),
    .A2(_08354_),
    .A3(_08419_),
    .ZN(_08420_));
 NOR2_X4 _30892_ (.A1(_08206_),
    .A2(_08213_),
    .ZN(_08421_));
 OAI221_X2 _30893_ (.A(_08230_),
    .B1(_08319_),
    .B2(_08224_),
    .C1(_06757_),
    .C2(_00414_),
    .ZN(_08422_));
 BUF_X4 _30894_ (.A(_08422_),
    .Z(_08423_));
 NOR4_X1 _30895_ (.A1(_08421_),
    .A2(_08412_),
    .A3(_08423_),
    .A4(_08409_),
    .ZN(_08424_));
 OAI21_X1 _30896_ (.A(_08395_),
    .B1(_08420_),
    .B2(_08424_),
    .ZN(_08425_));
 NOR4_X2 _30897_ (.A1(_08308_),
    .A2(_08419_),
    .A3(_08333_),
    .A4(_08290_),
    .ZN(_08426_));
 NOR2_X4 _30898_ (.A1(_08280_),
    .A2(_08290_),
    .ZN(_08427_));
 NOR3_X4 _30899_ (.A1(_08412_),
    .A2(_08422_),
    .A3(_08408_),
    .ZN(_08428_));
 NOR2_X2 _30900_ (.A1(_08331_),
    .A2(_08418_),
    .ZN(_08429_));
 NOR2_X1 _30901_ (.A1(_08273_),
    .A2(_08256_),
    .ZN(_08430_));
 AOI221_X2 _30902_ (.A(_08426_),
    .B1(_08427_),
    .B2(_08428_),
    .C1(_08429_),
    .C2(_08430_),
    .ZN(_08431_));
 OAI33_X1 _30903_ (.A1(_08331_),
    .A2(_08333_),
    .A3(_08346_),
    .B1(_08215_),
    .B2(_08417_),
    .B3(_08361_),
    .ZN(_08432_));
 NOR4_X2 _30904_ (.A1(_08331_),
    .A2(_08346_),
    .A3(_08372_),
    .A4(_08405_),
    .ZN(_08433_));
 NOR2_X2 _30905_ (.A1(_08215_),
    .A2(_08256_),
    .ZN(_08434_));
 NOR3_X4 _30906_ (.A1(_08419_),
    .A2(_08412_),
    .A3(_08408_),
    .ZN(_08435_));
 AOI211_X2 _30907_ (.A(_08432_),
    .B(_08433_),
    .C1(_08434_),
    .C2(_08435_),
    .ZN(_08436_));
 AND4_X1 _30908_ (.A1(_08416_),
    .A2(_08425_),
    .A3(_08431_),
    .A4(_08436_),
    .ZN(_08437_));
 NAND4_X4 _30909_ (.A1(_08353_),
    .A2(_08376_),
    .A3(_08404_),
    .A4(_08437_),
    .ZN(_08438_));
 NAND2_X1 _30910_ (.A1(_08295_),
    .A2(_08301_),
    .ZN(_08439_));
 NAND2_X2 _30911_ (.A1(_08280_),
    .A2(_08379_),
    .ZN(_08440_));
 NOR2_X1 _30912_ (.A1(_08234_),
    .A2(_08267_),
    .ZN(_08441_));
 OAI33_X1 _30913_ (.A1(_08309_),
    .A2(_08343_),
    .A3(_08346_),
    .B1(_08439_),
    .B2(_08440_),
    .B3(_08441_),
    .ZN(_08442_));
 NAND2_X2 _30914_ (.A1(_08232_),
    .A2(_08230_),
    .ZN(_08443_));
 OAI21_X1 _30915_ (.A(_08334_),
    .B1(_08399_),
    .B2(_08443_),
    .ZN(_08444_));
 OAI221_X2 _30916_ (.A(_08343_),
    .B1(_08368_),
    .B2(_08366_),
    .C1(_08280_),
    .C2(_08341_),
    .ZN(_08445_));
 AOI221_X2 _30917_ (.A(_08442_),
    .B1(_08444_),
    .B2(_08358_),
    .C1(_08355_),
    .C2(_08445_),
    .ZN(_08446_));
 NOR3_X4 _30918_ (.A1(_08412_),
    .A2(_08370_),
    .A3(_08408_),
    .ZN(_08447_));
 MUX2_X1 _30919_ (.A(_08373_),
    .B(_08447_),
    .S(_08273_),
    .Z(_08448_));
 AOI22_X4 _30920_ (.A1(_08194_),
    .A2(_08191_),
    .B1(_08310_),
    .B2(_08311_),
    .ZN(_08449_));
 NAND2_X2 _30921_ (.A1(_08322_),
    .A2(_08449_),
    .ZN(_08450_));
 NOR2_X1 _30922_ (.A1(_08450_),
    .A2(_08269_),
    .ZN(_08451_));
 AOI21_X1 _30923_ (.A(_08421_),
    .B1(_08358_),
    .B2(_08308_),
    .ZN(_08452_));
 NAND2_X1 _30924_ (.A1(_08366_),
    .A2(_08357_),
    .ZN(_08453_));
 OAI33_X1 _30925_ (.A1(_08309_),
    .A2(_08342_),
    .A3(_08355_),
    .B1(_08439_),
    .B2(_08452_),
    .B3(_08453_),
    .ZN(_08454_));
 NAND4_X1 _30926_ (.A1(_08261_),
    .A2(_08322_),
    .A3(_08267_),
    .A4(_08197_),
    .ZN(_08455_));
 NAND2_X1 _30927_ (.A1(_08320_),
    .A2(_08385_),
    .ZN(_08456_));
 OAI221_X2 _30928_ (.A(_08455_),
    .B1(_08456_),
    .B2(_08338_),
    .C1(_08450_),
    .C2(_08368_),
    .ZN(_08457_));
 NOR4_X4 _30929_ (.A1(_08448_),
    .A2(_08451_),
    .A3(_08454_),
    .A4(_08457_),
    .ZN(_08458_));
 NOR2_X4 _30930_ (.A1(_08270_),
    .A2(_08272_),
    .ZN(_08459_));
 BUF_X4 _30931_ (.A(_08456_),
    .Z(_08460_));
 NOR2_X1 _30932_ (.A1(_08421_),
    .A2(_08256_),
    .ZN(_08461_));
 OAI21_X2 _30933_ (.A(_08459_),
    .B1(_08460_),
    .B2(_08461_),
    .ZN(_08462_));
 NAND3_X1 _30934_ (.A1(_08281_),
    .A2(_08359_),
    .A3(_08268_),
    .ZN(_08463_));
 AOI22_X4 _30935_ (.A1(_08355_),
    .A2(_08460_),
    .B1(_08463_),
    .B2(_08322_),
    .ZN(_08464_));
 AOI22_X2 _30936_ (.A1(_08261_),
    .A2(_08304_),
    .B1(_08386_),
    .B2(_08235_),
    .ZN(_08465_));
 OAI22_X2 _30937_ (.A1(_08343_),
    .A2(_08348_),
    .B1(_08291_),
    .B2(_08465_),
    .ZN(_08466_));
 BUF_X4 _30938_ (.A(_08309_),
    .Z(_08467_));
 AOI22_X4 _30939_ (.A1(_08462_),
    .A2(_08464_),
    .B1(_08466_),
    .B2(_08467_),
    .ZN(_08468_));
 NAND3_X4 _30940_ (.A1(_08320_),
    .A2(_08295_),
    .A3(_08302_),
    .ZN(_08469_));
 AOI21_X1 _30941_ (.A(_08309_),
    .B1(_08421_),
    .B2(_08312_),
    .ZN(_08470_));
 NOR3_X2 _30942_ (.A1(_08367_),
    .A2(_08469_),
    .A3(_08470_),
    .ZN(_08471_));
 NAND3_X1 _30943_ (.A1(_08357_),
    .A2(_08261_),
    .A3(_08379_),
    .ZN(_08472_));
 NAND4_X1 _30944_ (.A1(_08443_),
    .A2(_08354_),
    .A3(_08295_),
    .A4(_08302_),
    .ZN(_08473_));
 XNOR2_X1 _30945_ (.A(_08366_),
    .B(_08361_),
    .ZN(_08474_));
 OAI221_X2 _30946_ (.A(_08472_),
    .B1(_08473_),
    .B2(_08474_),
    .C1(_08393_),
    .C2(_08440_),
    .ZN(_08475_));
 NAND3_X1 _30947_ (.A1(_08366_),
    .A2(_08235_),
    .A3(_08251_),
    .ZN(_08476_));
 NOR4_X4 _30948_ (.A1(_08270_),
    .A2(_08272_),
    .A3(_08254_),
    .A4(_08184_),
    .ZN(_08477_));
 NAND4_X1 _30949_ (.A1(_08377_),
    .A2(_08362_),
    .A3(_08302_),
    .A4(_08477_),
    .ZN(_08478_));
 AOI21_X2 _30950_ (.A(_08350_),
    .B1(_08476_),
    .B2(_08478_),
    .ZN(_08479_));
 NOR3_X4 _30951_ (.A1(_08366_),
    .A2(_08342_),
    .A3(_08351_),
    .ZN(_08480_));
 NOR4_X4 _30952_ (.A1(_08471_),
    .A2(_08475_),
    .A3(_08479_),
    .A4(_08480_),
    .ZN(_08481_));
 NAND4_X4 _30953_ (.A1(_08446_),
    .A2(_08458_),
    .A3(_08468_),
    .A4(_08481_),
    .ZN(_08482_));
 OAI21_X4 _30954_ (.A(_08314_),
    .B1(_08438_),
    .B2(_08482_),
    .ZN(_08483_));
 BUF_X4 _30955_ (.A(_08345_),
    .Z(_08484_));
 BUF_X4 _30956_ (.A(_08484_),
    .Z(_08485_));
 BUF_X4 _30957_ (.A(_08459_),
    .Z(_08486_));
 BUF_X4 _30958_ (.A(_08486_),
    .Z(_08487_));
 BUF_X4 _30959_ (.A(_08356_),
    .Z(_08488_));
 NOR3_X1 _30960_ (.A1(_08487_),
    .A2(_08488_),
    .A3(_08460_),
    .ZN(_08489_));
 NOR2_X4 _30961_ (.A1(_08419_),
    .A2(_08399_),
    .ZN(_08490_));
 BUF_X4 _30962_ (.A(_08421_),
    .Z(_08491_));
 BUF_X4 _30963_ (.A(_08491_),
    .Z(_08492_));
 MUX2_X1 _30964_ (.A(_08490_),
    .B(_08447_),
    .S(_08492_),
    .Z(_08493_));
 AOI21_X1 _30965_ (.A(_08489_),
    .B1(_08493_),
    .B2(_08487_),
    .ZN(_08494_));
 NOR2_X2 _30966_ (.A1(_08485_),
    .A2(_08494_),
    .ZN(_08495_));
 OAI221_X2 _30967_ (.A(_08311_),
    .B1(_08279_),
    .B2(_08277_),
    .C1(_08253_),
    .C2(_07486_),
    .ZN(_08496_));
 BUF_X4 _30968_ (.A(_08496_),
    .Z(_08497_));
 CLKBUF_X3 _30969_ (.A(_08497_),
    .Z(_08498_));
 AOI22_X1 _30970_ (.A1(_08377_),
    .A2(_08315_),
    .B1(_08384_),
    .B2(_08379_),
    .ZN(_08499_));
 OR3_X1 _30971_ (.A1(_08498_),
    .A2(_08439_),
    .A3(_08499_),
    .ZN(_08500_));
 NOR2_X1 _30972_ (.A1(_08491_),
    .A2(_08477_),
    .ZN(_08501_));
 OAI22_X4 _30973_ (.A1(_08277_),
    .A2(_08279_),
    .B1(_08254_),
    .B2(_08184_),
    .ZN(_08502_));
 BUF_X4 _30974_ (.A(_08502_),
    .Z(_08503_));
 OAI21_X1 _30975_ (.A(_08501_),
    .B1(_08503_),
    .B2(_08486_),
    .ZN(_08504_));
 NOR2_X2 _30976_ (.A1(_08419_),
    .A2(_08334_),
    .ZN(_08505_));
 NOR2_X4 _30977_ (.A1(_08333_),
    .A2(_08370_),
    .ZN(_08506_));
 AOI22_X4 _30978_ (.A1(_08286_),
    .A2(_08204_),
    .B1(_08310_),
    .B2(_08311_),
    .ZN(_08507_));
 OR2_X1 _30979_ (.A1(_08381_),
    .A2(_08507_),
    .ZN(_08508_));
 AOI21_X1 _30980_ (.A(_08505_),
    .B1(_08506_),
    .B2(_08508_),
    .ZN(_08509_));
 NAND2_X4 _30981_ (.A1(_08261_),
    .A2(_08304_),
    .ZN(_08510_));
 NAND2_X4 _30982_ (.A1(_08304_),
    .A2(_08386_),
    .ZN(_08511_));
 MUX2_X1 _30983_ (.A(_08510_),
    .B(_08511_),
    .S(_08257_),
    .Z(_08512_));
 OAI221_X2 _30984_ (.A(_08500_),
    .B1(_08504_),
    .B2(_08509_),
    .C1(_08512_),
    .C2(_08306_),
    .ZN(_08513_));
 BUF_X4 _30985_ (.A(_08381_),
    .Z(_08514_));
 BUF_X4 _30986_ (.A(_08514_),
    .Z(_08515_));
 BUF_X4 _30987_ (.A(_08418_),
    .Z(_08516_));
 BUF_X4 _30988_ (.A(_08419_),
    .Z(_08517_));
 BUF_X4 _30989_ (.A(_08334_),
    .Z(_08518_));
 BUF_X4 _30990_ (.A(_08423_),
    .Z(_08519_));
 BUF_X4 _30991_ (.A(_08367_),
    .Z(_08520_));
 OAI33_X1 _30992_ (.A1(_08515_),
    .A2(_08516_),
    .A3(_08517_),
    .B1(_08518_),
    .B2(_08519_),
    .B3(_08520_),
    .ZN(_08521_));
 NAND2_X1 _30993_ (.A1(_08488_),
    .A2(_08521_),
    .ZN(_08522_));
 BUF_X4 _30994_ (.A(_08379_),
    .Z(_08523_));
 NOR3_X1 _30995_ (.A1(_08283_),
    .A2(_08402_),
    .A3(_08516_),
    .ZN(_08524_));
 OAI21_X1 _30996_ (.A(_08523_),
    .B1(_08524_),
    .B2(_08506_),
    .ZN(_08525_));
 AOI21_X1 _30997_ (.A(_08485_),
    .B1(_08522_),
    .B2(_08525_),
    .ZN(_08526_));
 OR2_X2 _30998_ (.A1(_08513_),
    .A2(_08526_),
    .ZN(_08527_));
 AND2_X1 _30999_ (.A1(_08431_),
    .A2(_08436_),
    .ZN(_08528_));
 NAND2_X1 _31000_ (.A1(_08356_),
    .A2(_08484_),
    .ZN(_08529_));
 OAI33_X1 _31001_ (.A1(_08485_),
    .A2(_08252_),
    .A3(_08306_),
    .B1(_08511_),
    .B2(_08529_),
    .B3(_08487_),
    .ZN(_08530_));
 OAI22_X2 _31002_ (.A1(_08283_),
    .A2(_08469_),
    .B1(_08305_),
    .B2(_08485_),
    .ZN(_08531_));
 AOI22_X4 _31003_ (.A1(_08283_),
    .A2(_08530_),
    .B1(_08531_),
    .B2(_08322_),
    .ZN(_08532_));
 NAND4_X1 _31004_ (.A1(_08357_),
    .A2(_08359_),
    .A3(_08197_),
    .A4(_08523_),
    .ZN(_08533_));
 CLKBUF_X3 _31005_ (.A(_08405_),
    .Z(_08534_));
 OR2_X1 _31006_ (.A1(_08290_),
    .A2(_08534_),
    .ZN(_08535_));
 OAI221_X2 _31007_ (.A(_08533_),
    .B1(_08535_),
    .B2(_08460_),
    .C1(_08396_),
    .C2(_08469_),
    .ZN(_08536_));
 NOR3_X4 _31008_ (.A1(_08331_),
    .A2(_08412_),
    .A3(_08408_),
    .ZN(_08537_));
 OAI222_X2 _31009_ (.A1(_08242_),
    .A2(_08371_),
    .B1(_08297_),
    .B2(_08332_),
    .C1(_08254_),
    .C2(_08184_),
    .ZN(_08538_));
 NOR2_X2 _31010_ (.A1(_08401_),
    .A2(_08538_),
    .ZN(_08539_));
 NOR2_X4 _31011_ (.A1(_08423_),
    .A2(_08399_),
    .ZN(_08540_));
 OR3_X1 _31012_ (.A1(_08537_),
    .A2(_08539_),
    .A3(_08540_),
    .ZN(_08541_));
 BUF_X4 _31013_ (.A(_08281_),
    .Z(_08542_));
 NOR2_X4 _31014_ (.A1(_08542_),
    .A2(_08274_),
    .ZN(_08543_));
 NOR3_X2 _31015_ (.A1(_08309_),
    .A2(_08419_),
    .A3(_08399_),
    .ZN(_08544_));
 BUF_X4 _31016_ (.A(_08412_),
    .Z(_08545_));
 NOR4_X1 _31017_ (.A1(_08545_),
    .A2(_08497_),
    .A3(_08370_),
    .A4(_08409_),
    .ZN(_08546_));
 OR2_X1 _31018_ (.A1(_08544_),
    .A2(_08546_),
    .ZN(_08547_));
 AOI221_X2 _31019_ (.A(_08536_),
    .B1(_08541_),
    .B2(_08543_),
    .C1(_08322_),
    .C2(_08547_),
    .ZN(_08548_));
 AOI21_X1 _31020_ (.A(_08379_),
    .B1(_08315_),
    .B2(_08345_),
    .ZN(_08549_));
 NOR3_X1 _31021_ (.A1(_08542_),
    .A2(_08510_),
    .A3(_08549_),
    .ZN(_08550_));
 BUF_X4 _31022_ (.A(_08347_),
    .Z(_08551_));
 NOR2_X1 _31023_ (.A1(_08467_),
    .A2(_08551_),
    .ZN(_08552_));
 BUF_X4 _31024_ (.A(_08345_),
    .Z(_08553_));
 OAI21_X1 _31025_ (.A(_08342_),
    .B1(_08553_),
    .B2(_08303_),
    .ZN(_08554_));
 BUF_X4 _31026_ (.A(_08327_),
    .Z(_08555_));
 NAND3_X4 _31027_ (.A1(_08295_),
    .A2(_08267_),
    .A3(_08302_),
    .ZN(_08556_));
 NAND2_X2 _31028_ (.A1(_08497_),
    .A2(_08256_),
    .ZN(_08557_));
 OAI22_X2 _31029_ (.A1(_08503_),
    .A2(_08368_),
    .B1(_08556_),
    .B2(_08557_),
    .ZN(_08558_));
 AOI221_X2 _31030_ (.A(_08550_),
    .B1(_08552_),
    .B2(_08554_),
    .C1(_08555_),
    .C2(_08558_),
    .ZN(_08559_));
 NAND4_X4 _31031_ (.A1(_08528_),
    .A2(_08532_),
    .A3(_08548_),
    .A4(_08559_),
    .ZN(_08560_));
 BUF_X4 _31032_ (.A(_08347_),
    .Z(_08561_));
 OAI33_X1 _31033_ (.A1(_08561_),
    .A2(_08198_),
    .A3(_08511_),
    .B1(_08313_),
    .B2(_08303_),
    .B3(_08217_),
    .ZN(_08562_));
 NAND3_X1 _31034_ (.A1(_08394_),
    .A2(_08268_),
    .A3(_08386_),
    .ZN(_08563_));
 BUF_X4 _31035_ (.A(_08394_),
    .Z(_08564_));
 AOI221_X2 _31036_ (.A(_08306_),
    .B1(_08303_),
    .B2(_08563_),
    .C1(_08564_),
    .C2(_08514_),
    .ZN(_08565_));
 NOR3_X2 _31037_ (.A1(_08342_),
    .A2(_08217_),
    .A3(_08337_),
    .ZN(_08566_));
 NOR3_X4 _31038_ (.A1(_08562_),
    .A2(_08565_),
    .A3(_08566_),
    .ZN(_08567_));
 OAI33_X1 _31039_ (.A1(_08516_),
    .A2(_08517_),
    .A3(_08350_),
    .B1(_08519_),
    .B2(_08334_),
    .B3(_08349_),
    .ZN(_08568_));
 AND2_X1 _31040_ (.A1(_08375_),
    .A2(_08568_),
    .ZN(_08569_));
 NAND4_X1 _31041_ (.A1(_08486_),
    .A2(_08542_),
    .A3(_08235_),
    .A4(_08359_),
    .ZN(_08570_));
 OAI21_X1 _31042_ (.A(_08570_),
    .B1(_08303_),
    .B2(_08398_),
    .ZN(_08571_));
 NOR2_X1 _31043_ (.A1(_08356_),
    .A2(_08564_),
    .ZN(_08572_));
 NAND4_X4 _31044_ (.A1(_08194_),
    .A2(_08191_),
    .A3(_08288_),
    .A4(_08289_),
    .ZN(_08573_));
 NAND2_X1 _31045_ (.A1(_08357_),
    .A2(_08356_),
    .ZN(_08574_));
 OAI33_X1 _31046_ (.A1(_08485_),
    .A2(_08573_),
    .A3(_08556_),
    .B1(_08574_),
    .B2(_08498_),
    .B3(_08516_),
    .ZN(_08575_));
 AOI221_X2 _31047_ (.A(_08569_),
    .B1(_08571_),
    .B2(_08572_),
    .C1(_08520_),
    .C2(_08575_),
    .ZN(_08576_));
 NOR3_X2 _31048_ (.A1(_08517_),
    .A2(_08334_),
    .A3(_08347_),
    .ZN(_08577_));
 AND2_X1 _31049_ (.A1(_08313_),
    .A2(_08577_),
    .ZN(_08578_));
 AOI21_X1 _31050_ (.A(_08337_),
    .B1(_08497_),
    .B2(_08366_),
    .ZN(_08579_));
 OAI33_X1 _31051_ (.A1(_08459_),
    .A2(_08460_),
    .A3(_08313_),
    .B1(_08579_),
    .B2(_08399_),
    .B3(_08401_),
    .ZN(_08580_));
 BUF_X4 _31052_ (.A(_08394_),
    .Z(_08581_));
 NAND3_X4 _31053_ (.A1(_08362_),
    .A2(_08304_),
    .A3(_08302_),
    .ZN(_08582_));
 OAI33_X1 _31054_ (.A1(_08581_),
    .A2(_08573_),
    .A3(_08510_),
    .B1(_08582_),
    .B2(_08502_),
    .B3(_08421_),
    .ZN(_08583_));
 AOI221_X2 _31055_ (.A(_08578_),
    .B1(_08580_),
    .B2(_08356_),
    .C1(_08520_),
    .C2(_08583_),
    .ZN(_08584_));
 OAI33_X1 _31056_ (.A1(_08561_),
    .A2(_08498_),
    .A3(_08556_),
    .B1(_08469_),
    .B2(_08367_),
    .B3(_08542_),
    .ZN(_08585_));
 NAND4_X2 _31057_ (.A1(_08355_),
    .A2(_08362_),
    .A3(_08384_),
    .A4(_08363_),
    .ZN(_08586_));
 NOR2_X2 _31058_ (.A1(_08366_),
    .A2(_08345_),
    .ZN(_08587_));
 NAND2_X1 _31059_ (.A1(_08581_),
    .A2(_08322_),
    .ZN(_08588_));
 OAI221_X2 _31060_ (.A(_08282_),
    .B1(_08586_),
    .B2(_08587_),
    .C1(_08588_),
    .C2(_08269_),
    .ZN(_08589_));
 NAND3_X1 _31061_ (.A1(_08268_),
    .A2(_08379_),
    .A3(_08386_),
    .ZN(_08590_));
 NAND2_X1 _31062_ (.A1(_08394_),
    .A2(_08315_),
    .ZN(_08591_));
 OAI221_X2 _31063_ (.A(_08467_),
    .B1(_08581_),
    .B2(_08590_),
    .C1(_08591_),
    .C2(_08276_),
    .ZN(_08592_));
 OAI22_X4 _31064_ (.A1(_08274_),
    .A2(_08252_),
    .B1(_08306_),
    .B2(_08460_),
    .ZN(_08593_));
 AOI221_X2 _31065_ (.A(_08585_),
    .B1(_08589_),
    .B2(_08592_),
    .C1(_08593_),
    .C2(_08198_),
    .ZN(_08594_));
 NAND4_X4 _31066_ (.A1(_08567_),
    .A2(_08576_),
    .A3(_08584_),
    .A4(_08594_),
    .ZN(_08595_));
 OR4_X4 _31067_ (.A1(_08495_),
    .A2(_08527_),
    .A3(_08560_),
    .A4(_08595_),
    .ZN(_08596_));
 NOR2_X2 _31068_ (.A1(_08483_),
    .A2(_08596_),
    .ZN(_08597_));
 NOR2_X2 _31069_ (.A1(_06707_),
    .A2(_08597_),
    .ZN(_08598_));
 CLKBUF_X3 _31070_ (.A(_07228_),
    .Z(_08599_));
 XOR2_X2 _31071_ (.A(_07338_),
    .B(_07237_),
    .Z(_08600_));
 XNOR2_X1 _31072_ (.A(_00361_),
    .B(_08165_),
    .ZN(_08601_));
 XNOR2_X1 _31073_ (.A(_08600_),
    .B(_08601_),
    .ZN(_08602_));
 XNOR2_X1 _31074_ (.A(_07234_),
    .B(_08602_),
    .ZN(_08603_));
 MUX2_X1 _31075_ (.A(_07238_),
    .B(_08603_),
    .S(_07242_),
    .Z(_08604_));
 AOI22_X1 _31076_ (.A1(\block_reg[0][16] ),
    .A2(_07806_),
    .B1(_08599_),
    .B2(_08604_),
    .ZN(_08605_));
 INV_X1 _31077_ (.A(_08605_),
    .ZN(_08606_));
 CLKBUF_X3 _31078_ (.A(_07247_),
    .Z(_08607_));
 CLKBUF_X3 _31079_ (.A(_07253_),
    .Z(_08608_));
 OAI22_X1 _31080_ (.A1(\block_reg[0][16] ),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_08604_),
    .ZN(_08609_));
 MUX2_X1 _31081_ (.A(_08606_),
    .B(_08609_),
    .S(_18870_),
    .Z(_08610_));
 NOR3_X1 _31082_ (.A1(_08177_),
    .A2(_08598_),
    .A3(_08610_),
    .ZN(_08611_));
 CLKBUF_X3 _31083_ (.A(\core.enc_block.block_w0_reg[16] ),
    .Z(_08612_));
 INV_X1 _31084_ (.A(_08612_),
    .ZN(_08613_));
 AOI21_X1 _31085_ (.A(_08611_),
    .B1(_06705_),
    .B2(_08613_),
    .ZN(_00709_));
 BUF_X2 _31086_ (.A(\core.enc_block.block_w0_reg[17] ),
    .Z(_08614_));
 INV_X1 _31087_ (.A(_08614_),
    .ZN(_08615_));
 NAND2_X2 _31088_ (.A1(_08322_),
    .A2(_08502_),
    .ZN(_08616_));
 OAI22_X4 _31089_ (.A1(_08450_),
    .A2(_08269_),
    .B1(_08616_),
    .B2(_08343_),
    .ZN(_08617_));
 NAND2_X1 _31090_ (.A1(_08258_),
    .A2(_08259_),
    .ZN(_08618_));
 NOR2_X4 _31091_ (.A1(_08347_),
    .A2(_08497_),
    .ZN(_08619_));
 OAI221_X2 _31092_ (.A(_08248_),
    .B1(_08224_),
    .B2(_08319_),
    .C1(_08299_),
    .C2(_06888_),
    .ZN(_08620_));
 OAI221_X2 _31093_ (.A(_08265_),
    .B1(_08297_),
    .B2(_08332_),
    .C1(_06888_),
    .C2(_08318_),
    .ZN(_08621_));
 NAND2_X1 _31094_ (.A1(_08620_),
    .A2(_08621_),
    .ZN(_08622_));
 AND4_X1 _31095_ (.A1(_08443_),
    .A2(_08618_),
    .A3(_08619_),
    .A4(_08622_),
    .ZN(_08623_));
 NAND4_X1 _31096_ (.A1(_08459_),
    .A2(_08449_),
    .A3(_08384_),
    .A4(_08386_),
    .ZN(_08624_));
 OR4_X1 _31097_ (.A1(_08309_),
    .A2(_08401_),
    .A3(_08418_),
    .A4(_08507_),
    .ZN(_08625_));
 AOI21_X2 _31098_ (.A(_08491_),
    .B1(_08624_),
    .B2(_08625_),
    .ZN(_08626_));
 NAND2_X4 _31099_ (.A1(_08268_),
    .A2(_08385_),
    .ZN(_08627_));
 NAND3_X4 _31100_ (.A1(_08377_),
    .A2(_08251_),
    .A3(_08197_),
    .ZN(_08628_));
 AOI21_X2 _31101_ (.A(_08274_),
    .B1(_08627_),
    .B2(_08628_),
    .ZN(_08629_));
 NOR4_X4 _31102_ (.A1(_08617_),
    .A2(_08623_),
    .A3(_08626_),
    .A4(_08629_),
    .ZN(_08630_));
 AOI22_X1 _31103_ (.A1(_08280_),
    .A2(_08268_),
    .B1(_08497_),
    .B2(_08235_),
    .ZN(_08631_));
 OAI33_X1 _31104_ (.A1(_08551_),
    .A2(_08498_),
    .A3(_08510_),
    .B1(_08216_),
    .B2(_08400_),
    .B3(_08631_),
    .ZN(_08632_));
 OAI22_X4 _31105_ (.A1(_08277_),
    .A2(_08279_),
    .B1(_08206_),
    .B2(_08213_),
    .ZN(_08633_));
 NOR2_X1 _31106_ (.A1(_08633_),
    .A2(_08587_),
    .ZN(_08634_));
 NOR2_X2 _31107_ (.A1(_08459_),
    .A2(_08312_),
    .ZN(_08635_));
 OAI21_X1 _31108_ (.A(_08305_),
    .B1(_08460_),
    .B2(_08635_),
    .ZN(_08636_));
 NAND4_X1 _31109_ (.A1(_08542_),
    .A2(_08359_),
    .A3(_08553_),
    .A4(_08377_),
    .ZN(_08637_));
 OAI21_X1 _31110_ (.A(_08637_),
    .B1(_08305_),
    .B2(_08484_),
    .ZN(_08638_));
 BUF_X4 _31111_ (.A(_08315_),
    .Z(_08639_));
 AOI221_X2 _31112_ (.A(_08632_),
    .B1(_08634_),
    .B2(_08636_),
    .C1(_08638_),
    .C2(_08639_),
    .ZN(_08640_));
 NOR2_X4 _31113_ (.A1(_08280_),
    .A2(_08215_),
    .ZN(_08641_));
 AOI222_X2 _31114_ (.A1(_08639_),
    .A2(_08435_),
    .B1(_08537_),
    .B2(_08427_),
    .C1(_08641_),
    .C2(_08335_),
    .ZN(_08642_));
 NAND3_X1 _31115_ (.A1(_08639_),
    .A2(_08374_),
    .A3(_08557_),
    .ZN(_08643_));
 MUX2_X1 _31116_ (.A(_08388_),
    .B(_08363_),
    .S(_08486_),
    .Z(_08644_));
 NOR4_X1 _31117_ (.A1(_08402_),
    .A2(_08488_),
    .A3(_08545_),
    .A4(_08534_),
    .ZN(_08645_));
 MUX2_X1 _31118_ (.A(_08388_),
    .B(_08363_),
    .S(_08491_),
    .Z(_08646_));
 NOR4_X1 _31119_ (.A1(_08487_),
    .A2(_08545_),
    .A3(_08519_),
    .A4(_08534_),
    .ZN(_08647_));
 AOI22_X1 _31120_ (.A1(_08644_),
    .A2(_08645_),
    .B1(_08646_),
    .B2(_08647_),
    .ZN(_08648_));
 NOR3_X4 _31121_ (.A1(_08518_),
    .A2(_08519_),
    .A3(_08216_),
    .ZN(_08649_));
 NOR4_X1 _31122_ (.A1(_08402_),
    .A2(_08485_),
    .A3(_08561_),
    .A4(_08400_),
    .ZN(_08650_));
 OAI21_X1 _31123_ (.A(_08283_),
    .B1(_08649_),
    .B2(_08650_),
    .ZN(_08651_));
 AND4_X1 _31124_ (.A1(_08642_),
    .A2(_08643_),
    .A3(_08648_),
    .A4(_08651_),
    .ZN(_08652_));
 NAND4_X4 _31125_ (.A1(_08594_),
    .A2(_08630_),
    .A3(_08640_),
    .A4(_08652_),
    .ZN(_08653_));
 NOR3_X1 _31126_ (.A1(_08485_),
    .A2(_08573_),
    .A3(_08393_),
    .ZN(_08654_));
 NOR3_X1 _31127_ (.A1(_08564_),
    .A2(_08349_),
    .A3(_08511_),
    .ZN(_08655_));
 NOR2_X1 _31128_ (.A1(_08356_),
    .A2(_08449_),
    .ZN(_08656_));
 OAI21_X1 _31129_ (.A(_08486_),
    .B1(_08343_),
    .B2(_08656_),
    .ZN(_08657_));
 NOR3_X1 _31130_ (.A1(_08356_),
    .A2(_08197_),
    .A3(_08460_),
    .ZN(_08658_));
 NOR2_X1 _31131_ (.A1(_08498_),
    .A2(_08586_),
    .ZN(_08659_));
 OAI33_X1 _31132_ (.A1(_08654_),
    .A2(_08655_),
    .A3(_08657_),
    .B1(_08658_),
    .B2(_08659_),
    .B3(_08486_),
    .ZN(_08660_));
 BUF_X4 _31133_ (.A(_08370_),
    .Z(_08661_));
 NOR2_X1 _31134_ (.A1(_08515_),
    .A2(_08661_),
    .ZN(_08662_));
 BUF_X4 _31135_ (.A(_08581_),
    .Z(_08663_));
 NOR3_X1 _31136_ (.A1(_08663_),
    .A2(_08518_),
    .A3(_08561_),
    .ZN(_08664_));
 NOR2_X1 _31137_ (.A1(_08345_),
    .A2(_08216_),
    .ZN(_08665_));
 NOR3_X2 _31138_ (.A1(_08242_),
    .A2(_08371_),
    .A3(_08411_),
    .ZN(_08666_));
 NOR2_X1 _31139_ (.A1(_08409_),
    .A2(_08666_),
    .ZN(_08667_));
 OAI221_X1 _31140_ (.A(_08662_),
    .B1(_08664_),
    .B2(_08665_),
    .C1(_08667_),
    .C2(_08251_),
    .ZN(_08668_));
 NOR2_X1 _31141_ (.A1(_08519_),
    .A2(_08538_),
    .ZN(_08669_));
 OAI21_X1 _31142_ (.A(_08523_),
    .B1(_08546_),
    .B2(_08669_),
    .ZN(_08670_));
 NOR2_X2 _31143_ (.A1(_08418_),
    .A2(_08370_),
    .ZN(_08671_));
 NOR2_X2 _31144_ (.A1(_08401_),
    .A2(_08399_),
    .ZN(_08672_));
 AOI22_X1 _31145_ (.A1(_08671_),
    .A2(_08543_),
    .B1(_08672_),
    .B2(_08427_),
    .ZN(_08673_));
 NOR2_X2 _31146_ (.A1(_08291_),
    .A2(_08534_),
    .ZN(_08674_));
 NOR2_X1 _31147_ (.A1(_08503_),
    .A2(_08217_),
    .ZN(_08675_));
 NOR2_X4 _31148_ (.A1(_08418_),
    .A2(_08419_),
    .ZN(_08676_));
 AOI22_X1 _31149_ (.A1(_08374_),
    .A2(_08674_),
    .B1(_08675_),
    .B2(_08676_),
    .ZN(_08677_));
 AND4_X1 _31150_ (.A1(_08668_),
    .A2(_08670_),
    .A3(_08673_),
    .A4(_08677_),
    .ZN(_08678_));
 NOR2_X1 _31151_ (.A1(_08467_),
    .A2(_08291_),
    .ZN(_08679_));
 NOR2_X2 _31152_ (.A1(_08355_),
    .A2(_08553_),
    .ZN(_08680_));
 AOI222_X2 _31153_ (.A1(_08676_),
    .A2(_08543_),
    .B1(_08679_),
    .B2(_08428_),
    .C1(_08447_),
    .C2(_08680_),
    .ZN(_08681_));
 OR2_X1 _31154_ (.A1(_08390_),
    .A2(_08391_),
    .ZN(_08682_));
 NOR2_X2 _31155_ (.A1(_08297_),
    .A2(_08332_),
    .ZN(_08683_));
 NOR4_X1 _31156_ (.A1(_08683_),
    .A2(_08484_),
    .A3(_08517_),
    .A4(_08573_),
    .ZN(_08684_));
 AOI22_X1 _31157_ (.A1(_08198_),
    .A2(_08649_),
    .B1(_08682_),
    .B2(_08684_),
    .ZN(_08685_));
 NOR4_X1 _31158_ (.A1(_08356_),
    .A2(_08484_),
    .A3(_08518_),
    .A4(_08661_),
    .ZN(_08686_));
 NOR4_X1 _31159_ (.A1(_08545_),
    .A2(_08503_),
    .A3(_08661_),
    .A4(_08409_),
    .ZN(_08687_));
 OAI21_X1 _31160_ (.A(_08487_),
    .B1(_08686_),
    .B2(_08687_),
    .ZN(_08688_));
 NOR2_X1 _31161_ (.A1(_08553_),
    .A2(_08273_),
    .ZN(_08689_));
 AOI211_X2 _31162_ (.A(_08281_),
    .B(_08418_),
    .C1(_08519_),
    .C2(_08401_),
    .ZN(_08690_));
 NOR3_X2 _31163_ (.A1(_08381_),
    .A2(_08517_),
    .A3(_08334_),
    .ZN(_08691_));
 OAI21_X1 _31164_ (.A(_08689_),
    .B1(_08690_),
    .B2(_08691_),
    .ZN(_08692_));
 AND4_X1 _31165_ (.A1(_08681_),
    .A2(_08685_),
    .A3(_08688_),
    .A4(_08692_),
    .ZN(_08693_));
 NAND4_X1 _31166_ (.A1(_08359_),
    .A2(_08449_),
    .A3(_08384_),
    .A4(_08555_),
    .ZN(_08694_));
 NAND2_X1 _31167_ (.A1(_08197_),
    .A2(_08327_),
    .ZN(_08695_));
 OAI21_X1 _31168_ (.A(_08359_),
    .B1(_08268_),
    .B2(_08235_),
    .ZN(_08696_));
 AOI221_X2 _31169_ (.A(_08184_),
    .B1(_08289_),
    .B2(_08288_),
    .C1(_08195_),
    .C2(_07108_),
    .ZN(_08697_));
 NAND2_X1 _31170_ (.A1(_08697_),
    .A2(_08395_),
    .ZN(_08698_));
 OAI221_X2 _31171_ (.A(_08694_),
    .B1(_08695_),
    .B2(_08696_),
    .C1(_08269_),
    .C2(_08698_),
    .ZN(_08699_));
 AOI22_X2 _31172_ (.A1(_08520_),
    .A2(_08449_),
    .B1(_08477_),
    .B2(_08282_),
    .ZN(_08700_));
 NAND3_X1 _31173_ (.A1(_08487_),
    .A2(_08498_),
    .A3(_08257_),
    .ZN(_08701_));
 OAI22_X2 _31174_ (.A1(_08276_),
    .A2(_08700_),
    .B1(_08701_),
    .B2(_08368_),
    .ZN(_08702_));
 AOI211_X2 _31175_ (.A(_08457_),
    .B(_08699_),
    .C1(_08702_),
    .C2(_08492_),
    .ZN(_08703_));
 NAND4_X4 _31176_ (.A1(_08660_),
    .A2(_08678_),
    .A3(_08693_),
    .A4(_08703_),
    .ZN(_08704_));
 OR2_X4 _31177_ (.A1(_08653_),
    .A2(_08704_),
    .ZN(_08705_));
 NOR3_X1 _31178_ (.A1(_08556_),
    .A2(_08507_),
    .A3(_08633_),
    .ZN(_08706_));
 NOR2_X1 _31179_ (.A1(_08303_),
    .A2(_08616_),
    .ZN(_08707_));
 NOR2_X1 _31180_ (.A1(_08706_),
    .A2(_08707_),
    .ZN(_08708_));
 AOI21_X1 _31181_ (.A(_08197_),
    .B1(_08394_),
    .B2(_08459_),
    .ZN(_08709_));
 OAI33_X1 _31182_ (.A1(_08486_),
    .A2(_08467_),
    .A3(_08627_),
    .B1(_08709_),
    .B2(_08402_),
    .B3(_08518_),
    .ZN(_08710_));
 NAND4_X2 _31183_ (.A1(_08345_),
    .A2(_08377_),
    .A3(_08362_),
    .A4(_08302_),
    .ZN(_08711_));
 AOI221_X2 _31184_ (.A(_08459_),
    .B1(_08510_),
    .B2(_08469_),
    .C1(_08711_),
    .C2(_08381_),
    .ZN(_08712_));
 OAI21_X2 _31185_ (.A(_08492_),
    .B1(_08710_),
    .B2(_08712_),
    .ZN(_08713_));
 AND2_X1 _31186_ (.A1(_08708_),
    .A2(_08713_),
    .ZN(_08714_));
 OAI21_X4 _31187_ (.A(_08714_),
    .B1(_08438_),
    .B2(_08482_),
    .ZN(_08715_));
 OAI21_X4 _31188_ (.A(_07662_),
    .B1(_08705_),
    .B2(_08715_),
    .ZN(_08716_));
 XNOR2_X1 _31189_ (.A(_08165_),
    .B(_07238_),
    .ZN(_08717_));
 XNOR2_X2 _31190_ (.A(_07292_),
    .B(_08717_),
    .ZN(_08718_));
 XOR2_X1 _31191_ (.A(_00343_),
    .B(_00364_),
    .Z(_08719_));
 XNOR2_X1 _31192_ (.A(_08600_),
    .B(_08719_),
    .ZN(_08720_));
 XNOR2_X1 _31193_ (.A(_08718_),
    .B(_08720_),
    .ZN(_08721_));
 BUF_X4 _31194_ (.A(_07231_),
    .Z(_08722_));
 MUX2_X1 _31195_ (.A(_08187_),
    .B(_08721_),
    .S(_08722_),
    .Z(_08723_));
 OAI22_X1 _31196_ (.A1(\block_reg[0][17] ),
    .A2(_07787_),
    .B1(_07788_),
    .B2(_08723_),
    .ZN(_08724_));
 OR2_X1 _31197_ (.A1(_19191_),
    .A2(_08724_),
    .ZN(_08725_));
 AOI22_X1 _31198_ (.A1(\block_reg[0][17] ),
    .A2(_07807_),
    .B1(_08117_),
    .B2(_08723_),
    .ZN(_08726_));
 NAND2_X1 _31199_ (.A1(_19191_),
    .A2(_08726_),
    .ZN(_08727_));
 AOI21_X2 _31200_ (.A(_06704_),
    .B1(_08725_),
    .B2(_08727_),
    .ZN(_08728_));
 AOI22_X1 _31201_ (.A1(_08615_),
    .A2(_07661_),
    .B1(_08716_),
    .B2(_08728_),
    .ZN(_00710_));
 CLKBUF_X3 _31202_ (.A(\core.enc_block.block_w0_reg[18] ),
    .Z(_08729_));
 INV_X1 _31203_ (.A(_08729_),
    .ZN(_08730_));
 NOR2_X4 _31204_ (.A1(_08418_),
    .A2(_08423_),
    .ZN(_08731_));
 OAI33_X1 _31205_ (.A1(_08519_),
    .A2(_08573_),
    .A3(_08538_),
    .B1(_08633_),
    .B2(_08400_),
    .B3(_08517_),
    .ZN(_08732_));
 AOI22_X4 _31206_ (.A1(_08731_),
    .A2(_08543_),
    .B1(_08732_),
    .B2(_08487_),
    .ZN(_08733_));
 AND3_X1 _31207_ (.A1(_08416_),
    .A2(_08425_),
    .A3(_08733_),
    .ZN(_08734_));
 OAI33_X1 _31208_ (.A1(_08510_),
    .A2(_08306_),
    .A3(_08534_),
    .B1(_08582_),
    .B2(_08484_),
    .B3(_08573_),
    .ZN(_08735_));
 AOI22_X1 _31209_ (.A1(_08251_),
    .A2(_08268_),
    .B1(_08386_),
    .B2(_08235_),
    .ZN(_08736_));
 OAI21_X1 _31210_ (.A(_08325_),
    .B1(_08257_),
    .B2(_08736_),
    .ZN(_08737_));
 NAND4_X1 _31211_ (.A1(_08514_),
    .A2(_08356_),
    .A3(_08251_),
    .A4(_08268_),
    .ZN(_08738_));
 OAI21_X1 _31212_ (.A(_08738_),
    .B1(_08582_),
    .B2(_08515_),
    .ZN(_08739_));
 AOI221_X2 _31213_ (.A(_08735_),
    .B1(_08737_),
    .B2(_08520_),
    .C1(_08739_),
    .C2(_08477_),
    .ZN(_08740_));
 NOR3_X4 _31214_ (.A1(_08394_),
    .A2(_08370_),
    .A3(_08399_),
    .ZN(_08741_));
 MUX2_X1 _31215_ (.A(_08669_),
    .B(_08741_),
    .S(_08514_),
    .Z(_08742_));
 NOR2_X1 _31216_ (.A1(_08443_),
    .A2(_08553_),
    .ZN(_08743_));
 AOI221_X2 _31217_ (.A(_08184_),
    .B1(_08230_),
    .B2(_08232_),
    .C1(_08195_),
    .C2(_07108_),
    .ZN(_08744_));
 OAI33_X1 _31218_ (.A1(_08270_),
    .A2(_08272_),
    .A3(_08574_),
    .B1(_08743_),
    .B2(_08744_),
    .B3(_08551_),
    .ZN(_08745_));
 NOR3_X2 _31219_ (.A1(_08282_),
    .A2(_08358_),
    .A3(_08516_),
    .ZN(_08746_));
 OAI22_X4 _31220_ (.A1(_08350_),
    .A2(_08368_),
    .B1(_08556_),
    .B2(_08380_),
    .ZN(_08747_));
 AOI222_X2 _31221_ (.A1(_08555_),
    .A2(_08742_),
    .B1(_08745_),
    .B2(_08746_),
    .C1(_08747_),
    .C2(_08663_),
    .ZN(_08748_));
 NAND2_X1 _31222_ (.A1(_08235_),
    .A2(_08362_),
    .ZN(_08749_));
 OR2_X1 _31223_ (.A1(_08484_),
    .A2(_08633_),
    .ZN(_08750_));
 MUX2_X1 _31224_ (.A(_08683_),
    .B(_08409_),
    .S(_08367_),
    .Z(_08751_));
 OAI211_X2 _31225_ (.A(_08362_),
    .B(_08384_),
    .C1(_08363_),
    .C2(_08388_),
    .ZN(_08752_));
 OAI33_X1 _31226_ (.A1(_08749_),
    .A2(_08750_),
    .A3(_08751_),
    .B1(_08752_),
    .B2(_08274_),
    .B3(_08257_),
    .ZN(_08753_));
 NAND3_X1 _31227_ (.A1(_08359_),
    .A2(_08564_),
    .A3(_08384_),
    .ZN(_08754_));
 AOI21_X1 _31228_ (.A(_08639_),
    .B1(_08523_),
    .B2(_08514_),
    .ZN(_08755_));
 AOI22_X2 _31229_ (.A1(_08282_),
    .A2(_08639_),
    .B1(_08498_),
    .B2(_08327_),
    .ZN(_08756_));
 OAI22_X2 _31230_ (.A1(_08754_),
    .A2(_08755_),
    .B1(_08756_),
    .B2(_08627_),
    .ZN(_08757_));
 NOR4_X1 _31231_ (.A1(_08402_),
    .A2(_08581_),
    .A3(_08545_),
    .A4(_08409_),
    .ZN(_08758_));
 MUX2_X1 _31232_ (.A(_08539_),
    .B(_08758_),
    .S(_08514_),
    .Z(_08759_));
 AOI211_X2 _31233_ (.A(_08753_),
    .B(_08757_),
    .C1(_08555_),
    .C2(_08759_),
    .ZN(_08760_));
 NAND4_X2 _31234_ (.A1(_08734_),
    .A2(_08740_),
    .A3(_08748_),
    .A4(_08760_),
    .ZN(_08761_));
 NOR2_X1 _31235_ (.A1(_08457_),
    .A2(_08699_),
    .ZN(_08762_));
 OAI33_X1 _31236_ (.A1(_08343_),
    .A2(_08551_),
    .A3(_08257_),
    .B1(_08511_),
    .B2(_08274_),
    .B3(_08498_),
    .ZN(_08763_));
 NAND4_X1 _31237_ (.A1(_08235_),
    .A2(_08362_),
    .A3(_08497_),
    .A4(_08363_),
    .ZN(_08764_));
 AOI21_X1 _31238_ (.A(_08291_),
    .B1(_08628_),
    .B2(_08764_),
    .ZN(_08765_));
 NAND3_X1 _31239_ (.A1(_08542_),
    .A2(_08251_),
    .A3(_08384_),
    .ZN(_08766_));
 NAND4_X1 _31240_ (.A1(_08381_),
    .A2(_08359_),
    .A3(_08553_),
    .A4(_08384_),
    .ZN(_08767_));
 AOI21_X1 _31241_ (.A(_08217_),
    .B1(_08766_),
    .B2(_08767_),
    .ZN(_08768_));
 NOR3_X1 _31242_ (.A1(_08763_),
    .A2(_08765_),
    .A3(_08768_),
    .ZN(_08769_));
 AND2_X1 _31243_ (.A1(_08683_),
    .A2(_08620_),
    .ZN(_08770_));
 NAND3_X1 _31244_ (.A1(_08357_),
    .A2(_08618_),
    .A3(_08523_),
    .ZN(_08771_));
 OAI22_X1 _31245_ (.A1(_08269_),
    .A2(_08588_),
    .B1(_08770_),
    .B2(_08771_),
    .ZN(_08772_));
 MUX2_X1 _31246_ (.A(_08561_),
    .B(_08217_),
    .S(_08564_),
    .Z(_08773_));
 NOR2_X1 _31247_ (.A1(_08556_),
    .A2(_08773_),
    .ZN(_08774_));
 OAI21_X1 _31248_ (.A(_08515_),
    .B1(_08772_),
    .B2(_08774_),
    .ZN(_08775_));
 NAND4_X2 _31249_ (.A1(_08532_),
    .A2(_08762_),
    .A3(_08769_),
    .A4(_08775_),
    .ZN(_08776_));
 NOR3_X1 _31250_ (.A1(_08281_),
    .A2(_08361_),
    .A3(_08334_),
    .ZN(_08777_));
 OAI21_X1 _31251_ (.A(_08292_),
    .B1(_08777_),
    .B2(_08490_),
    .ZN(_08778_));
 AOI21_X1 _31252_ (.A(_08283_),
    .B1(_08511_),
    .B2(_08711_),
    .ZN(_08779_));
 NOR2_X1 _31253_ (.A1(_08741_),
    .A2(_08779_),
    .ZN(_08780_));
 AOI22_X2 _31254_ (.A1(_08375_),
    .A2(_08335_),
    .B1(_08523_),
    .B2(_08435_),
    .ZN(_08781_));
 OAI221_X2 _31255_ (.A(_08778_),
    .B1(_08780_),
    .B2(_08306_),
    .C1(_08257_),
    .C2(_08781_),
    .ZN(_08782_));
 NOR2_X1 _31256_ (.A1(_08439_),
    .A2(_08441_),
    .ZN(_08783_));
 NOR2_X1 _31257_ (.A1(_08561_),
    .A2(_08511_),
    .ZN(_08784_));
 OAI221_X2 _31258_ (.A(_08283_),
    .B1(_08374_),
    .B2(_08783_),
    .C1(_08784_),
    .C2(_08555_),
    .ZN(_08785_));
 NOR2_X4 _31259_ (.A1(_08347_),
    .A2(_08502_),
    .ZN(_08786_));
 NOR3_X4 _31260_ (.A1(_08331_),
    .A2(_08421_),
    .A3(_08372_),
    .ZN(_08787_));
 AOI22_X4 _31261_ (.A1(_08786_),
    .A2(_08335_),
    .B1(_08787_),
    .B2(_08198_),
    .ZN(_08788_));
 NAND3_X1 _31262_ (.A1(_08663_),
    .A2(_08384_),
    .A3(_08363_),
    .ZN(_08789_));
 MUX2_X1 _31263_ (.A(_08443_),
    .B(_08358_),
    .S(_08485_),
    .Z(_08790_));
 OAI21_X1 _31264_ (.A(_08789_),
    .B1(_08790_),
    .B2(_08683_),
    .ZN(_08791_));
 NOR2_X1 _31265_ (.A1(_08545_),
    .A2(_08339_),
    .ZN(_08792_));
 NAND3_X1 _31266_ (.A1(_08342_),
    .A2(_08511_),
    .A3(_08582_),
    .ZN(_08793_));
 AOI22_X2 _31267_ (.A1(_08791_),
    .A2(_08792_),
    .B1(_08793_),
    .B2(_08619_),
    .ZN(_08794_));
 NAND2_X1 _31268_ (.A1(_08375_),
    .A2(_08498_),
    .ZN(_08795_));
 OAI22_X4 _31269_ (.A1(_08342_),
    .A2(_08795_),
    .B1(_08628_),
    .B2(_08520_),
    .ZN(_08796_));
 AOI21_X1 _31270_ (.A(_08467_),
    .B1(_08377_),
    .B2(_08386_),
    .ZN(_08797_));
 OAI21_X2 _31271_ (.A(_08487_),
    .B1(_08564_),
    .B2(_08797_),
    .ZN(_08798_));
 NAND4_X1 _31272_ (.A1(_08377_),
    .A2(_08362_),
    .A3(_08348_),
    .A4(_08363_),
    .ZN(_08799_));
 AOI221_X2 _31273_ (.A(_08491_),
    .B1(_08460_),
    .B2(_08469_),
    .C1(_08799_),
    .C2(_08467_),
    .ZN(_08800_));
 AOI22_X4 _31274_ (.A1(_08488_),
    .A2(_08796_),
    .B1(_08798_),
    .B2(_08800_),
    .ZN(_08801_));
 NAND4_X2 _31275_ (.A1(_08785_),
    .A2(_08788_),
    .A3(_08794_),
    .A4(_08801_),
    .ZN(_08802_));
 NOR4_X4 _31276_ (.A1(_08761_),
    .A2(_08776_),
    .A3(_08782_),
    .A4(_08802_),
    .ZN(_08803_));
 OR2_X2 _31277_ (.A1(_06706_),
    .A2(_08803_),
    .ZN(_08804_));
 XNOR2_X1 _31278_ (.A(_07274_),
    .B(_08187_),
    .ZN(_08805_));
 XNOR2_X1 _31279_ (.A(_00367_),
    .B(_08805_),
    .ZN(_08806_));
 XOR2_X1 _31280_ (.A(_07643_),
    .B(_07292_),
    .Z(_08807_));
 XNOR2_X1 _31281_ (.A(_08806_),
    .B(_08807_),
    .ZN(_08808_));
 BUF_X4 _31282_ (.A(_07231_),
    .Z(_08809_));
 MUX2_X2 _31283_ (.A(_07644_),
    .B(_08808_),
    .S(_08809_),
    .Z(_08810_));
 OAI221_X2 _31284_ (.A(_19384_),
    .B1(_07893_),
    .B2(_08810_),
    .C1(_07906_),
    .C2(\block_reg[0][18] ),
    .ZN(_08811_));
 NAND2_X1 _31285_ (.A1(_07908_),
    .A2(_08810_),
    .ZN(_08812_));
 INV_X1 _31286_ (.A(\block_reg[0][18] ),
    .ZN(_08813_));
 OAI21_X1 _31287_ (.A(_08812_),
    .B1(_07787_),
    .B2(_08813_),
    .ZN(_08814_));
 OR2_X1 _31288_ (.A1(_19384_),
    .A2(_08814_),
    .ZN(_08815_));
 AOI21_X2 _31289_ (.A(_06704_),
    .B1(_08811_),
    .B2(_08815_),
    .ZN(_08816_));
 AOI22_X1 _31290_ (.A1(_08730_),
    .A2(_07661_),
    .B1(_08804_),
    .B2(_08816_),
    .ZN(_00711_));
 XNOR2_X2 _31291_ (.A(_08491_),
    .B(_08484_),
    .ZN(_08817_));
 NOR2_X1 _31292_ (.A1(_08511_),
    .A2(_08817_),
    .ZN(_08818_));
 NOR2_X1 _31293_ (.A1(_08663_),
    .A2(_08510_),
    .ZN(_08819_));
 AOI21_X1 _31294_ (.A(_08818_),
    .B1(_08819_),
    .B2(_08492_),
    .ZN(_08820_));
 OAI221_X2 _31295_ (.A(_08487_),
    .B1(_08510_),
    .B2(_08633_),
    .C1(_08820_),
    .C2(_08515_),
    .ZN(_08821_));
 NOR3_X1 _31296_ (.A1(_08488_),
    .A2(_08663_),
    .A3(_08469_),
    .ZN(_08822_));
 AOI21_X1 _31297_ (.A(_08822_),
    .B1(_08374_),
    .B2(_08663_),
    .ZN(_08823_));
 AOI21_X1 _31298_ (.A(_08676_),
    .B1(_08374_),
    .B2(_08515_),
    .ZN(_08824_));
 AOI21_X1 _31299_ (.A(_08506_),
    .B1(_08435_),
    .B2(_08492_),
    .ZN(_08825_));
 OAI222_X2 _31300_ (.A1(_08283_),
    .A2(_08823_),
    .B1(_08824_),
    .B2(_08492_),
    .C1(_08257_),
    .C2(_08825_),
    .ZN(_08826_));
 OAI21_X4 _31301_ (.A(_08821_),
    .B1(_08826_),
    .B2(_08487_),
    .ZN(_08827_));
 NOR4_X4 _31302_ (.A1(_08553_),
    .A2(_08545_),
    .A3(_08370_),
    .A4(_08409_),
    .ZN(_08828_));
 AND2_X1 _31303_ (.A1(_08322_),
    .A2(_08828_),
    .ZN(_08829_));
 OAI21_X2 _31304_ (.A(_08515_),
    .B1(_08649_),
    .B2(_08829_),
    .ZN(_08830_));
 OAI21_X2 _31305_ (.A(_08679_),
    .B1(_08539_),
    .B2(_08676_),
    .ZN(_08831_));
 NOR2_X4 _31306_ (.A1(_08347_),
    .A2(_08405_),
    .ZN(_08832_));
 NAND2_X1 _31307_ (.A1(_08355_),
    .A2(_08394_),
    .ZN(_08833_));
 MUX2_X1 _31308_ (.A(_08374_),
    .B(_08428_),
    .S(_08833_),
    .Z(_08834_));
 AOI22_X4 _31309_ (.A1(_08447_),
    .A2(_08832_),
    .B1(_08834_),
    .B2(_08395_),
    .ZN(_08835_));
 NAND4_X4 _31310_ (.A1(_08733_),
    .A2(_08830_),
    .A3(_08831_),
    .A4(_08835_),
    .ZN(_08836_));
 NOR2_X1 _31311_ (.A1(_08486_),
    .A2(_08534_),
    .ZN(_08837_));
 AND2_X1 _31312_ (.A1(_08459_),
    .A2(_08534_),
    .ZN(_08838_));
 AOI22_X1 _31313_ (.A1(_08374_),
    .A2(_08837_),
    .B1(_08838_),
    .B2(_08335_),
    .ZN(_08839_));
 NOR2_X1 _31314_ (.A1(_08488_),
    .A2(_08839_),
    .ZN(_08840_));
 OAI33_X1 _31315_ (.A1(_08375_),
    .A2(_08556_),
    .A3(_08337_),
    .B1(_08393_),
    .B2(_08398_),
    .B3(_08553_),
    .ZN(_08841_));
 AND2_X1 _31316_ (.A1(_08492_),
    .A2(_08841_),
    .ZN(_08842_));
 NOR4_X1 _31317_ (.A1(_08542_),
    .A2(_08401_),
    .A3(_08516_),
    .A4(_08216_),
    .ZN(_08843_));
 NOR3_X1 _31318_ (.A1(_08459_),
    .A2(_08518_),
    .A3(_08519_),
    .ZN(_08844_));
 OAI21_X1 _31319_ (.A(_08564_),
    .B1(_08843_),
    .B2(_08844_),
    .ZN(_08845_));
 NOR2_X4 _31320_ (.A1(_08333_),
    .A2(_08423_),
    .ZN(_08846_));
 OAI221_X2 _31321_ (.A(_08846_),
    .B1(_08213_),
    .B2(_08206_),
    .C1(_08375_),
    .C2(_08542_),
    .ZN(_08847_));
 NOR2_X2 _31322_ (.A1(_08290_),
    .A2(_08256_),
    .ZN(_08848_));
 AOI222_X2 _31323_ (.A1(_08786_),
    .A2(_08671_),
    .B1(_08537_),
    .B2(_08848_),
    .C1(_08832_),
    .C2(_08731_),
    .ZN(_08849_));
 NOR3_X1 _31324_ (.A1(_08358_),
    .A2(_08551_),
    .A3(_08534_),
    .ZN(_08850_));
 NOR4_X1 _31325_ (.A1(_08281_),
    .A2(_08361_),
    .A3(_08291_),
    .A4(_08744_),
    .ZN(_08851_));
 OAI21_X1 _31326_ (.A(_08386_),
    .B1(_08850_),
    .B2(_08851_),
    .ZN(_08852_));
 NAND4_X1 _31327_ (.A1(_08845_),
    .A2(_08847_),
    .A3(_08849_),
    .A4(_08852_),
    .ZN(_08853_));
 AOI21_X1 _31328_ (.A(_08366_),
    .B1(_08355_),
    .B2(_08312_),
    .ZN(_08854_));
 AOI21_X1 _31329_ (.A(_08401_),
    .B1(_08418_),
    .B2(_08334_),
    .ZN(_08855_));
 AOI222_X2 _31330_ (.A1(_08505_),
    .A2(_08523_),
    .B1(_08672_),
    .B2(_08854_),
    .C1(_08855_),
    .C2(_08315_),
    .ZN(_08856_));
 OAI221_X1 _31331_ (.A(_08778_),
    .B1(_08856_),
    .B2(_08282_),
    .C1(_08257_),
    .C2(_08781_),
    .ZN(_08857_));
 OR4_X2 _31332_ (.A1(_08840_),
    .A2(_08842_),
    .A3(_08853_),
    .A4(_08857_),
    .ZN(_08858_));
 NAND3_X1 _31333_ (.A1(_08235_),
    .A2(_08359_),
    .A3(_08379_),
    .ZN(_08859_));
 AOI21_X1 _31334_ (.A(_08498_),
    .B1(_08378_),
    .B2(_08859_),
    .ZN(_08860_));
 OAI33_X1 _31335_ (.A1(_08381_),
    .A2(_08368_),
    .A3(_08216_),
    .B1(_08256_),
    .B2(_08303_),
    .B3(_08273_),
    .ZN(_08861_));
 OAI22_X1 _31336_ (.A1(_08450_),
    .A2(_08627_),
    .B1(_08698_),
    .B2(_08582_),
    .ZN(_08862_));
 OR3_X2 _31337_ (.A1(_08860_),
    .A2(_08861_),
    .A3(_08862_),
    .ZN(_08863_));
 NOR2_X2 _31338_ (.A1(_08551_),
    .A2(_08257_),
    .ZN(_08864_));
 AOI21_X1 _31339_ (.A(_08864_),
    .B1(_08557_),
    .B2(_08555_),
    .ZN(_08865_));
 NOR2_X1 _31340_ (.A1(_08627_),
    .A2(_08865_),
    .ZN(_08866_));
 NOR2_X1 _31341_ (.A1(_08274_),
    .A2(_08534_),
    .ZN(_08867_));
 AOI22_X2 _31342_ (.A1(_08619_),
    .A2(_08506_),
    .B1(_08867_),
    .B2(_08435_),
    .ZN(_08868_));
 AOI21_X1 _31343_ (.A(_08544_),
    .B1(_08672_),
    .B2(_08467_),
    .ZN(_08869_));
 OAI21_X1 _31344_ (.A(_08691_),
    .B1(_08587_),
    .B2(_08635_),
    .ZN(_08870_));
 OAI221_X1 _31345_ (.A(_08868_),
    .B1(_08869_),
    .B2(_08591_),
    .C1(_08491_),
    .C2(_08870_),
    .ZN(_08871_));
 OAI33_X1 _31346_ (.A1(_08402_),
    .A2(_08518_),
    .A3(_08216_),
    .B1(_08303_),
    .B2(_08551_),
    .B3(_08281_),
    .ZN(_08872_));
 AND2_X1 _31347_ (.A1(_08564_),
    .A2(_08872_),
    .ZN(_08873_));
 OR4_X2 _31348_ (.A1(_08863_),
    .A2(_08866_),
    .A3(_08871_),
    .A4(_08873_),
    .ZN(_08874_));
 AOI22_X1 _31349_ (.A1(_08543_),
    .A2(_08490_),
    .B1(_08506_),
    .B2(_08555_),
    .ZN(_08875_));
 AND2_X1 _31350_ (.A1(_08377_),
    .A2(_08390_),
    .ZN(_08876_));
 AND3_X1 _31351_ (.A1(_08402_),
    .A2(_08519_),
    .A3(_08391_),
    .ZN(_08877_));
 OAI221_X2 _31352_ (.A(_08324_),
    .B1(_08876_),
    .B2(_08877_),
    .C1(_08332_),
    .C2(_08297_),
    .ZN(_08878_));
 AND3_X1 _31353_ (.A1(_08485_),
    .A2(_08875_),
    .A3(_08878_),
    .ZN(_08879_));
 OAI22_X2 _31354_ (.A1(_08349_),
    .A2(_08517_),
    .B1(_08350_),
    .B2(_08661_),
    .ZN(_08880_));
 NOR2_X1 _31355_ (.A1(_08367_),
    .A2(_08516_),
    .ZN(_08881_));
 OAI22_X1 _31356_ (.A1(_08269_),
    .A2(_08217_),
    .B1(_08469_),
    .B2(_08367_),
    .ZN(_08882_));
 AOI221_X2 _31357_ (.A(_08484_),
    .B1(_08880_),
    .B2(_08881_),
    .C1(_08882_),
    .C2(_08514_),
    .ZN(_08883_));
 OAI211_X2 _31358_ (.A(_08559_),
    .B(_08630_),
    .C1(_08879_),
    .C2(_08883_),
    .ZN(_08884_));
 NOR4_X4 _31359_ (.A1(_08836_),
    .A2(_08858_),
    .A3(_08874_),
    .A4(_08884_),
    .ZN(_08885_));
 AND2_X2 _31360_ (.A1(_08827_),
    .A2(_08885_),
    .ZN(_08886_));
 OR2_X2 _31361_ (.A1(_06706_),
    .A2(_08886_),
    .ZN(_08887_));
 CLKBUF_X3 _31362_ (.A(_07904_),
    .Z(_08888_));
 CLKBUF_X3 _31363_ (.A(_07253_),
    .Z(_08889_));
 XNOR2_X1 _31364_ (.A(_07283_),
    .B(_08165_),
    .ZN(_08890_));
 XNOR2_X1 _31365_ (.A(_07338_),
    .B(_08890_),
    .ZN(_08891_));
 XOR2_X2 _31366_ (.A(_00370_),
    .B(_07644_),
    .Z(_08892_));
 XOR2_X2 _31367_ (.A(_00347_),
    .B(_07274_),
    .Z(_08893_));
 XNOR2_X1 _31368_ (.A(_08892_),
    .B(_08893_),
    .ZN(_08894_));
 XNOR2_X1 _31369_ (.A(_08891_),
    .B(_08894_),
    .ZN(_08895_));
 BUF_X4 _31370_ (.A(_07231_),
    .Z(_08896_));
 MUX2_X1 _31371_ (.A(_07794_),
    .B(_08895_),
    .S(_08896_),
    .Z(_08897_));
 OAI22_X1 _31372_ (.A1(\block_reg[0][19] ),
    .A2(_08888_),
    .B1(_08889_),
    .B2(_08897_),
    .ZN(_08898_));
 NOR2_X1 _31373_ (.A1(_03286_),
    .A2(_08898_),
    .ZN(_08899_));
 BUF_X4 _31374_ (.A(_07805_),
    .Z(_08900_));
 CLKBUF_X3 _31375_ (.A(_07228_),
    .Z(_08901_));
 AOI22_X1 _31376_ (.A1(\block_reg[0][19] ),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_08897_),
    .ZN(_08902_));
 AND2_X1 _31377_ (.A1(_03286_),
    .A2(_08902_),
    .ZN(_08903_));
 OAI21_X1 _31378_ (.A(_08887_),
    .B1(_08899_),
    .B2(_08903_),
    .ZN(_08904_));
 BUF_X2 _31379_ (.A(\core.enc_block.block_w0_reg[19] ),
    .Z(_08905_));
 BUF_X4 _31380_ (.A(_06703_),
    .Z(_08906_));
 MUX2_X1 _31381_ (.A(_08904_),
    .B(_08905_),
    .S(_08906_),
    .Z(_00712_));
 OR4_X4 _31382_ (.A1(_06918_),
    .A2(_06994_),
    .A3(_07010_),
    .A4(_07043_),
    .ZN(_08907_));
 NOR2_X4 _31383_ (.A1(_06921_),
    .A2(_06968_),
    .ZN(_08908_));
 AOI21_X1 _31384_ (.A(_07070_),
    .B1(_07078_),
    .B2(_07098_),
    .ZN(_08909_));
 AOI22_X2 _31385_ (.A1(_06991_),
    .A2(_07082_),
    .B1(_08908_),
    .B2(_08909_),
    .ZN(_08910_));
 BUF_X4 _31386_ (.A(_06855_),
    .Z(_08911_));
 OAI221_X1 _31387_ (.A(_07074_),
    .B1(_07052_),
    .B2(_06876_),
    .C1(_08911_),
    .C2(_07077_),
    .ZN(_08912_));
 OAI21_X1 _31388_ (.A(_08912_),
    .B1(_06906_),
    .B2(_07074_),
    .ZN(_08913_));
 OAI33_X1 _31389_ (.A1(_06855_),
    .A2(_06872_),
    .A3(_06856_),
    .B1(_06909_),
    .B2(_07025_),
    .B3(_07035_),
    .ZN(_08914_));
 AOI221_X2 _31390_ (.A(_07135_),
    .B1(_08914_),
    .B2(_06808_),
    .C1(_07020_),
    .C2(_07159_),
    .ZN(_08915_));
 OAI221_X2 _31391_ (.A(_08910_),
    .B1(_08913_),
    .B2(_07028_),
    .C1(_08915_),
    .C2(_07102_),
    .ZN(_08916_));
 INV_X1 _31392_ (.A(_08916_),
    .ZN(_08917_));
 AOI21_X1 _31393_ (.A(_07106_),
    .B1(_07146_),
    .B2(_06847_),
    .ZN(_08918_));
 AOI221_X1 _31394_ (.A(_06853_),
    .B1(_06827_),
    .B2(_06833_),
    .C1(_06847_),
    .C2(_07055_),
    .ZN(_08919_));
 NOR3_X1 _31395_ (.A1(_07060_),
    .A2(_08918_),
    .A3(_08919_),
    .ZN(_08920_));
 NOR2_X1 _31396_ (.A1(_06816_),
    .A2(_07125_),
    .ZN(_08921_));
 MUX2_X1 _31397_ (.A(_06981_),
    .B(_07211_),
    .S(_06880_),
    .Z(_08922_));
 NOR2_X2 _31398_ (.A1(_06921_),
    .A2(_06944_),
    .ZN(_08923_));
 NAND4_X1 _31399_ (.A1(_06971_),
    .A2(_08921_),
    .A3(_08922_),
    .A4(_08923_),
    .ZN(_08924_));
 NAND2_X1 _31400_ (.A1(_07122_),
    .A2(_07130_),
    .ZN(_08925_));
 NOR2_X4 _31401_ (.A1(_06898_),
    .A2(_06808_),
    .ZN(_08926_));
 NOR3_X4 _31402_ (.A1(_06815_),
    .A2(_06759_),
    .A3(_06872_),
    .ZN(_08927_));
 AOI22_X1 _31403_ (.A1(_08926_),
    .A2(_07023_),
    .B1(_08927_),
    .B2(_06964_),
    .ZN(_08928_));
 OAI221_X1 _31404_ (.A(_08924_),
    .B1(_07186_),
    .B2(_08925_),
    .C1(_07067_),
    .C2(_08928_),
    .ZN(_08929_));
 NAND2_X1 _31405_ (.A1(_07138_),
    .A2(_07172_),
    .ZN(_08930_));
 AOI21_X1 _31406_ (.A(_06877_),
    .B1(_06928_),
    .B2(_07057_),
    .ZN(_08931_));
 OAI22_X2 _31407_ (.A1(_06874_),
    .A2(_07028_),
    .B1(_07088_),
    .B2(_06921_),
    .ZN(_08932_));
 AOI222_X2 _31408_ (.A1(_06945_),
    .A2(_07146_),
    .B1(_07178_),
    .B2(_08931_),
    .C1(_08932_),
    .C2(_07005_),
    .ZN(_08933_));
 NOR3_X2 _31409_ (.A1(_06730_),
    .A2(_06932_),
    .A3(_07052_),
    .ZN(_08934_));
 NOR2_X1 _31410_ (.A1(_06891_),
    .A2(_06955_),
    .ZN(_08935_));
 AOI222_X2 _31411_ (.A1(_06973_),
    .A2(_07048_),
    .B1(_08934_),
    .B2(_08935_),
    .C1(_08908_),
    .C2(_06989_),
    .ZN(_08936_));
 NAND4_X1 _31412_ (.A1(_07150_),
    .A2(_08930_),
    .A3(_08933_),
    .A4(_08936_),
    .ZN(_08937_));
 OAI221_X2 _31413_ (.A(_06924_),
    .B1(_06728_),
    .B2(_06712_),
    .C1(_06859_),
    .C2(_06888_),
    .ZN(_08938_));
 OAI221_X2 _31414_ (.A(_06953_),
    .B1(_06832_),
    .B2(_06830_),
    .C1(_06796_),
    .C2(_06887_),
    .ZN(_08939_));
 AOI21_X1 _31415_ (.A(_08938_),
    .B1(_07017_),
    .B2(_08939_),
    .ZN(_08940_));
 OAI21_X2 _31416_ (.A(_06991_),
    .B1(_07030_),
    .B2(_08940_),
    .ZN(_08941_));
 NOR2_X4 _31417_ (.A1(_07028_),
    .A2(_07093_),
    .ZN(_08942_));
 BUF_X4 _31418_ (.A(_06839_),
    .Z(_08943_));
 AOI22_X2 _31419_ (.A1(_07178_),
    .A2(_08908_),
    .B1(_08942_),
    .B2(_08943_),
    .ZN(_08944_));
 NAND4_X2 _31420_ (.A1(_07194_),
    .A2(_07197_),
    .A3(_08941_),
    .A4(_08944_),
    .ZN(_08945_));
 OR4_X2 _31421_ (.A1(_08920_),
    .A2(_08929_),
    .A3(_08937_),
    .A4(_08945_),
    .ZN(_08946_));
 NOR3_X1 _31422_ (.A1(_07066_),
    .A2(_07097_),
    .A3(_07140_),
    .ZN(_08947_));
 OAI221_X2 _31423_ (.A(_07074_),
    .B1(_08947_),
    .B2(_06829_),
    .C1(_06832_),
    .C2(_06830_),
    .ZN(_08948_));
 NOR4_X1 _31424_ (.A1(_07057_),
    .A2(_07090_),
    .A3(_07119_),
    .A4(_07140_),
    .ZN(_08949_));
 NOR4_X2 _31425_ (.A1(_06900_),
    .A2(_07104_),
    .A3(_08911_),
    .A4(_07090_),
    .ZN(_08950_));
 OAI21_X2 _31426_ (.A(_07076_),
    .B1(_08949_),
    .B2(_08950_),
    .ZN(_08951_));
 AOI21_X4 _31427_ (.A(_07079_),
    .B1(_07077_),
    .B2(_07090_),
    .ZN(_08952_));
 NOR3_X1 _31428_ (.A1(_08911_),
    .A2(_07098_),
    .A3(_07119_),
    .ZN(_08953_));
 OAI21_X2 _31429_ (.A(_07195_),
    .B1(_08952_),
    .B2(_08953_),
    .ZN(_08954_));
 NAND4_X4 _31430_ (.A1(_07160_),
    .A2(_08948_),
    .A3(_08951_),
    .A4(_08954_),
    .ZN(_08955_));
 NOR3_X2 _31431_ (.A1(_06894_),
    .A2(_06876_),
    .A3(_07140_),
    .ZN(_08956_));
 AOI22_X1 _31432_ (.A1(_07112_),
    .A2(_07138_),
    .B1(_07020_),
    .B2(_08956_),
    .ZN(_08957_));
 NOR2_X1 _31433_ (.A1(_07069_),
    .A2(_08957_),
    .ZN(_08958_));
 NAND2_X1 _31434_ (.A1(_07144_),
    .A2(_07155_),
    .ZN(_08959_));
 OAI22_X2 _31435_ (.A1(_07090_),
    .A2(_07092_),
    .B1(_07079_),
    .B2(_07087_),
    .ZN(_08960_));
 AOI21_X2 _31436_ (.A(_07055_),
    .B1(_08960_),
    .B2(_07061_),
    .ZN(_08961_));
 NOR3_X4 _31437_ (.A1(_06922_),
    .A2(_07140_),
    .A3(_06885_),
    .ZN(_08962_));
 NOR2_X1 _31438_ (.A1(_07059_),
    .A2(_08962_),
    .ZN(_08963_));
 AOI221_X2 _31439_ (.A(_07119_),
    .B1(_06950_),
    .B2(_06905_),
    .C1(_07159_),
    .C2(_07168_),
    .ZN(_08964_));
 OAI22_X2 _31440_ (.A1(_08959_),
    .A2(_08961_),
    .B1(_08963_),
    .B2(_08964_),
    .ZN(_08965_));
 OR4_X2 _31441_ (.A1(_07029_),
    .A2(_08955_),
    .A3(_08958_),
    .A4(_08965_),
    .ZN(_08966_));
 OAI33_X1 _31442_ (.A1(_07063_),
    .A2(_07099_),
    .A3(_07046_),
    .B1(_07053_),
    .B2(_07120_),
    .B3(_07050_),
    .ZN(_08967_));
 NAND2_X2 _31443_ (.A1(_07057_),
    .A2(_07104_),
    .ZN(_08968_));
 NOR2_X1 _31444_ (.A1(_07165_),
    .A2(_07074_),
    .ZN(_08969_));
 NAND2_X1 _31445_ (.A1(_07129_),
    .A2(_07122_),
    .ZN(_08970_));
 OAI33_X1 _31446_ (.A1(_07060_),
    .A2(_07204_),
    .A3(_08968_),
    .B1(_08969_),
    .B2(_08970_),
    .B3(_07086_),
    .ZN(_08971_));
 AOI22_X4 _31447_ (.A1(_07155_),
    .A2(_08967_),
    .B1(_08971_),
    .B2(_07067_),
    .ZN(_08972_));
 NOR3_X2 _31448_ (.A1(_06899_),
    .A2(_06876_),
    .A3(_07091_),
    .ZN(_08973_));
 NOR3_X1 _31449_ (.A1(_07057_),
    .A2(_07077_),
    .A3(_07070_),
    .ZN(_08974_));
 OAI221_X1 _31450_ (.A(_07088_),
    .B1(_08973_),
    .B2(_08974_),
    .C1(_06728_),
    .C2(_06712_),
    .ZN(_08975_));
 AOI22_X1 _31451_ (.A1(_07045_),
    .A2(_07172_),
    .B1(_07156_),
    .B2(_07155_),
    .ZN(_08976_));
 NOR2_X1 _31452_ (.A1(_07098_),
    .A2(_07102_),
    .ZN(_08977_));
 OAI221_X2 _31453_ (.A(_06812_),
    .B1(_06860_),
    .B2(_06870_),
    .C1(_06888_),
    .C2(_06776_),
    .ZN(_08978_));
 OAI22_X1 _31454_ (.A1(_07080_),
    .A2(_07046_),
    .B1(_08978_),
    .B2(_07061_),
    .ZN(_08979_));
 AOI221_X2 _31455_ (.A(_07131_),
    .B1(_07119_),
    .B2(_06971_),
    .C1(_06953_),
    .C2(_06799_),
    .ZN(_08980_));
 OAI21_X1 _31456_ (.A(_08977_),
    .B1(_08979_),
    .B2(_08980_),
    .ZN(_08981_));
 NOR4_X1 _31457_ (.A1(_07057_),
    .A2(_07105_),
    .A3(_08911_),
    .A4(_07090_),
    .ZN(_08982_));
 NOR3_X1 _31458_ (.A1(_07068_),
    .A2(_07107_),
    .A3(_07053_),
    .ZN(_08983_));
 OAI21_X1 _31459_ (.A(_07110_),
    .B1(_08982_),
    .B2(_08983_),
    .ZN(_08984_));
 AND4_X2 _31460_ (.A1(_08975_),
    .A2(_08976_),
    .A3(_08981_),
    .A4(_08984_),
    .ZN(_08985_));
 OAI21_X1 _31461_ (.A(_06829_),
    .B1(_07165_),
    .B2(_07069_),
    .ZN(_08986_));
 NOR3_X1 _31462_ (.A1(_07107_),
    .A2(_07046_),
    .A3(_07053_),
    .ZN(_08987_));
 OAI21_X1 _31463_ (.A(_07069_),
    .B1(_07054_),
    .B2(_08987_),
    .ZN(_08988_));
 NAND4_X2 _31464_ (.A1(_06787_),
    .A2(_06845_),
    .A3(_06799_),
    .A4(_06953_),
    .ZN(_08989_));
 OAI33_X1 _31465_ (.A1(_07063_),
    .A2(_07078_),
    .A3(_08989_),
    .B1(_07017_),
    .B2(_07053_),
    .B3(_07087_),
    .ZN(_08990_));
 NOR3_X1 _31466_ (.A1(_06853_),
    .A2(_07097_),
    .A3(_07052_),
    .ZN(_08991_));
 OAI21_X1 _31467_ (.A(_07060_),
    .B1(_08990_),
    .B2(_08991_),
    .ZN(_08992_));
 AND3_X1 _31468_ (.A1(_08986_),
    .A2(_08988_),
    .A3(_08992_),
    .ZN(_08993_));
 OAI211_X4 _31469_ (.A(_08972_),
    .B(_08985_),
    .C1(_08993_),
    .C2(_07085_),
    .ZN(_08994_));
 NOR3_X2 _31470_ (.A1(_08946_),
    .A2(_08966_),
    .A3(_08994_),
    .ZN(_08995_));
 NAND3_X4 _31471_ (.A1(_08907_),
    .A2(_08917_),
    .A3(_08995_),
    .ZN(_08996_));
 NAND2_X2 _31472_ (.A1(_07260_),
    .A2(_08996_),
    .ZN(_08997_));
 XOR2_X2 _31473_ (.A(\core.enc_block.block_w3_reg[0] ),
    .B(_07791_),
    .Z(_08998_));
 BUF_X2 _31474_ (.A(\core.enc_block.block_w0_reg[25] ),
    .Z(_08999_));
 XOR2_X1 _31475_ (.A(_08187_),
    .B(_08999_),
    .Z(_09000_));
 XNOR2_X1 _31476_ (.A(_08998_),
    .B(_09000_),
    .ZN(_09001_));
 XNOR2_X1 _31477_ (.A(_00312_),
    .B(_07236_),
    .ZN(_09002_));
 XNOR2_X1 _31478_ (.A(_09001_),
    .B(_09002_),
    .ZN(_09003_));
 MUX2_X1 _31479_ (.A(_00364_),
    .B(_09003_),
    .S(_07242_),
    .Z(_09004_));
 BUF_X4 _31480_ (.A(_07805_),
    .Z(_09005_));
 AOI221_X2 _31481_ (.A(_03509_),
    .B1(_07808_),
    .B2(_09004_),
    .C1(_09005_),
    .C2(_06504_),
    .ZN(_09006_));
 CLKBUF_X3 _31482_ (.A(_07252_),
    .Z(_09007_));
 NOR2_X1 _31483_ (.A1(_09007_),
    .A2(_09004_),
    .ZN(_09008_));
 AOI21_X1 _31484_ (.A(_09008_),
    .B1(_08900_),
    .B2(\block_reg[0][1] ),
    .ZN(_09009_));
 AND2_X1 _31485_ (.A1(_03509_),
    .A2(_09009_),
    .ZN(_09010_));
 OAI21_X2 _31486_ (.A(_08997_),
    .B1(_09006_),
    .B2(_09010_),
    .ZN(_09011_));
 MUX2_X1 _31487_ (.A(_09011_),
    .B(\core.enc_block.block_w0_reg[1] ),
    .S(_08906_),
    .Z(_00713_));
 BUF_X2 _31488_ (.A(\core.enc_block.block_w0_reg[20] ),
    .Z(_09012_));
 INV_X1 _31489_ (.A(_09012_),
    .ZN(_09013_));
 NOR4_X2 _31490_ (.A1(_08502_),
    .A2(_08423_),
    .A3(_08291_),
    .A4(_08399_),
    .ZN(_09014_));
 AOI221_X2 _31491_ (.A(_09014_),
    .B1(_08832_),
    .B2(_08435_),
    .C1(_08671_),
    .C2(_08434_),
    .ZN(_09015_));
 AOI21_X2 _31492_ (.A(_08552_),
    .B1(_08555_),
    .B2(_08503_),
    .ZN(_09016_));
 AND2_X1 _31493_ (.A1(_08581_),
    .A2(_08395_),
    .ZN(_09017_));
 AOI22_X2 _31494_ (.A1(_08731_),
    .A2(_08198_),
    .B1(_09017_),
    .B2(_08429_),
    .ZN(_09018_));
 OAI221_X2 _31495_ (.A(_09015_),
    .B1(_09016_),
    .B2(_08305_),
    .C1(_08488_),
    .C2(_09018_),
    .ZN(_09019_));
 AND2_X1 _31496_ (.A1(_08492_),
    .A2(_08777_),
    .ZN(_09020_));
 AOI221_X2 _31497_ (.A(_08491_),
    .B1(_08360_),
    .B2(_08364_),
    .C1(_08230_),
    .C2(_08232_),
    .ZN(_09021_));
 OAI21_X2 _31498_ (.A(_08520_),
    .B1(_09020_),
    .B2(_09021_),
    .ZN(_09022_));
 MUX2_X1 _31499_ (.A(_08335_),
    .B(_08672_),
    .S(_08553_),
    .Z(_09023_));
 OAI22_X1 _31500_ (.A1(_08556_),
    .A2(_08339_),
    .B1(_08303_),
    .B2(_08561_),
    .ZN(_09024_));
 AOI222_X2 _31501_ (.A1(_08198_),
    .A2(_08593_),
    .B1(_09023_),
    .B2(_08427_),
    .C1(_09024_),
    .C2(_08503_),
    .ZN(_09025_));
 NAND4_X4 _31502_ (.A1(_08584_),
    .A2(net14),
    .A3(_09022_),
    .A4(_09025_),
    .ZN(_09026_));
 OR3_X4 _31503_ (.A1(_08836_),
    .A2(_09019_),
    .A3(_09026_),
    .ZN(_09027_));
 NAND2_X1 _31504_ (.A1(_08555_),
    .A2(_08742_),
    .ZN(_09028_));
 AOI22_X2 _31505_ (.A1(_08745_),
    .A2(_08746_),
    .B1(_08747_),
    .B2(_08663_),
    .ZN(_09029_));
 NAND2_X2 _31506_ (.A1(_09028_),
    .A2(_09029_),
    .ZN(_09030_));
 MUX2_X1 _31507_ (.A(_08414_),
    .B(_08412_),
    .S(_08443_),
    .Z(_09031_));
 NOR4_X1 _31508_ (.A1(_08361_),
    .A2(_08683_),
    .A3(_08535_),
    .A4(_09031_),
    .ZN(_09032_));
 OAI221_X1 _31509_ (.A(_08337_),
    .B1(_08373_),
    .B2(_08447_),
    .C1(_08327_),
    .C2(_08322_),
    .ZN(_09033_));
 MUX2_X1 _31510_ (.A(_08388_),
    .B(_08302_),
    .S(_08354_),
    .Z(_09034_));
 NOR3_X1 _31511_ (.A1(_08381_),
    .A2(_08401_),
    .A3(_08412_),
    .ZN(_09035_));
 NAND3_X1 _31512_ (.A1(_08477_),
    .A2(_09034_),
    .A3(_09035_),
    .ZN(_09036_));
 NAND2_X1 _31513_ (.A1(_09033_),
    .A2(_09036_),
    .ZN(_09037_));
 OR4_X2 _31514_ (.A1(_08479_),
    .A2(_08480_),
    .A3(_09032_),
    .A4(_09037_),
    .ZN(_09038_));
 AOI222_X2 _31515_ (.A1(_08676_),
    .A2(_08832_),
    .B1(_08846_),
    .B2(_08864_),
    .C1(_08506_),
    .C2(_08639_),
    .ZN(_09039_));
 NOR2_X1 _31516_ (.A1(_08198_),
    .A2(_08469_),
    .ZN(_09040_));
 OAI21_X1 _31517_ (.A(_08639_),
    .B1(_08539_),
    .B2(_09040_),
    .ZN(_09041_));
 OAI21_X1 _31518_ (.A(_08641_),
    .B1(_08540_),
    .B2(_08731_),
    .ZN(_09042_));
 OAI22_X1 _31519_ (.A1(_08402_),
    .A2(_08414_),
    .B1(_08545_),
    .B2(_08423_),
    .ZN(_09043_));
 NAND3_X1 _31520_ (.A1(_08786_),
    .A2(_08363_),
    .A3(_09043_),
    .ZN(_09044_));
 OAI21_X1 _31521_ (.A(_08619_),
    .B1(_08540_),
    .B2(_08505_),
    .ZN(_09045_));
 OAI21_X1 _31522_ (.A(_08335_),
    .B1(_08665_),
    .B2(_08619_),
    .ZN(_09046_));
 AND4_X1 _31523_ (.A1(_09042_),
    .A2(_09044_),
    .A3(_09045_),
    .A4(_09046_),
    .ZN(_09047_));
 NAND3_X2 _31524_ (.A1(_09039_),
    .A2(_09041_),
    .A3(_09047_),
    .ZN(_09048_));
 NAND3_X1 _31525_ (.A1(_08459_),
    .A2(_08581_),
    .A3(_08537_),
    .ZN(_09049_));
 NAND2_X1 _31526_ (.A1(_08635_),
    .A2(_08846_),
    .ZN(_09050_));
 AOI21_X1 _31527_ (.A(_08633_),
    .B1(_09049_),
    .B2(_09050_),
    .ZN(_09051_));
 NAND2_X1 _31528_ (.A1(_08553_),
    .A2(_08537_),
    .ZN(_09052_));
 OAI21_X1 _31529_ (.A(_08281_),
    .B1(_08537_),
    .B2(_08846_),
    .ZN(_09053_));
 AOI21_X1 _31530_ (.A(_08291_),
    .B1(_09052_),
    .B2(_09053_),
    .ZN(_09054_));
 NOR3_X1 _31531_ (.A1(_08291_),
    .A2(_08469_),
    .A3(_08313_),
    .ZN(_09055_));
 OAI33_X1 _31532_ (.A1(_08216_),
    .A2(_08556_),
    .A3(_08256_),
    .B1(_08627_),
    .B2(_08273_),
    .B3(_08197_),
    .ZN(_09056_));
 OR4_X2 _31533_ (.A1(_09051_),
    .A2(_09054_),
    .A3(_09055_),
    .A4(_09056_),
    .ZN(_09057_));
 OR4_X4 _31534_ (.A1(_09030_),
    .A2(_09038_),
    .A3(_09048_),
    .A4(_09057_),
    .ZN(_09058_));
 OAI21_X4 _31535_ (.A(_07260_),
    .B1(_09027_),
    .B2(_09058_),
    .ZN(_09059_));
 XNOR2_X1 _31536_ (.A(_07317_),
    .B(_07794_),
    .ZN(_09060_));
 XNOR2_X1 _31537_ (.A(_00330_),
    .B(_00350_),
    .ZN(_09061_));
 XNOR2_X1 _31538_ (.A(_09060_),
    .B(_09061_),
    .ZN(_09062_));
 XNOR2_X1 _31539_ (.A(_08891_),
    .B(_09062_),
    .ZN(_09063_));
 MUX2_X1 _31540_ (.A(_07895_),
    .B(_09063_),
    .S(_07243_),
    .Z(_09064_));
 OAI221_X2 _31541_ (.A(_03723_),
    .B1(_07893_),
    .B2(_09064_),
    .C1(_07906_),
    .C2(\block_reg[0][20] ),
    .ZN(_09065_));
 AOI22_X1 _31542_ (.A1(\block_reg[0][20] ),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_09064_),
    .ZN(_09066_));
 OAI21_X1 _31543_ (.A(_09066_),
    .B1(_03722_),
    .B2(_03721_),
    .ZN(_09067_));
 AOI21_X2 _31544_ (.A(_06704_),
    .B1(_09065_),
    .B2(_09067_),
    .ZN(_09068_));
 AOI22_X1 _31545_ (.A1(_09013_),
    .A2(_07661_),
    .B1(_09059_),
    .B2(_09068_),
    .ZN(_00714_));
 NOR2_X1 _31546_ (.A1(_08520_),
    .A2(_08429_),
    .ZN(_09069_));
 NOR3_X1 _31547_ (.A1(_08486_),
    .A2(_08490_),
    .A3(_08435_),
    .ZN(_09070_));
 NOR3_X1 _31548_ (.A1(_08750_),
    .A2(_09069_),
    .A3(_09070_),
    .ZN(_09071_));
 NOR2_X1 _31549_ (.A1(_08358_),
    .A2(_08400_),
    .ZN(_09072_));
 NOR2_X1 _31550_ (.A1(_08282_),
    .A2(_08491_),
    .ZN(_09073_));
 AOI21_X1 _31551_ (.A(_09073_),
    .B1(_08743_),
    .B2(_08573_),
    .ZN(_09074_));
 OAI22_X1 _31552_ (.A1(_08357_),
    .A2(_08633_),
    .B1(_09074_),
    .B2(_08520_),
    .ZN(_09075_));
 AOI21_X1 _31553_ (.A(_09071_),
    .B1(_09072_),
    .B2(_09075_),
    .ZN(_09076_));
 NOR3_X2 _31554_ (.A1(_08516_),
    .A2(_08517_),
    .A3(_08347_),
    .ZN(_09077_));
 NAND2_X1 _31555_ (.A1(_08663_),
    .A2(_09077_),
    .ZN(_09078_));
 NOR2_X1 _31556_ (.A1(_08581_),
    .A2(_08217_),
    .ZN(_09079_));
 OAI21_X1 _31557_ (.A(_09079_),
    .B1(_08428_),
    .B2(_08676_),
    .ZN(_09080_));
 AOI21_X1 _31558_ (.A(_08515_),
    .B1(_09078_),
    .B2(_09080_),
    .ZN(_09081_));
 NOR3_X1 _31559_ (.A1(_08471_),
    .A2(_08475_),
    .A3(_09081_),
    .ZN(_09082_));
 AOI21_X1 _31560_ (.A(_08577_),
    .B1(_08523_),
    .B2(_08428_),
    .ZN(_09083_));
 NOR3_X1 _31561_ (.A1(_08676_),
    .A2(_08428_),
    .A3(_08335_),
    .ZN(_09084_));
 NAND2_X1 _31562_ (.A1(_08639_),
    .A2(_08337_),
    .ZN(_09085_));
 OAI22_X2 _31563_ (.A1(_08503_),
    .A2(_09083_),
    .B1(_09084_),
    .B2(_09085_),
    .ZN(_09086_));
 OAI21_X1 _31564_ (.A(_08641_),
    .B1(_08846_),
    .B2(_08828_),
    .ZN(_09087_));
 NAND2_X1 _31565_ (.A1(_08868_),
    .A2(_09087_),
    .ZN(_09088_));
 NOR3_X2 _31566_ (.A1(_08513_),
    .A2(_09086_),
    .A3(_09088_),
    .ZN(_09089_));
 NOR3_X1 _31567_ (.A1(_08342_),
    .A2(_08564_),
    .A3(_08339_),
    .ZN(_09090_));
 AOI21_X1 _31568_ (.A(_08252_),
    .B1(_08339_),
    .B2(_08217_),
    .ZN(_09091_));
 AOI21_X1 _31569_ (.A(_09090_),
    .B1(_09091_),
    .B2(_08663_),
    .ZN(_09092_));
 NOR3_X2 _31570_ (.A1(_08418_),
    .A2(_08423_),
    .A3(_08216_),
    .ZN(_09093_));
 NOR3_X1 _31571_ (.A1(_08484_),
    .A2(_08306_),
    .A3(_08305_),
    .ZN(_09094_));
 OAI21_X1 _31572_ (.A(_08283_),
    .B1(_09093_),
    .B2(_09094_),
    .ZN(_09095_));
 AOI21_X1 _31573_ (.A(_08561_),
    .B1(_08276_),
    .B2(_08342_),
    .ZN(_09096_));
 OAI21_X1 _31574_ (.A(_08313_),
    .B1(_08649_),
    .B2(_09096_),
    .ZN(_09097_));
 AND3_X1 _31575_ (.A1(_09092_),
    .A2(_09095_),
    .A3(_09097_),
    .ZN(_09098_));
 NAND4_X2 _31576_ (.A1(_09076_),
    .A2(_09082_),
    .A3(_09089_),
    .A4(_09098_),
    .ZN(_09099_));
 OR3_X1 _31577_ (.A1(_08763_),
    .A2(_08765_),
    .A3(_08768_),
    .ZN(_09100_));
 MUX2_X1 _31578_ (.A(_08556_),
    .B(_08276_),
    .S(_08557_),
    .Z(_09101_));
 AOI21_X2 _31579_ (.A(_09093_),
    .B1(_08846_),
    .B2(_08523_),
    .ZN(_09102_));
 OAI22_X4 _31580_ (.A1(_08561_),
    .A2(_09101_),
    .B1(_09102_),
    .B2(_08503_),
    .ZN(_09103_));
 AOI22_X2 _31581_ (.A1(_08639_),
    .A2(_08671_),
    .B1(_08641_),
    .B2(_08540_),
    .ZN(_09104_));
 OAI222_X2 _31582_ (.A1(_08342_),
    .A2(_08440_),
    .B1(_08627_),
    .B2(_08338_),
    .C1(_09104_),
    .C2(_08581_),
    .ZN(_09105_));
 NAND2_X1 _31583_ (.A1(_08683_),
    .A2(_08400_),
    .ZN(_09106_));
 NOR4_X1 _31584_ (.A1(_08551_),
    .A2(_08502_),
    .A3(_08370_),
    .A4(_08666_),
    .ZN(_09107_));
 AOI22_X1 _31585_ (.A1(_08198_),
    .A2(_09077_),
    .B1(_09106_),
    .B2(_09107_),
    .ZN(_09108_));
 NOR3_X1 _31586_ (.A1(_08350_),
    .A2(_08661_),
    .A3(_08400_),
    .ZN(_09109_));
 NOR4_X1 _31587_ (.A1(_08516_),
    .A2(_08394_),
    .A3(_08349_),
    .A4(_08423_),
    .ZN(_09110_));
 OAI21_X1 _31588_ (.A(_08375_),
    .B1(_09109_),
    .B2(_09110_),
    .ZN(_09111_));
 NOR2_X1 _31589_ (.A1(_08381_),
    .A2(_08491_),
    .ZN(_09112_));
 AOI22_X2 _31590_ (.A1(_08540_),
    .A2(_08674_),
    .B1(_08741_),
    .B2(_09112_),
    .ZN(_09113_));
 OAI33_X1 _31591_ (.A1(_08297_),
    .A2(_08661_),
    .A3(_08300_),
    .B1(_08621_),
    .B2(_08394_),
    .B3(_08443_),
    .ZN(_09114_));
 NAND3_X1 _31592_ (.A1(_08618_),
    .A2(_08641_),
    .A3(_09114_),
    .ZN(_09115_));
 NAND4_X1 _31593_ (.A1(_09108_),
    .A2(_09111_),
    .A3(_09113_),
    .A4(_09115_),
    .ZN(_09116_));
 NOR4_X1 _31594_ (.A1(_09100_),
    .A2(_09103_),
    .A3(_09105_),
    .A4(_09116_),
    .ZN(_09117_));
 NAND2_X1 _31595_ (.A1(_08514_),
    .A2(_08672_),
    .ZN(_09118_));
 NOR2_X2 _31596_ (.A1(_08367_),
    .A2(_08467_),
    .ZN(_09119_));
 AOI222_X2 _31597_ (.A1(_08395_),
    .A2(_08490_),
    .B1(_08435_),
    .B2(_09119_),
    .C1(_08537_),
    .C2(_08375_),
    .ZN(_09120_));
 MUX2_X1 _31598_ (.A(_09118_),
    .B(_09120_),
    .S(_08488_),
    .Z(_09121_));
 OAI21_X1 _31599_ (.A(_09117_),
    .B1(_09121_),
    .B2(_08663_),
    .ZN(_09122_));
 OR3_X4 _31600_ (.A1(_08715_),
    .A2(_09099_),
    .A3(_09122_),
    .ZN(_09123_));
 NAND2_X4 _31601_ (.A1(_07662_),
    .A2(_09123_),
    .ZN(_09124_));
 CLKBUF_X3 _31602_ (.A(_07805_),
    .Z(_09125_));
 CLKBUF_X3 _31603_ (.A(_07228_),
    .Z(_09126_));
 XNOR2_X2 _31604_ (.A(_07317_),
    .B(_07895_),
    .ZN(_09127_));
 XOR2_X1 _31605_ (.A(_07306_),
    .B(_08041_),
    .Z(_09128_));
 XNOR2_X1 _31606_ (.A(_09127_),
    .B(_09128_),
    .ZN(_09129_));
 XNOR2_X1 _31607_ (.A(_00353_),
    .B(_09129_),
    .ZN(_09130_));
 BUF_X4 _31608_ (.A(_07231_),
    .Z(_09131_));
 MUX2_X1 _31609_ (.A(_08040_),
    .B(_09130_),
    .S(_09131_),
    .Z(_09132_));
 AOI22_X1 _31610_ (.A1(\block_reg[0][21] ),
    .A2(_09125_),
    .B1(_09126_),
    .B2(_09132_),
    .ZN(_09133_));
 CLKBUF_X3 _31611_ (.A(_07246_),
    .Z(_09134_));
 OAI22_X1 _31612_ (.A1(\block_reg[0][21] ),
    .A2(_09134_),
    .B1(_09007_),
    .B2(_09132_),
    .ZN(_09135_));
 INV_X1 _31613_ (.A(_09135_),
    .ZN(_09136_));
 MUX2_X1 _31614_ (.A(_09133_),
    .B(_09136_),
    .S(_03856_),
    .Z(_09137_));
 NAND2_X1 _31615_ (.A1(_09124_),
    .A2(_09137_),
    .ZN(_09138_));
 BUF_X2 _31616_ (.A(\core.enc_block.block_w0_reg[21] ),
    .Z(_09139_));
 MUX2_X1 _31617_ (.A(_09138_),
    .B(_09139_),
    .S(_08906_),
    .Z(_00715_));
 NAND3_X1 _31618_ (.A1(_09111_),
    .A2(_09113_),
    .A3(_09115_),
    .ZN(_09140_));
 NOR4_X2 _31619_ (.A1(_08347_),
    .A2(_08370_),
    .A3(_08256_),
    .A4(_08372_),
    .ZN(_09141_));
 AOI221_X2 _31620_ (.A(_09141_),
    .B1(_08537_),
    .B2(_08641_),
    .C1(_08676_),
    .C2(_08848_),
    .ZN(_09142_));
 NAND3_X1 _31621_ (.A1(_08561_),
    .A2(_08350_),
    .A3(_08828_),
    .ZN(_09143_));
 OAI21_X1 _31622_ (.A(_08691_),
    .B1(_08507_),
    .B2(_09079_),
    .ZN(_09144_));
 NOR4_X1 _31623_ (.A1(_08542_),
    .A2(_08551_),
    .A3(_08661_),
    .A4(_08400_),
    .ZN(_09145_));
 OAI21_X1 _31624_ (.A(_08485_),
    .B1(_09093_),
    .B2(_09145_),
    .ZN(_09146_));
 NAND4_X1 _31625_ (.A1(_09142_),
    .A2(_09143_),
    .A3(_09144_),
    .A4(_09146_),
    .ZN(_09147_));
 OR4_X1 _31626_ (.A1(_08454_),
    .A2(_08861_),
    .A3(_09055_),
    .A4(_09056_),
    .ZN(_09148_));
 NOR2_X1 _31627_ (.A1(_08312_),
    .A2(_08290_),
    .ZN(_09149_));
 AOI221_X2 _31628_ (.A(_08281_),
    .B1(_08506_),
    .B2(_09149_),
    .C1(_08787_),
    .C2(_08367_),
    .ZN(_09150_));
 AOI22_X1 _31629_ (.A1(_08635_),
    .A2(_08335_),
    .B1(_08374_),
    .B2(_08665_),
    .ZN(_09151_));
 AOI21_X1 _31630_ (.A(_09150_),
    .B1(_09151_),
    .B2(_08282_),
    .ZN(_09152_));
 OR4_X1 _31631_ (.A1(_09140_),
    .A2(_09147_),
    .A3(_09148_),
    .A4(_09152_),
    .ZN(_09153_));
 OAI21_X1 _31632_ (.A(_08754_),
    .B1(_08582_),
    .B2(_08529_),
    .ZN(_09154_));
 AOI22_X1 _31633_ (.A1(_08555_),
    .A2(_08819_),
    .B1(_09154_),
    .B2(_08520_),
    .ZN(_09155_));
 NOR2_X1 _31634_ (.A1(_08515_),
    .A2(_09155_),
    .ZN(_09156_));
 AOI22_X2 _31635_ (.A1(_08786_),
    .A2(_08506_),
    .B1(_08674_),
    .B2(_09072_),
    .ZN(_09157_));
 AOI21_X1 _31636_ (.A(_09077_),
    .B1(_08490_),
    .B2(_08523_),
    .ZN(_09158_));
 OR2_X1 _31637_ (.A1(_08503_),
    .A2(_09158_),
    .ZN(_09159_));
 NOR2_X1 _31638_ (.A1(_08486_),
    .A2(_08542_),
    .ZN(_09160_));
 AOI22_X2 _31639_ (.A1(_09119_),
    .A2(_08374_),
    .B1(_08537_),
    .B2(_09160_),
    .ZN(_09161_));
 OR2_X1 _31640_ (.A1(_08488_),
    .A2(_09161_),
    .ZN(_09162_));
 NAND4_X1 _31641_ (.A1(_08801_),
    .A2(_09157_),
    .A3(_09159_),
    .A4(_09162_),
    .ZN(_09163_));
 NAND2_X1 _31642_ (.A1(_08492_),
    .A2(_08841_),
    .ZN(_09164_));
 AND4_X1 _31643_ (.A1(_08845_),
    .A2(_08847_),
    .A3(_08849_),
    .A4(_08852_),
    .ZN(_09165_));
 OAI33_X1 _31644_ (.A1(_08282_),
    .A2(_08343_),
    .A3(_08348_),
    .B1(_08269_),
    .B2(_08557_),
    .B3(_08375_),
    .ZN(_09166_));
 OAI33_X1 _31645_ (.A1(_08514_),
    .A2(_08402_),
    .A3(_08518_),
    .B1(_08398_),
    .B2(_08460_),
    .B3(_08581_),
    .ZN(_09167_));
 OAI21_X1 _31646_ (.A(_08492_),
    .B1(_09166_),
    .B2(_09167_),
    .ZN(_09168_));
 NAND4_X2 _31647_ (.A1(_08640_),
    .A2(_09164_),
    .A3(_09165_),
    .A4(_09168_),
    .ZN(_09169_));
 OR4_X4 _31648_ (.A1(_09153_),
    .A2(_09156_),
    .A3(_09163_),
    .A4(_09169_),
    .ZN(_09170_));
 NOR2_X4 _31649_ (.A1(_08483_),
    .A2(_09170_),
    .ZN(_09171_));
 NOR2_X4 _31650_ (.A1(_06707_),
    .A2(_09171_),
    .ZN(_09172_));
 XNOR2_X2 _31651_ (.A(_07306_),
    .B(_08040_),
    .ZN(_09173_));
 XOR2_X1 _31652_ (.A(_07329_),
    .B(_08107_),
    .Z(_09174_));
 XNOR2_X1 _31653_ (.A(_09173_),
    .B(_09174_),
    .ZN(_09175_));
 XNOR2_X1 _31654_ (.A(_00356_),
    .B(_09175_),
    .ZN(_09176_));
 MUX2_X1 _31655_ (.A(_08106_),
    .B(_09176_),
    .S(_07242_),
    .Z(_09177_));
 AOI22_X1 _31656_ (.A1(\block_reg[0][22] ),
    .A2(_07806_),
    .B1(_08599_),
    .B2(_09177_),
    .ZN(_09178_));
 INV_X1 _31657_ (.A(_09178_),
    .ZN(_09179_));
 OAI22_X1 _31658_ (.A1(\block_reg[0][22] ),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_09177_),
    .ZN(_09180_));
 MUX2_X1 _31659_ (.A(_09179_),
    .B(_09180_),
    .S(_03914_),
    .Z(_09181_));
 NOR3_X1 _31660_ (.A1(_08177_),
    .A2(_09172_),
    .A3(_09181_),
    .ZN(_09182_));
 BUF_X2 _31661_ (.A(\core.enc_block.block_w0_reg[22] ),
    .Z(_09183_));
 INV_X1 _31662_ (.A(_09183_),
    .ZN(_09184_));
 AOI21_X1 _31663_ (.A(_09182_),
    .B1(_06705_),
    .B2(_09184_),
    .ZN(_00716_));
 OAI33_X1 _31664_ (.A1(_08443_),
    .A2(_08545_),
    .A3(_08409_),
    .B1(_08399_),
    .B2(_08423_),
    .B3(_08312_),
    .ZN(_09185_));
 AOI221_X1 _31665_ (.A(_08787_),
    .B1(_08689_),
    .B2(_08676_),
    .C1(_09185_),
    .C2(_08639_),
    .ZN(_09186_));
 OR2_X1 _31666_ (.A1(_08515_),
    .A2(_09186_),
    .ZN(_09187_));
 AND4_X2 _31667_ (.A1(_08353_),
    .A2(_08567_),
    .A3(_08693_),
    .A4(_09187_),
    .ZN(_09188_));
 OAI221_X2 _31668_ (.A(_09157_),
    .B1(_09158_),
    .B2(_08503_),
    .C1(_09161_),
    .C2(_08488_),
    .ZN(_09189_));
 NOR2_X1 _31669_ (.A1(_08467_),
    .A2(_08443_),
    .ZN(_09190_));
 XNOR2_X1 _31670_ (.A(_08375_),
    .B(_09190_),
    .ZN(_09191_));
 NOR4_X2 _31671_ (.A1(_08361_),
    .A2(_08518_),
    .A3(_08833_),
    .A4(_09191_),
    .ZN(_09192_));
 NOR4_X4 _31672_ (.A1(_08863_),
    .A2(_09019_),
    .A3(_09189_),
    .A4(_09192_),
    .ZN(_09193_));
 AOI21_X1 _31673_ (.A(_08544_),
    .B1(_08505_),
    .B2(_08514_),
    .ZN(_09194_));
 AOI22_X2 _31674_ (.A1(_08680_),
    .A2(_08435_),
    .B1(_08540_),
    .B2(_08817_),
    .ZN(_09195_));
 OAI221_X2 _31675_ (.A(_08788_),
    .B1(_09194_),
    .B2(_08217_),
    .C1(_09195_),
    .C2(_08398_),
    .ZN(_09196_));
 NOR4_X2 _31676_ (.A1(_08516_),
    .A2(_08517_),
    .A3(_08306_),
    .A4(_08534_),
    .ZN(_09197_));
 NOR4_X2 _31677_ (.A1(_08282_),
    .A2(_08518_),
    .A3(_08274_),
    .A4(_08661_),
    .ZN(_09198_));
 NOR4_X2 _31678_ (.A1(_08517_),
    .A2(_08551_),
    .A3(_08256_),
    .A4(_08400_),
    .ZN(_09199_));
 NOR4_X2 _31679_ (.A1(_08661_),
    .A2(_08400_),
    .A3(_08507_),
    .A4(_08633_),
    .ZN(_09200_));
 NOR4_X2 _31680_ (.A1(_09197_),
    .A2(_09198_),
    .A3(_09199_),
    .A4(_09200_),
    .ZN(_09201_));
 OAI33_X1 _31681_ (.A1(_08414_),
    .A2(_08683_),
    .A3(_08661_),
    .B1(_08409_),
    .B2(_08545_),
    .B3(_08519_),
    .ZN(_09202_));
 AOI22_X2 _31682_ (.A1(_08337_),
    .A2(_08846_),
    .B1(_09202_),
    .B2(_08198_),
    .ZN(_09203_));
 NAND4_X2 _31683_ (.A1(_08232_),
    .A2(_08230_),
    .A3(_08258_),
    .A4(_08411_),
    .ZN(_09204_));
 AOI211_X2 _31684_ (.A(_08274_),
    .B(_09204_),
    .C1(_08620_),
    .C2(_08621_),
    .ZN(_09205_));
 AOI22_X2 _31685_ (.A1(_08697_),
    .A2(_08447_),
    .B1(_09205_),
    .B2(_08564_),
    .ZN(_09206_));
 OAI221_X2 _31686_ (.A(_09201_),
    .B1(_09203_),
    .B2(_08306_),
    .C1(_08283_),
    .C2(_09206_),
    .ZN(_09207_));
 NOR4_X4 _31687_ (.A1(_09103_),
    .A2(_09105_),
    .A3(_09196_),
    .A4(_09207_),
    .ZN(_09208_));
 NAND3_X4 _31688_ (.A1(_09188_),
    .A2(_09193_),
    .A3(_09208_),
    .ZN(_09209_));
 NAND2_X2 _31689_ (.A1(_07662_),
    .A2(_09209_),
    .ZN(_09210_));
 CLKBUF_X3 _31690_ (.A(_07228_),
    .Z(_09211_));
 NOR2_X1 _31691_ (.A1(_08165_),
    .A2(_08722_),
    .ZN(_09212_));
 XNOR2_X1 _31692_ (.A(_08106_),
    .B(_07235_),
    .ZN(_09213_));
 XNOR2_X1 _31693_ (.A(_07329_),
    .B(_07338_),
    .ZN(_09214_));
 XNOR2_X1 _31694_ (.A(_09213_),
    .B(_09214_),
    .ZN(_09215_));
 XNOR2_X1 _31695_ (.A(_06742_),
    .B(_09215_),
    .ZN(_09216_));
 BUF_X4 _31696_ (.A(_07651_),
    .Z(_09217_));
 AOI21_X2 _31697_ (.A(_09212_),
    .B1(_09216_),
    .B2(_09217_),
    .ZN(_09218_));
 AOI22_X1 _31698_ (.A1(\block_reg[0][23] ),
    .A2(_09005_),
    .B1(_09211_),
    .B2(_09218_),
    .ZN(_09219_));
 NAND2_X1 _31699_ (.A1(_03975_),
    .A2(_09219_),
    .ZN(_09220_));
 BUF_X4 _31700_ (.A(_09134_),
    .Z(_09221_));
 CLKBUF_X3 _31701_ (.A(_07253_),
    .Z(_09222_));
 BUF_X4 _31702_ (.A(_09222_),
    .Z(_09223_));
 OAI22_X1 _31703_ (.A1(\block_reg[0][23] ),
    .A2(_09221_),
    .B1(_09223_),
    .B2(_09218_),
    .ZN(_09224_));
 OAI21_X2 _31704_ (.A(_09220_),
    .B1(_09224_),
    .B2(_03975_),
    .ZN(_09225_));
 NAND2_X1 _31705_ (.A1(_09210_),
    .A2(_09225_),
    .ZN(_09226_));
 CLKBUF_X3 _31706_ (.A(\core.enc_block.block_w0_reg[23] ),
    .Z(_09227_));
 MUX2_X1 _31707_ (.A(_09226_),
    .B(_09227_),
    .S(_08906_),
    .Z(_00717_));
 INV_X1 _31708_ (.A(_07234_),
    .ZN(_09228_));
 BUF_X4 _31709_ (.A(_00346_),
    .Z(_09229_));
 OR2_X4 _31710_ (.A1(_09229_),
    .A2(_06919_),
    .ZN(_09230_));
 CLKBUF_X3 _31711_ (.A(\core.enc_block.block_w2_reg[27] ),
    .Z(_09231_));
 AOI21_X1 _31712_ (.A(_06866_),
    .B1(_09231_),
    .B2(_07264_),
    .ZN(_09232_));
 BUF_X2 _31713_ (.A(\core.enc_block.block_w1_reg[27] ),
    .Z(_09233_));
 INV_X1 _31714_ (.A(_09233_),
    .ZN(_09234_));
 OAI221_X2 _31715_ (.A(_09232_),
    .B1(_07266_),
    .B2(_09234_),
    .C1(_00348_),
    .C2(_16252_),
    .ZN(_09235_));
 NAND2_X2 _31716_ (.A1(_06702_),
    .A2(_00347_),
    .ZN(_09236_));
 NAND4_X4 _31717_ (.A1(_06698_),
    .A2(_07419_),
    .A3(_09235_),
    .A4(_09236_),
    .ZN(_09237_));
 BUF_X4 _31718_ (.A(_00345_),
    .Z(_09238_));
 OR2_X4 _31719_ (.A1(_09238_),
    .A2(_06919_),
    .ZN(_09239_));
 CLKBUF_X3 _31720_ (.A(\core.enc_block.block_w1_reg[26] ),
    .Z(_09240_));
 AOI21_X1 _31721_ (.A(_06725_),
    .B1(_09240_),
    .B2(_06718_),
    .ZN(_09241_));
 INV_X1 _31722_ (.A(_07264_),
    .ZN(_09242_));
 BUF_X2 _31723_ (.A(\core.enc_block.block_w2_reg[26] ),
    .Z(_09243_));
 INV_X1 _31724_ (.A(_09243_),
    .ZN(_09244_));
 INV_X2 _31725_ (.A(\core.enc_block.block_w3_reg[26] ),
    .ZN(_09245_));
 OAI221_X2 _31726_ (.A(_09241_),
    .B1(_09242_),
    .B2(_09244_),
    .C1(_09245_),
    .C2(_16251_),
    .ZN(_09246_));
 INV_X1 _31727_ (.A(_07643_),
    .ZN(_09247_));
 NAND2_X1 _31728_ (.A1(_06866_),
    .A2(_09247_),
    .ZN(_09248_));
 NAND4_X4 _31729_ (.A1(_06698_),
    .A2(_06822_),
    .A3(_09246_),
    .A4(_09248_),
    .ZN(_09249_));
 AOI22_X4 _31730_ (.A1(_09230_),
    .A2(_09237_),
    .B1(_09239_),
    .B2(_09249_),
    .ZN(_09250_));
 BUF_X4 _31731_ (.A(_09250_),
    .Z(_09251_));
 NAND2_X2 _31732_ (.A1(_06702_),
    .A2(_00339_),
    .ZN(_09252_));
 BUF_X4 _31733_ (.A(\core.enc_block.block_w1_reg[31] ),
    .Z(_09253_));
 AOI21_X1 _31734_ (.A(_06866_),
    .B1(_09253_),
    .B2(_06718_),
    .ZN(_09254_));
 BUF_X4 _31735_ (.A(\core.enc_block.block_w2_reg[31] ),
    .Z(_09255_));
 INV_X1 _31736_ (.A(_09255_),
    .ZN(_09256_));
 OAI221_X2 _31737_ (.A(_09254_),
    .B1(_09242_),
    .B2(_09256_),
    .C1(_00340_),
    .C2(_16252_),
    .ZN(_09257_));
 NAND4_X4 _31738_ (.A1(_06698_),
    .A2(_06837_),
    .A3(_09252_),
    .A4(_09257_),
    .ZN(_09258_));
 NAND2_X1 _31739_ (.A1(_06702_),
    .A2(_00336_),
    .ZN(_09259_));
 BUF_X2 _31740_ (.A(\core.enc_block.block_w1_reg[30] ),
    .Z(_09260_));
 AOI21_X1 _31741_ (.A(_06701_),
    .B1(_09260_),
    .B2(_06718_),
    .ZN(_09261_));
 BUF_X2 _31742_ (.A(\core.enc_block.block_w2_reg[30] ),
    .Z(_09262_));
 INV_X1 _31743_ (.A(_09262_),
    .ZN(_09263_));
 OAI221_X2 _31744_ (.A(_09261_),
    .B1(_09242_),
    .B2(_09263_),
    .C1(_00337_),
    .C2(_16252_),
    .ZN(_09264_));
 AND4_X2 _31745_ (.A1(_06697_),
    .A2(_07315_),
    .A3(_09259_),
    .A4(_09264_),
    .ZN(_09265_));
 BUF_X4 _31746_ (.A(_09265_),
    .Z(_09266_));
 NOR2_X4 _31747_ (.A1(_00335_),
    .A2(_06837_),
    .ZN(_09267_));
 CLKBUF_X3 _31748_ (.A(\core.keymem.prev_key1_reg[31] ),
    .Z(_09268_));
 INV_X1 _31749_ (.A(_09268_),
    .ZN(_09269_));
 OAI221_X2 _31750_ (.A(_09258_),
    .B1(_09266_),
    .B2(_09267_),
    .C1(_07486_),
    .C2(_09269_),
    .ZN(_09270_));
 BUF_X4 _31751_ (.A(_09270_),
    .Z(_09271_));
 BUF_X4 _31752_ (.A(_09271_),
    .Z(_09272_));
 INV_X2 _31753_ (.A(_00332_),
    .ZN(_09273_));
 NAND2_X4 _31754_ (.A1(_09273_),
    .A2(_06938_),
    .ZN(_09274_));
 CLKBUF_X3 _31755_ (.A(\core.enc_block.block_w2_reg[29] ),
    .Z(_09275_));
 AOI21_X1 _31756_ (.A(_06701_),
    .B1(_09275_),
    .B2(_07264_),
    .ZN(_09276_));
 CLKBUF_X3 _31757_ (.A(\core.enc_block.block_w1_reg[29] ),
    .Z(_09277_));
 INV_X1 _31758_ (.A(_09277_),
    .ZN(_09278_));
 OAI221_X2 _31759_ (.A(_09276_),
    .B1(_07266_),
    .B2(_09278_),
    .C1(_00334_),
    .C2(_16252_),
    .ZN(_09279_));
 NAND2_X1 _31760_ (.A1(_06702_),
    .A2(_00333_),
    .ZN(_09280_));
 NAND4_X4 _31761_ (.A1(_06843_),
    .A2(_06837_),
    .A3(_09279_),
    .A4(_09280_),
    .ZN(_09281_));
 CLKBUF_X3 _31762_ (.A(\core.keymem.prev_key1_reg[28] ),
    .Z(_09282_));
 NAND2_X4 _31763_ (.A1(_09282_),
    .A2(_06936_),
    .ZN(_09283_));
 AOI21_X1 _31764_ (.A(_06725_),
    .B1(_07264_),
    .B2(\core.enc_block.block_w2_reg[28] ),
    .ZN(_09284_));
 CLKBUF_X2 _31765_ (.A(\core.enc_block.block_w1_reg[28] ),
    .Z(_09285_));
 INV_X1 _31766_ (.A(_09285_),
    .ZN(_09286_));
 OAI221_X2 _31767_ (.A(_09284_),
    .B1(_07266_),
    .B2(_09286_),
    .C1(_00331_),
    .C2(_16252_),
    .ZN(_09287_));
 NAND2_X2 _31768_ (.A1(_00330_),
    .A2(_06702_),
    .ZN(_09288_));
 NAND4_X4 _31769_ (.A1(_06698_),
    .A2(_06822_),
    .A3(_09287_),
    .A4(_09288_),
    .ZN(_09289_));
 NAND4_X4 _31770_ (.A1(_09274_),
    .A2(_09281_),
    .A3(_09283_),
    .A4(_09289_),
    .ZN(_09290_));
 BUF_X4 _31771_ (.A(_09290_),
    .Z(_09291_));
 NOR2_X4 _31772_ (.A1(_09272_),
    .A2(_09291_),
    .ZN(_09292_));
 BUF_X4 _31773_ (.A(_09292_),
    .Z(_09293_));
 BUF_X4 _31774_ (.A(_09271_),
    .Z(_09294_));
 CLKBUF_X3 _31775_ (.A(_09294_),
    .Z(_09295_));
 NOR2_X4 _31776_ (.A1(_00332_),
    .A2(_07419_),
    .ZN(_09296_));
 AND4_X2 _31777_ (.A1(_06697_),
    .A2(_06820_),
    .A3(_09279_),
    .A4(_09280_),
    .ZN(_09297_));
 BUF_X4 _31778_ (.A(_09297_),
    .Z(_09298_));
 INV_X2 _31779_ (.A(_09282_),
    .ZN(_09299_));
 NOR2_X4 _31780_ (.A1(_09299_),
    .A2(_07419_),
    .ZN(_09300_));
 AND4_X2 _31781_ (.A1(_06697_),
    .A2(_06820_),
    .A3(_09287_),
    .A4(_09288_),
    .ZN(_09301_));
 BUF_X4 _31782_ (.A(_09301_),
    .Z(_09302_));
 OAI22_X4 _31783_ (.A1(_09296_),
    .A2(_09298_),
    .B1(_09300_),
    .B2(_09302_),
    .ZN(_09303_));
 BUF_X4 _31784_ (.A(_09303_),
    .Z(_09304_));
 BUF_X4 _31785_ (.A(_09304_),
    .Z(_09305_));
 BUF_X4 _31786_ (.A(_09305_),
    .Z(_09306_));
 BUF_X4 _31787_ (.A(_09306_),
    .Z(_09307_));
 CLKBUF_X3 _31788_ (.A(_00342_),
    .Z(_09308_));
 NOR2_X4 _31789_ (.A1(_09308_),
    .A2(_07419_),
    .ZN(_09309_));
 CLKBUF_X3 _31790_ (.A(\core.enc_block.block_w2_reg[25] ),
    .Z(_09310_));
 AOI21_X1 _31791_ (.A(_06866_),
    .B1(_09310_),
    .B2(_07264_),
    .ZN(_09311_));
 BUF_X4 _31792_ (.A(\core.enc_block.block_w1_reg[25] ),
    .Z(_09312_));
 INV_X1 _31793_ (.A(_09312_),
    .ZN(_09313_));
 OAI221_X2 _31794_ (.A(_09311_),
    .B1(_07266_),
    .B2(_09313_),
    .C1(_00344_),
    .C2(_16252_),
    .ZN(_09314_));
 NAND2_X2 _31795_ (.A1(_06702_),
    .A2(_00343_),
    .ZN(_09315_));
 AND4_X4 _31796_ (.A1(_06697_),
    .A2(_07315_),
    .A3(_09314_),
    .A4(_09315_),
    .ZN(_09316_));
 BUF_X8 _31797_ (.A(_09316_),
    .Z(_09317_));
 CLKBUF_X3 _31798_ (.A(\core.keymem.prev_key1_reg[24] ),
    .Z(_09318_));
 INV_X1 _31799_ (.A(_09318_),
    .ZN(_09319_));
 NOR2_X4 _31800_ (.A1(_09319_),
    .A2(_06837_),
    .ZN(_09320_));
 CLKBUF_X3 _31801_ (.A(\core.enc_block.block_w2_reg[24] ),
    .Z(_09321_));
 AOI21_X1 _31802_ (.A(_06701_),
    .B1(_09321_),
    .B2(_07264_),
    .ZN(_09322_));
 BUF_X4 _31803_ (.A(\core.enc_block.block_w1_reg[24] ),
    .Z(_09323_));
 INV_X1 _31804_ (.A(_09323_),
    .ZN(_09324_));
 OAI221_X2 _31805_ (.A(_09322_),
    .B1(_07266_),
    .B2(_09324_),
    .C1(_00341_),
    .C2(_16252_),
    .ZN(_09325_));
 NAND2_X2 _31806_ (.A1(_06702_),
    .A2(_09228_),
    .ZN(_09326_));
 AND4_X2 _31807_ (.A1(_06697_),
    .A2(_06820_),
    .A3(_09325_),
    .A4(_09326_),
    .ZN(_09327_));
 BUF_X4 _31808_ (.A(_09327_),
    .Z(_09328_));
 NOR4_X4 _31809_ (.A1(_09309_),
    .A2(_09317_),
    .A3(_09320_),
    .A4(_09328_),
    .ZN(_09329_));
 BUF_X4 _31810_ (.A(_09329_),
    .Z(_09330_));
 NOR3_X2 _31811_ (.A1(_09295_),
    .A2(_09307_),
    .A3(_09330_),
    .ZN(_09331_));
 NOR2_X4 _31812_ (.A1(_09320_),
    .A2(_09328_),
    .ZN(_09332_));
 BUF_X4 _31813_ (.A(_09332_),
    .Z(_09333_));
 BUF_X4 _31814_ (.A(_09333_),
    .Z(_09334_));
 BUF_X4 _31815_ (.A(_09334_),
    .Z(_09335_));
 NOR2_X4 _31816_ (.A1(_09309_),
    .A2(_09317_),
    .ZN(_09336_));
 BUF_X4 _31817_ (.A(_09336_),
    .Z(_09337_));
 BUF_X4 _31818_ (.A(_09337_),
    .Z(_09338_));
 OAI221_X1 _31819_ (.A(_09251_),
    .B1(_09293_),
    .B2(_09331_),
    .C1(_09335_),
    .C2(_09338_),
    .ZN(_09339_));
 NAND2_X4 _31820_ (.A1(_09318_),
    .A2(_06936_),
    .ZN(_09340_));
 NAND4_X4 _31821_ (.A1(_06698_),
    .A2(_06886_),
    .A3(_09325_),
    .A4(_09326_),
    .ZN(_09341_));
 NAND2_X1 _31822_ (.A1(_09340_),
    .A2(_09341_),
    .ZN(_09342_));
 BUF_X4 _31823_ (.A(_09342_),
    .Z(_09343_));
 NAND4_X4 _31824_ (.A1(_09230_),
    .A2(_09237_),
    .A3(_09239_),
    .A4(_09249_),
    .ZN(_09344_));
 BUF_X4 _31825_ (.A(_09344_),
    .Z(_09345_));
 NOR2_X2 _31826_ (.A1(_09343_),
    .A2(_09345_),
    .ZN(_09346_));
 AOI22_X4 _31827_ (.A1(_09274_),
    .A2(_09281_),
    .B1(_09283_),
    .B2(_09289_),
    .ZN(_09347_));
 NAND4_X4 _31828_ (.A1(_06698_),
    .A2(_06837_),
    .A3(_09259_),
    .A4(_09264_),
    .ZN(_09348_));
 BUF_X2 _31829_ (.A(\core.keymem.prev_key1_reg[30] ),
    .Z(_09349_));
 NAND2_X2 _31830_ (.A1(_09349_),
    .A2(_06938_),
    .ZN(_09350_));
 NAND2_X4 _31831_ (.A1(_09268_),
    .A2(_06938_),
    .ZN(_09351_));
 AND4_X1 _31832_ (.A1(_09258_),
    .A2(_09348_),
    .A3(_09350_),
    .A4(_09351_),
    .ZN(_09352_));
 CLKBUF_X3 _31833_ (.A(_09352_),
    .Z(_09353_));
 NAND2_X1 _31834_ (.A1(_09347_),
    .A2(_09353_),
    .ZN(_09354_));
 NOR2_X1 _31835_ (.A1(_09338_),
    .A2(_09354_),
    .ZN(_09355_));
 NOR2_X4 _31836_ (.A1(_00338_),
    .A2(_07419_),
    .ZN(_09356_));
 AND4_X4 _31837_ (.A1(_06843_),
    .A2(_06757_),
    .A3(_09252_),
    .A4(_09257_),
    .ZN(_09357_));
 INV_X2 _31838_ (.A(_09349_),
    .ZN(_09358_));
 OAI221_X2 _31839_ (.A(_09348_),
    .B1(_09356_),
    .B2(_09357_),
    .C1(_09358_),
    .C2(_06934_),
    .ZN(_09359_));
 BUF_X4 _31840_ (.A(_09359_),
    .Z(_09360_));
 BUF_X8 _31841_ (.A(_09360_),
    .Z(_09361_));
 NOR2_X4 _31842_ (.A1(_09361_),
    .A2(_09304_),
    .ZN(_09362_));
 OAI21_X1 _31843_ (.A(_09346_),
    .B1(_09355_),
    .B2(_09362_),
    .ZN(_09363_));
 BUF_X4 _31844_ (.A(_09360_),
    .Z(_09364_));
 NOR4_X4 _31845_ (.A1(_09336_),
    .A2(_09364_),
    .A3(_09305_),
    .A4(_09345_),
    .ZN(_09365_));
 NOR2_X4 _31846_ (.A1(_09229_),
    .A2(_07419_),
    .ZN(_09366_));
 AND4_X2 _31847_ (.A1(_06697_),
    .A2(_07315_),
    .A3(_09235_),
    .A4(_09236_),
    .ZN(_09367_));
 BUF_X4 _31848_ (.A(_09367_),
    .Z(_09368_));
 OAI22_X4 _31849_ (.A1(_09366_),
    .A2(_09368_),
    .B1(_09309_),
    .B2(_09317_),
    .ZN(_09369_));
 BUF_X4 _31850_ (.A(_09369_),
    .Z(_09370_));
 OAI221_X2 _31851_ (.A(_09249_),
    .B1(_09320_),
    .B2(_09328_),
    .C1(_06888_),
    .C2(_09238_),
    .ZN(_09371_));
 NOR2_X2 _31852_ (.A1(_09370_),
    .A2(_09371_),
    .ZN(_09372_));
 NOR2_X2 _31853_ (.A1(_09271_),
    .A2(_09304_),
    .ZN(_09373_));
 BUF_X4 _31854_ (.A(_09373_),
    .Z(_09374_));
 OAI22_X4 _31855_ (.A1(_09357_),
    .A2(_09356_),
    .B1(_09266_),
    .B2(_09267_),
    .ZN(_09375_));
 NOR2_X4 _31856_ (.A1(_09304_),
    .A2(_09375_),
    .ZN(_09376_));
 INV_X2 _31857_ (.A(_09308_),
    .ZN(_09377_));
 NAND2_X4 _31858_ (.A1(_09377_),
    .A2(_06936_),
    .ZN(_09378_));
 NAND4_X4 _31859_ (.A1(_06698_),
    .A2(_07419_),
    .A3(_09314_),
    .A4(_09315_),
    .ZN(_09379_));
 NAND4_X4 _31860_ (.A1(_09230_),
    .A2(_09237_),
    .A3(_09378_),
    .A4(_09379_),
    .ZN(_09380_));
 NOR2_X4 _31861_ (.A1(_09380_),
    .A2(_09371_),
    .ZN(_09381_));
 AOI221_X2 _31862_ (.A(_09365_),
    .B1(_09372_),
    .B2(_09374_),
    .C1(_09376_),
    .C2(_09381_),
    .ZN(_09382_));
 BUF_X4 _31863_ (.A(_09343_),
    .Z(_09383_));
 BUF_X4 _31864_ (.A(_09383_),
    .Z(_09384_));
 NOR2_X4 _31865_ (.A1(_09366_),
    .A2(_09368_),
    .ZN(_09385_));
 NAND2_X2 _31866_ (.A1(_09239_),
    .A2(_09249_),
    .ZN(_09386_));
 NOR2_X4 _31867_ (.A1(_09385_),
    .A2(_09386_),
    .ZN(_09387_));
 NAND3_X1 _31868_ (.A1(_09384_),
    .A2(_09293_),
    .A3(_09387_),
    .ZN(_09388_));
 AND4_X2 _31869_ (.A1(_09339_),
    .A2(_09363_),
    .A3(_09382_),
    .A4(_09388_),
    .ZN(_09389_));
 BUF_X4 _31870_ (.A(_09386_),
    .Z(_09390_));
 NAND4_X4 _31871_ (.A1(_09258_),
    .A2(_09348_),
    .A3(_09350_),
    .A4(_09351_),
    .ZN(_09391_));
 BUF_X4 _31872_ (.A(_09391_),
    .Z(_09392_));
 NOR4_X2 _31873_ (.A1(_09390_),
    .A2(_09304_),
    .A3(_09392_),
    .A4(_09380_),
    .ZN(_09393_));
 NOR2_X4 _31874_ (.A1(_09238_),
    .A2(_06757_),
    .ZN(_09394_));
 AND4_X2 _31875_ (.A1(_06733_),
    .A2(_06711_),
    .A3(_09246_),
    .A4(_09248_),
    .ZN(_09395_));
 BUF_X4 _31876_ (.A(_09395_),
    .Z(_09396_));
 OAI221_X2 _31877_ (.A(_09237_),
    .B1(_09394_),
    .B2(_09396_),
    .C1(_06934_),
    .C2(_09229_),
    .ZN(_09397_));
 BUF_X4 _31878_ (.A(_09397_),
    .Z(_09398_));
 NAND4_X4 _31879_ (.A1(_09378_),
    .A2(_09379_),
    .A3(_09340_),
    .A4(_09341_),
    .ZN(_09399_));
 NOR2_X4 _31880_ (.A1(_09398_),
    .A2(_09399_),
    .ZN(_09400_));
 NOR2_X4 _31881_ (.A1(_09375_),
    .A2(_09290_),
    .ZN(_09401_));
 OAI22_X4 _31882_ (.A1(_09366_),
    .A2(_09368_),
    .B1(_09394_),
    .B2(_09396_),
    .ZN(_09402_));
 NOR2_X2 _31883_ (.A1(_09336_),
    .A2(_09402_),
    .ZN(_09403_));
 AOI221_X2 _31884_ (.A(_09393_),
    .B1(_09400_),
    .B2(_09401_),
    .C1(_09292_),
    .C2(_09403_),
    .ZN(_09404_));
 NOR2_X4 _31885_ (.A1(_09361_),
    .A2(_09291_),
    .ZN(_09405_));
 BUF_X4 _31886_ (.A(_09375_),
    .Z(_09406_));
 BUF_X4 _31887_ (.A(_09406_),
    .Z(_09407_));
 BUF_X4 _31888_ (.A(_09291_),
    .Z(_09408_));
 NOR3_X2 _31889_ (.A1(_09407_),
    .A2(_09408_),
    .A3(_09330_),
    .ZN(_09409_));
 AOI22_X4 _31890_ (.A1(_09239_),
    .A2(_09249_),
    .B1(_09378_),
    .B2(_09379_),
    .ZN(_09410_));
 NOR3_X2 _31891_ (.A1(_09364_),
    .A2(_09408_),
    .A3(_09410_),
    .ZN(_09411_));
 BUF_X4 _31892_ (.A(_09385_),
    .Z(_09412_));
 BUF_X4 _31893_ (.A(_09412_),
    .Z(_09413_));
 OAI22_X4 _31894_ (.A1(_09405_),
    .A2(_09409_),
    .B1(_09411_),
    .B2(_09413_),
    .ZN(_09414_));
 BUF_X4 _31895_ (.A(_09390_),
    .Z(_09415_));
 AOI221_X2 _31896_ (.A(_09328_),
    .B1(_09379_),
    .B2(_09378_),
    .C1(_09318_),
    .C2(_07108_),
    .ZN(_09416_));
 BUF_X4 _31897_ (.A(_09416_),
    .Z(_09417_));
 NAND2_X2 _31898_ (.A1(_09412_),
    .A2(_09417_),
    .ZN(_09418_));
 AOI21_X2 _31899_ (.A(_09415_),
    .B1(_09405_),
    .B2(_09418_),
    .ZN(_09419_));
 OAI21_X4 _31900_ (.A(_09404_),
    .B1(_09414_),
    .B2(_09419_),
    .ZN(_09420_));
 OAI221_X2 _31901_ (.A(_09379_),
    .B1(_09320_),
    .B2(_09328_),
    .C1(_07486_),
    .C2(_09308_),
    .ZN(_09421_));
 BUF_X4 _31902_ (.A(_09421_),
    .Z(_09422_));
 BUF_X4 _31903_ (.A(_09392_),
    .Z(_09423_));
 BUF_X4 _31904_ (.A(_09423_),
    .Z(_09424_));
 OAI221_X2 _31905_ (.A(_09249_),
    .B1(_09368_),
    .B2(_09366_),
    .C1(_09238_),
    .C2(_06934_),
    .ZN(_09425_));
 BUF_X4 _31906_ (.A(_09425_),
    .Z(_09426_));
 BUF_X4 _31907_ (.A(_09426_),
    .Z(_09427_));
 NOR3_X1 _31908_ (.A1(_09424_),
    .A2(_09291_),
    .A3(_09427_),
    .ZN(_09428_));
 NOR4_X2 _31909_ (.A1(_09305_),
    .A2(_09406_),
    .A3(_09333_),
    .A4(_09398_),
    .ZN(_09429_));
 OAI21_X2 _31910_ (.A(_09422_),
    .B1(_09428_),
    .B2(_09429_),
    .ZN(_09430_));
 OAI221_X2 _31911_ (.A(_09289_),
    .B1(_09298_),
    .B2(_09296_),
    .C1(_09299_),
    .C2(_07486_),
    .ZN(_09431_));
 BUF_X4 _31912_ (.A(_09431_),
    .Z(_09432_));
 BUF_X4 _31913_ (.A(_09432_),
    .Z(_09433_));
 NOR4_X4 _31914_ (.A1(_09433_),
    .A2(_09423_),
    .A3(_09427_),
    .A4(_09329_),
    .ZN(_09434_));
 NOR3_X2 _31915_ (.A1(_09305_),
    .A2(_09423_),
    .A3(_09402_),
    .ZN(_09435_));
 NAND2_X2 _31916_ (.A1(_09230_),
    .A2(_09237_),
    .ZN(_09436_));
 BUF_X4 _31917_ (.A(_09436_),
    .Z(_09437_));
 NAND2_X2 _31918_ (.A1(_09274_),
    .A2(_09281_),
    .ZN(_09438_));
 BUF_X4 _31919_ (.A(_09438_),
    .Z(_09439_));
 NOR4_X4 _31920_ (.A1(_09437_),
    .A2(_09390_),
    .A3(_09439_),
    .A4(_09375_),
    .ZN(_09440_));
 NOR3_X4 _31921_ (.A1(_09361_),
    .A2(_09433_),
    .A3(_09369_),
    .ZN(_09441_));
 NOR4_X4 _31922_ (.A1(_09434_),
    .A2(_09435_),
    .A3(_09440_),
    .A4(_09441_),
    .ZN(_09442_));
 NOR2_X4 _31923_ (.A1(_09266_),
    .A2(_09267_),
    .ZN(_09443_));
 NAND4_X4 _31924_ (.A1(_09258_),
    .A2(_09283_),
    .A3(_09289_),
    .A4(_09351_),
    .ZN(_09444_));
 NOR2_X2 _31925_ (.A1(_09443_),
    .A2(_09444_),
    .ZN(_09445_));
 NOR4_X4 _31926_ (.A1(_09366_),
    .A2(_09368_),
    .A3(_09394_),
    .A4(_09396_),
    .ZN(_09446_));
 NAND3_X2 _31927_ (.A1(_09439_),
    .A2(_09445_),
    .A3(_09446_),
    .ZN(_09447_));
 NOR2_X4 _31928_ (.A1(_09300_),
    .A2(_09302_),
    .ZN(_09448_));
 AOI221_X2 _31929_ (.A(_09316_),
    .B1(_09274_),
    .B2(_09281_),
    .C1(_06936_),
    .C2(_09377_),
    .ZN(_09449_));
 NOR4_X2 _31930_ (.A1(_09448_),
    .A2(_09392_),
    .A3(_09426_),
    .A4(_09449_),
    .ZN(_09450_));
 NAND2_X2 _31931_ (.A1(_09378_),
    .A2(_09379_),
    .ZN(_09451_));
 NOR2_X4 _31932_ (.A1(_09451_),
    .A2(_09402_),
    .ZN(_09452_));
 OAI221_X2 _31933_ (.A(_09281_),
    .B1(_09300_),
    .B2(_09302_),
    .C1(_06934_),
    .C2(_00332_),
    .ZN(_09453_));
 BUF_X8 _31934_ (.A(_09453_),
    .Z(_09454_));
 NOR2_X4 _31935_ (.A1(_09454_),
    .A2(_09375_),
    .ZN(_09455_));
 NAND4_X2 _31936_ (.A1(_09283_),
    .A2(_09289_),
    .A3(_09348_),
    .A4(_09350_),
    .ZN(_09456_));
 OAI221_X2 _31937_ (.A(_09237_),
    .B1(_09300_),
    .B2(_09302_),
    .C1(_06888_),
    .C2(_09229_),
    .ZN(_09457_));
 OAI22_X2 _31938_ (.A1(_09385_),
    .A2(_09456_),
    .B1(_09457_),
    .B2(_09443_),
    .ZN(_09458_));
 OR2_X4 _31939_ (.A1(_00338_),
    .A2(_06886_),
    .ZN(_09459_));
 NAND2_X1 _31940_ (.A1(_09258_),
    .A2(_09459_),
    .ZN(_09460_));
 AND2_X1 _31941_ (.A1(_09460_),
    .A2(_09449_),
    .ZN(_09461_));
 AOI221_X2 _31942_ (.A(_09450_),
    .B1(_09452_),
    .B2(_09455_),
    .C1(_09458_),
    .C2(_09461_),
    .ZN(_09462_));
 NAND4_X4 _31943_ (.A1(_09430_),
    .A2(_09442_),
    .A3(_09447_),
    .A4(_09462_),
    .ZN(_09463_));
 BUF_X4 _31944_ (.A(_09432_),
    .Z(_09464_));
 NOR4_X1 _31945_ (.A1(_09412_),
    .A2(_09464_),
    .A3(_09343_),
    .A4(_09423_),
    .ZN(_09465_));
 NOR2_X4 _31946_ (.A1(_09394_),
    .A2(_09396_),
    .ZN(_09466_));
 NOR4_X2 _31947_ (.A1(_09437_),
    .A2(_09466_),
    .A3(_09305_),
    .A4(_09423_),
    .ZN(_09467_));
 OAI21_X2 _31948_ (.A(_09337_),
    .B1(_09465_),
    .B2(_09467_),
    .ZN(_09468_));
 OAI221_X2 _31949_ (.A(_09249_),
    .B1(_09309_),
    .B2(_09317_),
    .C1(_07486_),
    .C2(_09238_),
    .ZN(_09469_));
 OAI33_X1 _31950_ (.A1(_09466_),
    .A2(_09304_),
    .A3(_09375_),
    .B1(_09469_),
    .B2(_09360_),
    .B3(_09454_),
    .ZN(_09470_));
 NOR4_X4 _31951_ (.A1(_09394_),
    .A2(_09396_),
    .A3(_09309_),
    .A4(_09317_),
    .ZN(_09471_));
 BUF_X4 _31952_ (.A(_09451_),
    .Z(_09472_));
 NOR2_X4 _31953_ (.A1(_09466_),
    .A2(_09472_),
    .ZN(_09473_));
 NOR2_X4 _31954_ (.A1(_09271_),
    .A2(_09432_),
    .ZN(_09474_));
 AOI221_X2 _31955_ (.A(_09470_),
    .B1(_09471_),
    .B2(_09373_),
    .C1(_09473_),
    .C2(_09474_),
    .ZN(_09475_));
 BUF_X4 _31956_ (.A(_09412_),
    .Z(_09476_));
 OAI21_X2 _31957_ (.A(_09468_),
    .B1(_09475_),
    .B2(_09476_),
    .ZN(_09477_));
 NOR4_X2 _31958_ (.A1(_09392_),
    .A2(_09290_),
    .A3(_09426_),
    .A4(_09421_),
    .ZN(_09478_));
 NOR2_X4 _31959_ (.A1(_09336_),
    .A2(_09344_),
    .ZN(_09479_));
 NOR2_X2 _31960_ (.A1(_09454_),
    .A2(_09391_),
    .ZN(_09480_));
 NOR2_X1 _31961_ (.A1(_09448_),
    .A2(_09375_),
    .ZN(_09481_));
 AOI221_X2 _31962_ (.A(_09478_),
    .B1(_09479_),
    .B2(_09480_),
    .C1(_09387_),
    .C2(_09481_),
    .ZN(_09482_));
 OAI22_X2 _31963_ (.A1(_09271_),
    .A2(_09304_),
    .B1(_09432_),
    .B2(_09392_),
    .ZN(_09483_));
 NOR2_X4 _31964_ (.A1(_09375_),
    .A2(_09432_),
    .ZN(_09484_));
 OAI22_X4 _31965_ (.A1(_09309_),
    .A2(_09317_),
    .B1(_09320_),
    .B2(_09328_),
    .ZN(_09485_));
 NOR2_X2 _31966_ (.A1(_09436_),
    .A2(_09485_),
    .ZN(_09486_));
 NOR2_X4 _31967_ (.A1(_09436_),
    .A2(_09332_),
    .ZN(_09487_));
 NOR2_X4 _31968_ (.A1(_09303_),
    .A2(_09391_),
    .ZN(_09488_));
 AOI222_X2 _31969_ (.A1(_09437_),
    .A2(_09483_),
    .B1(_09484_),
    .B2(_09486_),
    .C1(_09487_),
    .C2(_09488_),
    .ZN(_09489_));
 BUF_X4 _31970_ (.A(_09466_),
    .Z(_09490_));
 BUF_X4 _31971_ (.A(_09490_),
    .Z(_09491_));
 BUF_X4 _31972_ (.A(_09437_),
    .Z(_09492_));
 OAI21_X1 _31973_ (.A(_09471_),
    .B1(_09291_),
    .B2(_09272_),
    .ZN(_09493_));
 OAI221_X2 _31974_ (.A(_09493_),
    .B1(_09469_),
    .B2(_09376_),
    .C1(_09490_),
    .C2(_09474_),
    .ZN(_09494_));
 OAI221_X2 _31975_ (.A(_09482_),
    .B1(_09489_),
    .B2(_09491_),
    .C1(_09492_),
    .C2(_09494_),
    .ZN(_09495_));
 OR4_X4 _31976_ (.A1(_09420_),
    .A2(_09463_),
    .A3(_09477_),
    .A4(_09495_),
    .ZN(_09496_));
 OAI221_X2 _31977_ (.A(_09341_),
    .B1(_09317_),
    .B2(_09309_),
    .C1(_09319_),
    .C2(_07486_),
    .ZN(_09497_));
 BUF_X8 _31978_ (.A(_09497_),
    .Z(_09498_));
 NOR2_X4 _31979_ (.A1(_09498_),
    .A2(_09398_),
    .ZN(_09499_));
 NOR3_X4 _31980_ (.A1(_09390_),
    .A2(_09454_),
    .A3(_09392_),
    .ZN(_09500_));
 NOR4_X4 _31981_ (.A1(_09366_),
    .A2(_09368_),
    .A3(_09309_),
    .A4(_09317_),
    .ZN(_09501_));
 NOR2_X4 _31982_ (.A1(_09498_),
    .A2(_09426_),
    .ZN(_09502_));
 AOI222_X2 _31983_ (.A1(_09484_),
    .A2(_09499_),
    .B1(_09500_),
    .B2(_09501_),
    .C1(_09502_),
    .C2(_09373_),
    .ZN(_09503_));
 BUF_X4 _31984_ (.A(_09472_),
    .Z(_09504_));
 NOR3_X4 _31985_ (.A1(_09272_),
    .A2(_09304_),
    .A3(_09333_),
    .ZN(_09505_));
 BUF_X4 _31986_ (.A(_09437_),
    .Z(_09506_));
 NOR3_X1 _31987_ (.A1(_09506_),
    .A2(_09305_),
    .A3(_09423_),
    .ZN(_09507_));
 OAI221_X2 _31988_ (.A(_09504_),
    .B1(_09505_),
    .B2(_09507_),
    .C1(_09334_),
    .C2(_09490_),
    .ZN(_09508_));
 NOR4_X4 _31989_ (.A1(_09360_),
    .A2(_09290_),
    .A3(_09498_),
    .A4(_09345_),
    .ZN(_09509_));
 NOR4_X4 _31990_ (.A1(_09466_),
    .A2(_09454_),
    .A3(_09375_),
    .A4(_09369_),
    .ZN(_09510_));
 NOR4_X2 _31991_ (.A1(_09305_),
    .A2(_09406_),
    .A3(_09498_),
    .A4(_09398_),
    .ZN(_09511_));
 NOR4_X2 _31992_ (.A1(_09472_),
    .A2(_09272_),
    .A3(_09433_),
    .A4(_09426_),
    .ZN(_09512_));
 NOR4_X4 _31993_ (.A1(_09509_),
    .A2(_09510_),
    .A3(_09511_),
    .A4(_09512_),
    .ZN(_09513_));
 NOR3_X2 _31994_ (.A1(_09412_),
    .A2(_09294_),
    .A3(_09291_),
    .ZN(_09514_));
 BUF_X4 _31995_ (.A(_09454_),
    .Z(_09515_));
 NOR4_X2 _31996_ (.A1(_09506_),
    .A2(_09515_),
    .A3(_09406_),
    .A4(_09343_),
    .ZN(_09516_));
 OAI21_X2 _31997_ (.A(_09473_),
    .B1(_09514_),
    .B2(_09516_),
    .ZN(_09517_));
 NAND4_X4 _31998_ (.A1(_09503_),
    .A2(_09508_),
    .A3(_09513_),
    .A4(_09517_),
    .ZN(_09518_));
 OAI21_X1 _31999_ (.A(_09472_),
    .B1(_09272_),
    .B2(_09433_),
    .ZN(_09519_));
 OAI221_X2 _32000_ (.A(_09250_),
    .B1(_09405_),
    .B2(_09519_),
    .C1(_09484_),
    .C2(_09504_),
    .ZN(_09520_));
 NOR2_X1 _32001_ (.A1(_09490_),
    .A2(_09485_),
    .ZN(_09521_));
 AOI21_X1 _32002_ (.A(_09483_),
    .B1(_09292_),
    .B2(_09521_),
    .ZN(_09522_));
 AOI221_X2 _32003_ (.A(_09298_),
    .B1(_09283_),
    .B2(_09289_),
    .C1(_07109_),
    .C2(_09273_),
    .ZN(_09523_));
 BUF_X4 _32004_ (.A(_09523_),
    .Z(_09524_));
 NOR3_X1 _32005_ (.A1(_09412_),
    .A2(_09472_),
    .A3(_09424_),
    .ZN(_09525_));
 OAI221_X2 _32006_ (.A(_09237_),
    .B1(_09309_),
    .B2(_09316_),
    .C1(_07486_),
    .C2(_09229_),
    .ZN(_09526_));
 NOR2_X1 _32007_ (.A1(_09406_),
    .A2(_09526_),
    .ZN(_09527_));
 OAI21_X1 _32008_ (.A(_09524_),
    .B1(_09525_),
    .B2(_09527_),
    .ZN(_09528_));
 OAI221_X2 _32009_ (.A(_09520_),
    .B1(_09522_),
    .B2(_09492_),
    .C1(_09528_),
    .C2(_09491_),
    .ZN(_09529_));
 NAND4_X4 _32010_ (.A1(_09239_),
    .A2(_09249_),
    .A3(_09274_),
    .A4(_09281_),
    .ZN(_09530_));
 NOR4_X2 _32011_ (.A1(_09443_),
    .A2(_09444_),
    .A3(_09526_),
    .A4(_09530_),
    .ZN(_09531_));
 OAI22_X4 _32012_ (.A1(_09394_),
    .A2(_09396_),
    .B1(_09309_),
    .B2(_09317_),
    .ZN(_09532_));
 OAI222_X2 _32013_ (.A1(_09366_),
    .A2(_09368_),
    .B1(_09296_),
    .B2(_09298_),
    .C1(_09300_),
    .C2(_09302_),
    .ZN(_09533_));
 OAI33_X1 _32014_ (.A1(_09385_),
    .A2(_09454_),
    .A3(_09271_),
    .B1(_09532_),
    .B2(_09533_),
    .B3(_09360_),
    .ZN(_09534_));
 NOR2_X4 _32015_ (.A1(_09357_),
    .A2(_09356_),
    .ZN(_09535_));
 OAI221_X2 _32016_ (.A(_09289_),
    .B1(_09266_),
    .B2(_09267_),
    .C1(_07486_),
    .C2(_09299_),
    .ZN(_09536_));
 NOR3_X1 _32017_ (.A1(_09385_),
    .A2(_09535_),
    .A3(_09536_),
    .ZN(_09537_));
 MUX2_X1 _32018_ (.A(_09471_),
    .B(_09410_),
    .S(_09438_),
    .Z(_09538_));
 AOI211_X2 _32019_ (.A(_09531_),
    .B(_09534_),
    .C1(_09537_),
    .C2(_09538_),
    .ZN(_09539_));
 OAI33_X1 _32020_ (.A1(_09439_),
    .A2(_09392_),
    .A3(_09398_),
    .B1(_09426_),
    .B2(_09303_),
    .B3(_09360_),
    .ZN(_09540_));
 NOR2_X2 _32021_ (.A1(_09345_),
    .A2(_09329_),
    .ZN(_09541_));
 NOR2_X4 _32022_ (.A1(_09392_),
    .A2(_09290_),
    .ZN(_09542_));
 BUF_X4 _32023_ (.A(_09480_),
    .Z(_09543_));
 AOI221_X2 _32024_ (.A(_09540_),
    .B1(_09541_),
    .B2(_09542_),
    .C1(_09403_),
    .C2(_09543_),
    .ZN(_09544_));
 NOR3_X2 _32025_ (.A1(_09412_),
    .A2(_09361_),
    .A3(_09305_),
    .ZN(_09545_));
 NOR3_X1 _32026_ (.A1(_09437_),
    .A2(_09406_),
    .A3(_09464_),
    .ZN(_09546_));
 OAI21_X2 _32027_ (.A(_09337_),
    .B1(_09545_),
    .B2(_09546_),
    .ZN(_09547_));
 NAND3_X2 _32028_ (.A1(_09539_),
    .A2(_09544_),
    .A3(_09547_),
    .ZN(_09548_));
 NOR2_X4 _32029_ (.A1(_09472_),
    .A2(_09426_),
    .ZN(_09549_));
 NOR2_X4 _32030_ (.A1(_09454_),
    .A2(_09361_),
    .ZN(_09550_));
 OAI21_X2 _32031_ (.A(_09549_),
    .B1(_09488_),
    .B2(_09550_),
    .ZN(_09551_));
 NOR2_X4 _32032_ (.A1(_09437_),
    .A2(_09466_),
    .ZN(_09552_));
 NAND3_X2 _32033_ (.A1(_09485_),
    .A2(_09292_),
    .A3(_09552_),
    .ZN(_09553_));
 NOR3_X4 _32034_ (.A1(_09392_),
    .A2(_09402_),
    .A3(_09290_),
    .ZN(_09554_));
 NOR2_X4 _32035_ (.A1(_09398_),
    .A2(_09421_),
    .ZN(_09555_));
 NOR2_X1 _32036_ (.A1(_09426_),
    .A2(_09449_),
    .ZN(_09556_));
 AOI221_X2 _32037_ (.A(_09554_),
    .B1(_09555_),
    .B2(_09455_),
    .C1(_09445_),
    .C2(_09556_),
    .ZN(_09557_));
 OAI221_X2 _32038_ (.A(_09348_),
    .B1(_09302_),
    .B2(_09300_),
    .C1(_09358_),
    .C2(_06887_),
    .ZN(_09558_));
 AOI221_X2 _32039_ (.A(_09438_),
    .B1(_09558_),
    .B2(_09536_),
    .C1(_09459_),
    .C2(_09258_),
    .ZN(_09559_));
 NOR2_X4 _32040_ (.A1(_09296_),
    .A2(_09298_),
    .ZN(_09560_));
 OAI21_X1 _32041_ (.A(_09369_),
    .B1(_09501_),
    .B2(_09560_),
    .ZN(_09561_));
 NOR3_X1 _32042_ (.A1(_09390_),
    .A2(_09535_),
    .A3(_09536_),
    .ZN(_09562_));
 OAI21_X1 _32043_ (.A(_09361_),
    .B1(_09272_),
    .B2(_09439_),
    .ZN(_09563_));
 NOR4_X4 _32044_ (.A1(_09296_),
    .A2(_09298_),
    .A3(_09300_),
    .A4(_09302_),
    .ZN(_09564_));
 NOR2_X1 _32045_ (.A1(_09437_),
    .A2(_09564_),
    .ZN(_09565_));
 AOI222_X2 _32046_ (.A1(_09250_),
    .A2(_09559_),
    .B1(_09561_),
    .B2(_09562_),
    .C1(_09563_),
    .C2(_09565_),
    .ZN(_09566_));
 NAND4_X4 _32047_ (.A1(_09551_),
    .A2(_09553_),
    .A3(_09557_),
    .A4(_09566_),
    .ZN(_09567_));
 OR4_X4 _32048_ (.A1(_09518_),
    .A2(_09529_),
    .A3(_09548_),
    .A4(_09567_),
    .ZN(_09568_));
 OAI21_X4 _32049_ (.A(_09389_),
    .B1(_09496_),
    .B2(_09568_),
    .ZN(_09569_));
 BUF_X4 _32050_ (.A(_09492_),
    .Z(_09570_));
 OAI21_X2 _32051_ (.A(_09482_),
    .B1(_09494_),
    .B2(_09570_),
    .ZN(_09571_));
 CLKBUF_X3 _32052_ (.A(_09343_),
    .Z(_09572_));
 NAND2_X4 _32053_ (.A1(_09258_),
    .A2(_09351_),
    .ZN(_09573_));
 NAND2_X2 _32054_ (.A1(_09348_),
    .A2(_09350_),
    .ZN(_09574_));
 OAI33_X1 _32055_ (.A1(_09515_),
    .A2(_09364_),
    .A3(_09572_),
    .B1(_09408_),
    .B2(_09573_),
    .B3(_09574_),
    .ZN(_09575_));
 AOI22_X4 _32056_ (.A1(_09488_),
    .A2(_09452_),
    .B1(_09479_),
    .B2(_09575_),
    .ZN(_09576_));
 NOR4_X1 _32057_ (.A1(_09413_),
    .A2(_09336_),
    .A3(_09424_),
    .A4(_09408_),
    .ZN(_09577_));
 AOI21_X2 _32058_ (.A(_09577_),
    .B1(_09487_),
    .B2(_09488_),
    .ZN(_09578_));
 BUF_X4 _32059_ (.A(_09415_),
    .Z(_09579_));
 BUF_X4 _32060_ (.A(_09579_),
    .Z(_09580_));
 AOI221_X2 _32061_ (.A(_09317_),
    .B1(_09340_),
    .B2(_09341_),
    .C1(_07109_),
    .C2(_09377_),
    .ZN(_09581_));
 BUF_X4 _32062_ (.A(_09581_),
    .Z(_09582_));
 CLKBUF_X3 _32063_ (.A(_09515_),
    .Z(_09583_));
 BUF_X4 _32064_ (.A(_09406_),
    .Z(_09584_));
 BUF_X4 _32065_ (.A(_09424_),
    .Z(_09585_));
 CLKBUF_X3 _32066_ (.A(_09408_),
    .Z(_09586_));
 OAI22_X1 _32067_ (.A1(_09583_),
    .A2(_09584_),
    .B1(_09585_),
    .B2(_09586_),
    .ZN(_09587_));
 AOI22_X2 _32068_ (.A1(_09582_),
    .A2(_09542_),
    .B1(_09587_),
    .B2(_09417_),
    .ZN(_09588_));
 BUF_X4 _32069_ (.A(_09402_),
    .Z(_09589_));
 OAI221_X2 _32070_ (.A(_09576_),
    .B1(_09578_),
    .B2(_09580_),
    .C1(_09588_),
    .C2(_09589_),
    .ZN(_09590_));
 NOR4_X4 _32071_ (.A1(_09466_),
    .A2(_09560_),
    .A3(_09361_),
    .A4(_09457_),
    .ZN(_09591_));
 BUF_X4 _32072_ (.A(_09498_),
    .Z(_09592_));
 AOI22_X2 _32073_ (.A1(_09550_),
    .A2(_09381_),
    .B1(_09591_),
    .B2(_09592_),
    .ZN(_09593_));
 BUF_X4 _32074_ (.A(_09472_),
    .Z(_09594_));
 NOR3_X1 _32075_ (.A1(_09464_),
    .A2(_09334_),
    .A3(_09424_),
    .ZN(_09595_));
 CLKBUF_X3 _32076_ (.A(_09464_),
    .Z(_09596_));
 NOR3_X1 _32077_ (.A1(_09407_),
    .A2(_09596_),
    .A3(_09572_),
    .ZN(_09597_));
 NOR3_X1 _32078_ (.A1(_09594_),
    .A2(_09595_),
    .A3(_09597_),
    .ZN(_09598_));
 BUF_X4 _32079_ (.A(_09484_),
    .Z(_09599_));
 NOR2_X2 _32080_ (.A1(_09433_),
    .A2(_09423_),
    .ZN(_09600_));
 BUF_X4 _32081_ (.A(_09600_),
    .Z(_09601_));
 OAI21_X1 _32082_ (.A(_09387_),
    .B1(_09599_),
    .B2(_09601_),
    .ZN(_09602_));
 NOR2_X4 _32083_ (.A1(_09515_),
    .A2(_09294_),
    .ZN(_09603_));
 NAND2_X2 _32084_ (.A1(_09383_),
    .A2(_09603_),
    .ZN(_09604_));
 NAND2_X2 _32085_ (.A1(_09338_),
    .A2(_09387_),
    .ZN(_09605_));
 OAI221_X2 _32086_ (.A(_09593_),
    .B1(_09598_),
    .B2(_09602_),
    .C1(_09604_),
    .C2(_09605_),
    .ZN(_09606_));
 NOR3_X1 _32087_ (.A1(_09407_),
    .A2(_09464_),
    .A3(_09380_),
    .ZN(_09607_));
 NOR4_X1 _32088_ (.A1(_09306_),
    .A2(_09406_),
    .A3(_09343_),
    .A4(_09369_),
    .ZN(_09608_));
 OAI21_X1 _32089_ (.A(_09579_),
    .B1(_09607_),
    .B2(_09608_),
    .ZN(_09609_));
 NAND2_X4 _32090_ (.A1(_09283_),
    .A2(_09289_),
    .ZN(_09610_));
 NOR2_X1 _32091_ (.A1(_09610_),
    .A2(_09424_),
    .ZN(_09611_));
 BUF_X4 _32092_ (.A(_09399_),
    .Z(_09612_));
 NOR2_X4 _32093_ (.A1(_09427_),
    .A2(_09612_),
    .ZN(_09613_));
 AOI22_X2 _32094_ (.A1(_09611_),
    .A2(_09555_),
    .B1(_09543_),
    .B2(_09613_),
    .ZN(_09614_));
 NAND2_X1 _32095_ (.A1(_09609_),
    .A2(_09614_),
    .ZN(_09615_));
 NOR4_X2 _32096_ (.A1(_09571_),
    .A2(_09590_),
    .A3(_09606_),
    .A4(_09615_),
    .ZN(_09616_));
 NOR3_X2 _32097_ (.A1(_09406_),
    .A2(_09433_),
    .A3(_09612_),
    .ZN(_09617_));
 OAI21_X1 _32098_ (.A(_09446_),
    .B1(_09505_),
    .B2(_09617_),
    .ZN(_09618_));
 NOR2_X4 _32099_ (.A1(_09402_),
    .A2(_09498_),
    .ZN(_09619_));
 MUX2_X1 _32100_ (.A(_09572_),
    .B(_09417_),
    .S(_09413_),
    .Z(_09620_));
 BUF_X4 _32101_ (.A(_09490_),
    .Z(_09621_));
 AOI21_X1 _32102_ (.A(_09619_),
    .B1(_09620_),
    .B2(_09621_),
    .ZN(_09622_));
 OR2_X2 _32103_ (.A1(_00335_),
    .A2(_06887_),
    .ZN(_09623_));
 AOI22_X4 _32104_ (.A1(_09258_),
    .A2(_09459_),
    .B1(_09348_),
    .B2(_09623_),
    .ZN(_09624_));
 NAND2_X2 _32105_ (.A1(_09624_),
    .A2(_09564_),
    .ZN(_09625_));
 BUF_X4 _32106_ (.A(_09455_),
    .Z(_09626_));
 NOR2_X1 _32107_ (.A1(_09492_),
    .A2(_09592_),
    .ZN(_09627_));
 MUX2_X1 _32108_ (.A(_09572_),
    .B(_09330_),
    .S(_09413_),
    .Z(_09628_));
 AOI22_X1 _32109_ (.A1(_09626_),
    .A2(_09627_),
    .B1(_09628_),
    .B2(_09405_),
    .ZN(_09629_));
 BUF_X4 _32110_ (.A(_09579_),
    .Z(_09630_));
 OAI221_X2 _32111_ (.A(_09618_),
    .B1(_09622_),
    .B2(_09625_),
    .C1(_09629_),
    .C2(_09630_),
    .ZN(_09631_));
 OAI21_X1 _32112_ (.A(_09580_),
    .B1(_09550_),
    .B2(_09601_),
    .ZN(_09632_));
 AOI21_X2 _32113_ (.A(_09370_),
    .B1(_09604_),
    .B2(_09632_),
    .ZN(_09633_));
 MUX2_X1 _32114_ (.A(_09583_),
    .B(_09596_),
    .S(_09492_),
    .Z(_09634_));
 AOI221_X2 _32115_ (.A(_09357_),
    .B1(_09348_),
    .B2(_09623_),
    .C1(_07109_),
    .C2(_09268_),
    .ZN(_09635_));
 NAND3_X2 _32116_ (.A1(_09621_),
    .A2(_09635_),
    .A3(_09592_),
    .ZN(_09636_));
 NOR3_X2 _32117_ (.A1(_09464_),
    .A2(_09343_),
    .A3(_09424_),
    .ZN(_09637_));
 AOI21_X2 _32118_ (.A(_09637_),
    .B1(_09626_),
    .B2(_09383_),
    .ZN(_09638_));
 NAND2_X2 _32119_ (.A1(_09337_),
    .A2(_09251_),
    .ZN(_09639_));
 OAI22_X4 _32120_ (.A1(_09634_),
    .A2(_09636_),
    .B1(_09638_),
    .B2(_09639_),
    .ZN(_09640_));
 NOR2_X4 _32121_ (.A1(_09361_),
    .A2(_09433_),
    .ZN(_09641_));
 AOI222_X2 _32122_ (.A1(_09455_),
    .A2(_09555_),
    .B1(_09641_),
    .B2(_09400_),
    .C1(_09452_),
    .C2(_09401_),
    .ZN(_09642_));
 NOR3_X1 _32123_ (.A1(_09407_),
    .A2(_09596_),
    .A3(_09371_),
    .ZN(_09643_));
 AOI21_X1 _32124_ (.A(_09643_),
    .B1(_09637_),
    .B2(_09579_),
    .ZN(_09644_));
 NAND3_X1 _32125_ (.A1(_09560_),
    .A2(_09353_),
    .A3(_09552_),
    .ZN(_09645_));
 NOR2_X1 _32126_ (.A1(_09448_),
    .A2(_09334_),
    .ZN(_09646_));
 XNOR2_X1 _32127_ (.A(_09594_),
    .B(_09646_),
    .ZN(_09647_));
 OAI221_X2 _32128_ (.A(_09642_),
    .B1(_09644_),
    .B2(_09526_),
    .C1(_09645_),
    .C2(_09647_),
    .ZN(_09648_));
 NOR4_X4 _32129_ (.A1(_09631_),
    .A2(_09633_),
    .A3(_09640_),
    .A4(_09648_),
    .ZN(_09649_));
 BUF_X4 _32130_ (.A(_09474_),
    .Z(_09650_));
 AOI22_X4 _32131_ (.A1(_09378_),
    .A2(_09379_),
    .B1(_09340_),
    .B2(_09341_),
    .ZN(_09651_));
 AOI22_X2 _32132_ (.A1(_09650_),
    .A2(_09651_),
    .B1(_09330_),
    .B2(_09374_),
    .ZN(_09652_));
 NOR2_X2 _32133_ (.A1(_09345_),
    .A2(_09652_),
    .ZN(_09653_));
 NOR2_X1 _32134_ (.A1(_09334_),
    .A2(_09589_),
    .ZN(_09654_));
 OAI21_X1 _32135_ (.A(_09654_),
    .B1(_09405_),
    .B2(_09599_),
    .ZN(_09655_));
 OAI21_X1 _32136_ (.A(_09400_),
    .B1(_09292_),
    .B2(_09376_),
    .ZN(_09656_));
 NOR4_X2 _32137_ (.A1(_09437_),
    .A2(_09360_),
    .A3(_09290_),
    .A4(_09416_),
    .ZN(_09657_));
 AOI221_X2 _32138_ (.A(_09509_),
    .B1(_09619_),
    .B2(_09474_),
    .C1(_09657_),
    .C2(_09390_),
    .ZN(_09658_));
 NAND3_X2 _32139_ (.A1(_09655_),
    .A2(_09656_),
    .A3(_09658_),
    .ZN(_09659_));
 BUF_X4 _32140_ (.A(_09413_),
    .Z(_09660_));
 NAND2_X1 _32141_ (.A1(_09524_),
    .A2(_09635_),
    .ZN(_09661_));
 NAND2_X1 _32142_ (.A1(_09601_),
    .A2(_09485_),
    .ZN(_09662_));
 OAI221_X2 _32143_ (.A(_09660_),
    .B1(_09532_),
    .B2(_09661_),
    .C1(_09662_),
    .C2(_09580_),
    .ZN(_09663_));
 BUF_X4 _32144_ (.A(_09506_),
    .Z(_09664_));
 AOI221_X2 _32145_ (.A(_09266_),
    .B1(_09459_),
    .B2(_09258_),
    .C1(_09349_),
    .C2(_07108_),
    .ZN(_09665_));
 NAND2_X1 _32146_ (.A1(_09665_),
    .A2(_09564_),
    .ZN(_09666_));
 AOI21_X1 _32147_ (.A(_09582_),
    .B1(_09592_),
    .B2(_09579_),
    .ZN(_09667_));
 OR2_X2 _32148_ (.A1(_09361_),
    .A2(_09464_),
    .ZN(_09668_));
 OAI221_X2 _32149_ (.A(_09664_),
    .B1(_09666_),
    .B2(_09532_),
    .C1(_09667_),
    .C2(_09668_),
    .ZN(_09669_));
 AOI211_X2 _32150_ (.A(_09653_),
    .B(_09659_),
    .C1(_09663_),
    .C2(_09669_),
    .ZN(_09670_));
 BUF_X4 _32151_ (.A(_09333_),
    .Z(_09671_));
 NOR4_X1 _32152_ (.A1(_09337_),
    .A2(_09307_),
    .A3(_09671_),
    .A4(_09585_),
    .ZN(_09672_));
 CLKBUF_X3 _32153_ (.A(_09364_),
    .Z(_09673_));
 NOR3_X1 _32154_ (.A1(_09673_),
    .A2(_09307_),
    .A3(_09612_),
    .ZN(_09674_));
 OAI21_X1 _32155_ (.A(_09251_),
    .B1(_09672_),
    .B2(_09674_),
    .ZN(_09675_));
 AOI222_X2 _32156_ (.A1(_09650_),
    .A2(_09381_),
    .B1(_09372_),
    .B2(_09543_),
    .C1(_09613_),
    .C2(_09488_),
    .ZN(_09676_));
 NOR3_X1 _32157_ (.A1(_09307_),
    .A2(_09585_),
    .A3(_09592_),
    .ZN(_09677_));
 OAI21_X1 _32158_ (.A(_09552_),
    .B1(_09505_),
    .B2(_09677_),
    .ZN(_09678_));
 AND3_X1 _32159_ (.A1(_09675_),
    .A2(_09676_),
    .A3(_09678_),
    .ZN(_09679_));
 NAND4_X4 _32160_ (.A1(_09616_),
    .A2(_09649_),
    .A3(_09670_),
    .A4(_09679_),
    .ZN(_09680_));
 OR2_X4 _32161_ (.A1(_09569_),
    .A2(_09680_),
    .ZN(_09681_));
 NAND2_X2 _32162_ (.A1(_07260_),
    .A2(_09681_),
    .ZN(_09682_));
 NOR2_X1 _32163_ (.A1(_07234_),
    .A2(_08722_),
    .ZN(_09683_));
 XNOR2_X1 _32164_ (.A(_07239_),
    .B(_08166_),
    .ZN(_09684_));
 XNOR2_X1 _32165_ (.A(_00361_),
    .B(_09684_),
    .ZN(_09685_));
 AOI21_X2 _32166_ (.A(_09683_),
    .B1(_09685_),
    .B2(_09217_),
    .ZN(_09686_));
 OAI221_X2 _32167_ (.A(_04262_),
    .B1(_09223_),
    .B2(_09686_),
    .C1(_09221_),
    .C2(\block_reg[0][24] ),
    .ZN(_09687_));
 NAND2_X1 _32168_ (.A1(_07908_),
    .A2(_09686_),
    .ZN(_09688_));
 INV_X1 _32169_ (.A(\block_reg[0][24] ),
    .ZN(_09689_));
 OAI21_X1 _32170_ (.A(_09688_),
    .B1(_07787_),
    .B2(_09689_),
    .ZN(_09690_));
 OR2_X1 _32171_ (.A1(_04262_),
    .A2(_09690_),
    .ZN(_09691_));
 AOI21_X2 _32172_ (.A(_06704_),
    .B1(_09687_),
    .B2(_09691_),
    .ZN(_09692_));
 AOI22_X1 _32173_ (.A1(_09228_),
    .A2(_07661_),
    .B1(_09682_),
    .B2(_09692_),
    .ZN(_00718_));
 INV_X1 _32174_ (.A(_08999_),
    .ZN(_09693_));
 NOR4_X1 _32175_ (.A1(_09673_),
    .A2(_09596_),
    .A3(_09671_),
    .A4(_09427_),
    .ZN(_09694_));
 OAI22_X1 _32176_ (.A1(_09583_),
    .A2(_09295_),
    .B1(_09596_),
    .B2(_09673_),
    .ZN(_09695_));
 AOI21_X2 _32177_ (.A(_09694_),
    .B1(_09695_),
    .B2(_09549_),
    .ZN(_09696_));
 NOR3_X1 _32178_ (.A1(_09584_),
    .A2(_09586_),
    .A3(_09612_),
    .ZN(_09697_));
 OAI21_X2 _32179_ (.A(_09251_),
    .B1(_09331_),
    .B2(_09697_),
    .ZN(_09698_));
 NOR3_X1 _32180_ (.A1(_09307_),
    .A2(_09671_),
    .A3(_09585_),
    .ZN(_09699_));
 NOR3_X1 _32181_ (.A1(_09673_),
    .A2(_09383_),
    .A3(_09586_),
    .ZN(_09700_));
 NOR3_X2 _32182_ (.A1(_09580_),
    .A2(_09699_),
    .A3(_09700_),
    .ZN(_09701_));
 NOR2_X4 _32183_ (.A1(_09385_),
    .A2(_09336_),
    .ZN(_09702_));
 NOR3_X1 _32184_ (.A1(_09673_),
    .A2(_09671_),
    .A3(_09586_),
    .ZN(_09703_));
 OAI21_X2 _32185_ (.A(_09702_),
    .B1(_09703_),
    .B2(_09621_),
    .ZN(_09704_));
 OAI211_X4 _32186_ (.A(_09696_),
    .B(_09698_),
    .C1(_09701_),
    .C2(_09704_),
    .ZN(_09705_));
 NOR4_X4 _32187_ (.A1(_09420_),
    .A2(_09463_),
    .A3(_09477_),
    .A4(_09495_),
    .ZN(_09706_));
 NOR4_X4 _32188_ (.A1(_09518_),
    .A2(_09529_),
    .A3(_09548_),
    .A4(_09567_),
    .ZN(_09707_));
 AOI21_X4 _32189_ (.A(_09705_),
    .B1(_09706_),
    .B2(_09707_),
    .ZN(_09708_));
 BUF_X4 _32190_ (.A(_09398_),
    .Z(_09709_));
 NOR2_X2 _32191_ (.A1(_09336_),
    .A2(_09709_),
    .ZN(_09710_));
 AOI222_X2 _32192_ (.A1(_09599_),
    .A2(_09502_),
    .B1(_09710_),
    .B2(_09455_),
    .C1(_09499_),
    .C2(_09543_),
    .ZN(_09711_));
 AOI22_X4 _32193_ (.A1(_09446_),
    .A2(_09362_),
    .B1(_09452_),
    .B2(_09626_),
    .ZN(_09712_));
 OAI21_X2 _32194_ (.A(_09711_),
    .B1(_09712_),
    .B2(_09384_),
    .ZN(_09713_));
 AOI22_X4 _32195_ (.A1(_09641_),
    .A2(_09479_),
    .B1(_09619_),
    .B2(_09293_),
    .ZN(_09714_));
 AOI222_X2 _32196_ (.A1(_09550_),
    .A2(_09251_),
    .B1(_09543_),
    .B2(_09400_),
    .C1(_09549_),
    .C2(_09484_),
    .ZN(_09715_));
 NOR2_X1 _32197_ (.A1(_09415_),
    .A2(_09485_),
    .ZN(_09716_));
 AOI22_X4 _32198_ (.A1(_09626_),
    .A2(_09381_),
    .B1(_09716_),
    .B2(_09401_),
    .ZN(_09717_));
 NAND3_X4 _32199_ (.A1(_09714_),
    .A2(_09715_),
    .A3(_09717_),
    .ZN(_09718_));
 NOR2_X2 _32200_ (.A1(_09466_),
    .A2(_09333_),
    .ZN(_09719_));
 NAND2_X1 _32201_ (.A1(_09524_),
    .A2(_09353_),
    .ZN(_09720_));
 NOR2_X1 _32202_ (.A1(_09358_),
    .A2(_06888_),
    .ZN(_09721_));
 NOR2_X1 _32203_ (.A1(_09266_),
    .A2(_09721_),
    .ZN(_09722_));
 NAND2_X1 _32204_ (.A1(_09348_),
    .A2(_09623_),
    .ZN(_09723_));
 MUX2_X1 _32205_ (.A(_09722_),
    .B(_09723_),
    .S(_09439_),
    .Z(_09724_));
 NOR3_X1 _32206_ (.A1(_09472_),
    .A2(_09535_),
    .A3(_09448_),
    .ZN(_09725_));
 AOI22_X1 _32207_ (.A1(_09611_),
    .A2(_09485_),
    .B1(_09724_),
    .B2(_09725_),
    .ZN(_09726_));
 OAI33_X1 _32208_ (.A1(_09370_),
    .A2(_09719_),
    .A3(_09720_),
    .B1(_09726_),
    .B2(_09492_),
    .B3(_09491_),
    .ZN(_09727_));
 AOI221_X2 _32209_ (.A(_09437_),
    .B1(_09274_),
    .B2(_09281_),
    .C1(_09610_),
    .C2(_09472_),
    .ZN(_09728_));
 NOR3_X1 _32210_ (.A1(_09490_),
    .A2(_09294_),
    .A3(_09572_),
    .ZN(_09729_));
 NOR2_X1 _32211_ (.A1(_09294_),
    .A2(_09371_),
    .ZN(_09730_));
 AND3_X1 _32212_ (.A1(_09506_),
    .A2(_09610_),
    .A3(_09449_),
    .ZN(_09731_));
 AOI22_X2 _32213_ (.A1(_09728_),
    .A2(_09729_),
    .B1(_09730_),
    .B2(_09731_),
    .ZN(_09732_));
 NAND4_X2 _32214_ (.A1(_09551_),
    .A2(_09553_),
    .A3(_09557_),
    .A4(_09732_),
    .ZN(_09733_));
 NOR4_X2 _32215_ (.A1(_09713_),
    .A2(_09718_),
    .A3(_09727_),
    .A4(_09733_),
    .ZN(_09734_));
 OAI21_X2 _32216_ (.A(_09576_),
    .B1(_09578_),
    .B2(_09630_),
    .ZN(_09735_));
 OAI33_X1 _32217_ (.A1(_09574_),
    .A2(_09573_),
    .A3(_09596_),
    .B1(_09334_),
    .B2(_09407_),
    .B3(_09515_),
    .ZN(_09736_));
 NAND3_X1 _32218_ (.A1(_09446_),
    .A2(_09422_),
    .A3(_09736_),
    .ZN(_09737_));
 NOR4_X4 _32219_ (.A1(_09413_),
    .A2(_09448_),
    .A3(_09407_),
    .A4(_09530_),
    .ZN(_09738_));
 OAI21_X4 _32220_ (.A(_09417_),
    .B1(_09591_),
    .B2(_09738_),
    .ZN(_09739_));
 NAND2_X1 _32221_ (.A1(_09476_),
    .A2(_09383_),
    .ZN(_09740_));
 NAND2_X1 _32222_ (.A1(_09491_),
    .A2(_09671_),
    .ZN(_09741_));
 NOR3_X1 _32223_ (.A1(_09336_),
    .A2(_09306_),
    .A3(_09407_),
    .ZN(_09742_));
 NAND3_X1 _32224_ (.A1(_09740_),
    .A2(_09741_),
    .A3(_09742_),
    .ZN(_09743_));
 NAND4_X2 _32225_ (.A1(_09658_),
    .A2(_09737_),
    .A3(_09739_),
    .A4(_09743_),
    .ZN(_09744_));
 OR2_X2 _32226_ (.A1(_09272_),
    .A2(_09432_),
    .ZN(_09745_));
 NAND2_X2 _32227_ (.A1(_09665_),
    .A2(_09347_),
    .ZN(_09746_));
 OAI33_X1 _32228_ (.A1(_09506_),
    .A2(_09745_),
    .A3(_09330_),
    .B1(_09746_),
    .B2(_09333_),
    .B3(_09369_),
    .ZN(_09747_));
 AND2_X2 _32229_ (.A1(_09491_),
    .A2(_09747_),
    .ZN(_09748_));
 NAND2_X2 _32230_ (.A1(_09582_),
    .A2(_09545_),
    .ZN(_09749_));
 NOR2_X1 _32231_ (.A1(_09506_),
    .A2(_09612_),
    .ZN(_09750_));
 AOI22_X4 _32232_ (.A1(_09486_),
    .A2(_09292_),
    .B1(_09603_),
    .B2(_09750_),
    .ZN(_09751_));
 AOI21_X4 _32233_ (.A(_09580_),
    .B1(_09749_),
    .B2(_09751_),
    .ZN(_09752_));
 NOR4_X4 _32234_ (.A1(_09735_),
    .A2(_09744_),
    .A3(_09748_),
    .A4(_09752_),
    .ZN(_09753_));
 BUF_X4 _32235_ (.A(_09594_),
    .Z(_09754_));
 NOR4_X2 _32236_ (.A1(_09294_),
    .A2(_09333_),
    .A3(_09291_),
    .A4(_09345_),
    .ZN(_09755_));
 AOI221_X2 _32237_ (.A(_09755_),
    .B1(_09346_),
    .B2(_09401_),
    .C1(_09719_),
    .C2(_09514_),
    .ZN(_09756_));
 AOI221_X2 _32238_ (.A(_09617_),
    .B1(_09651_),
    .B2(_09484_),
    .C1(_09488_),
    .C2(_09417_),
    .ZN(_09757_));
 OAI22_X4 _32239_ (.A1(_09754_),
    .A2(_09756_),
    .B1(_09757_),
    .B2(_09589_),
    .ZN(_09758_));
 OAI221_X1 _32240_ (.A(_09579_),
    .B1(_09306_),
    .B2(_09585_),
    .C1(_09586_),
    .C2(_09584_),
    .ZN(_09759_));
 OAI21_X1 _32241_ (.A(_09491_),
    .B1(_09295_),
    .B2(_09306_),
    .ZN(_09760_));
 NAND3_X1 _32242_ (.A1(_09487_),
    .A2(_09759_),
    .A3(_09760_),
    .ZN(_09761_));
 NOR4_X1 _32243_ (.A1(_09579_),
    .A2(_09515_),
    .A3(_09294_),
    .A4(_09572_),
    .ZN(_09762_));
 NOR4_X2 _32244_ (.A1(_09491_),
    .A2(_09515_),
    .A3(_09407_),
    .A4(_09334_),
    .ZN(_09763_));
 OAI21_X2 _32245_ (.A(_09702_),
    .B1(_09762_),
    .B2(_09763_),
    .ZN(_09764_));
 NOR3_X1 _32246_ (.A1(_09584_),
    .A2(_09586_),
    .A3(_09532_),
    .ZN(_09765_));
 NOR4_X2 _32247_ (.A1(_09415_),
    .A2(_09364_),
    .A3(_09408_),
    .A4(_09422_),
    .ZN(_09766_));
 OAI21_X2 _32248_ (.A(_09664_),
    .B1(_09765_),
    .B2(_09766_),
    .ZN(_09767_));
 NAND4_X4 _32249_ (.A1(_09503_),
    .A2(_09761_),
    .A3(_09764_),
    .A4(_09767_),
    .ZN(_09768_));
 NOR2_X1 _32250_ (.A1(_09416_),
    .A2(_09582_),
    .ZN(_09769_));
 MUX2_X1 _32251_ (.A(_09746_),
    .B(_09661_),
    .S(_09769_),
    .Z(_09770_));
 NOR4_X2 _32252_ (.A1(_09390_),
    .A2(_09304_),
    .A3(_09423_),
    .A4(_09498_),
    .ZN(_09771_));
 NOR3_X4 _32253_ (.A1(_09454_),
    .A2(_09272_),
    .A3(_09332_),
    .ZN(_09772_));
 AOI221_X2 _32254_ (.A(_09771_),
    .B1(_09772_),
    .B2(_09410_),
    .C1(_09582_),
    .C2(_09641_),
    .ZN(_09773_));
 OAI22_X2 _32255_ (.A1(_09589_),
    .A2(_09770_),
    .B1(_09773_),
    .B2(_09570_),
    .ZN(_09774_));
 NOR3_X2 _32256_ (.A1(_09758_),
    .A2(_09768_),
    .A3(_09774_),
    .ZN(_09775_));
 AND3_X2 _32257_ (.A1(_09734_),
    .A2(_09753_),
    .A3(_09775_),
    .ZN(_09776_));
 NAND2_X4 _32258_ (.A1(_09708_),
    .A2(_09776_),
    .ZN(_09777_));
 NAND2_X2 _32259_ (.A1(_07662_),
    .A2(_09777_),
    .ZN(_09778_));
 XNOR2_X1 _32260_ (.A(_08187_),
    .B(_07645_),
    .ZN(_09779_));
 XNOR2_X1 _32261_ (.A(_07236_),
    .B(_09779_),
    .ZN(_09780_));
 XNOR2_X1 _32262_ (.A(_08718_),
    .B(_09780_),
    .ZN(_09781_));
 NAND2_X1 _32263_ (.A1(_08039_),
    .A2(_09781_),
    .ZN(_09782_));
 OAI21_X2 _32264_ (.A(_09782_),
    .B1(_08048_),
    .B2(_00343_),
    .ZN(_09783_));
 OAI22_X1 _32265_ (.A1(\block_reg[0][25] ),
    .A2(_07251_),
    .B1(_07254_),
    .B2(_09783_),
    .ZN(_09784_));
 NAND2_X1 _32266_ (.A1(_07229_),
    .A2(_09783_),
    .ZN(_09785_));
 OAI21_X1 _32267_ (.A(_09785_),
    .B1(_07248_),
    .B2(_04539_),
    .ZN(_09786_));
 MUX2_X1 _32268_ (.A(_09784_),
    .B(_09786_),
    .S(_04550_),
    .Z(_09787_));
 NOR2_X1 _32269_ (.A1(_07224_),
    .A2(_09787_),
    .ZN(_09788_));
 AOI22_X1 _32270_ (.A1(_09693_),
    .A2(_07661_),
    .B1(_09778_),
    .B2(_09788_),
    .ZN(_00719_));
 AOI221_X2 _32271_ (.A(_09491_),
    .B1(_09600_),
    .B2(_09702_),
    .C1(_09641_),
    .C2(_09337_),
    .ZN(_09789_));
 BUF_X4 _32272_ (.A(_09621_),
    .Z(_09790_));
 OAI21_X1 _32273_ (.A(_09519_),
    .B1(_09599_),
    .B2(_09594_),
    .ZN(_09791_));
 AOI21_X1 _32274_ (.A(_09742_),
    .B1(_09455_),
    .B2(_09337_),
    .ZN(_09792_));
 MUX2_X1 _32275_ (.A(_09791_),
    .B(_09792_),
    .S(_09660_),
    .Z(_09793_));
 AOI221_X2 _32276_ (.A(_09789_),
    .B1(_09341_),
    .B2(_09340_),
    .C1(_09790_),
    .C2(_09793_),
    .ZN(_09794_));
 OAI33_X1 _32277_ (.A1(_09476_),
    .A2(_09584_),
    .A3(_09586_),
    .B1(_09709_),
    .B2(_09294_),
    .B3(_09515_),
    .ZN(_09795_));
 NAND2_X1 _32278_ (.A1(_09582_),
    .A2(_09795_),
    .ZN(_09796_));
 XNOR2_X1 _32279_ (.A(_09412_),
    .B(_09504_),
    .ZN(_09797_));
 AOI22_X2 _32280_ (.A1(_09641_),
    .A2(_09710_),
    .B1(_09797_),
    .B2(_09500_),
    .ZN(_09798_));
 NAND2_X1 _32281_ (.A1(_09621_),
    .A2(_09401_),
    .ZN(_09799_));
 OAI221_X2 _32282_ (.A(_09796_),
    .B1(_09798_),
    .B2(_09335_),
    .C1(_09370_),
    .C2(_09799_),
    .ZN(_09800_));
 OAI21_X1 _32283_ (.A(_09542_),
    .B1(_09502_),
    .B2(_09452_),
    .ZN(_09801_));
 NOR2_X1 _32284_ (.A1(_09589_),
    .A2(_09417_),
    .ZN(_09802_));
 AOI222_X2 _32285_ (.A1(_09550_),
    .A2(_09549_),
    .B1(_09502_),
    .B2(_09292_),
    .C1(_09802_),
    .C2(_09599_),
    .ZN(_09803_));
 OAI21_X2 _32286_ (.A(_09384_),
    .B1(_09554_),
    .B2(_09365_),
    .ZN(_09804_));
 NAND4_X4 _32287_ (.A1(_09739_),
    .A2(_09801_),
    .A3(_09803_),
    .A4(_09804_),
    .ZN(_09805_));
 NAND3_X1 _32288_ (.A1(_09675_),
    .A2(_09676_),
    .A3(_09678_),
    .ZN(_09806_));
 OR2_X1 _32289_ (.A1(_09420_),
    .A2(_09806_),
    .ZN(_09807_));
 NOR4_X4 _32290_ (.A1(_09794_),
    .A2(_09800_),
    .A3(_09805_),
    .A4(_09807_),
    .ZN(_09808_));
 NOR3_X1 _32291_ (.A1(_09506_),
    .A2(_09294_),
    .A3(_09291_),
    .ZN(_09809_));
 OAI221_X2 _32292_ (.A(_09379_),
    .B1(_09396_),
    .B2(_09394_),
    .C1(_09308_),
    .C2(_06888_),
    .ZN(_09810_));
 OAI22_X1 _32293_ (.A1(_09810_),
    .A2(_09333_),
    .B1(_09498_),
    .B2(_09415_),
    .ZN(_09811_));
 AND2_X1 _32294_ (.A1(_09809_),
    .A2(_09811_),
    .ZN(_09812_));
 OAI22_X2 _32295_ (.A1(_09709_),
    .A2(_09668_),
    .B1(_09746_),
    .B2(_09413_),
    .ZN(_09813_));
 MUX2_X1 _32296_ (.A(_09600_),
    .B(_09455_),
    .S(_09572_),
    .Z(_09814_));
 AOI221_X2 _32297_ (.A(_09812_),
    .B1(_09813_),
    .B2(_09417_),
    .C1(_09549_),
    .C2(_09814_),
    .ZN(_09815_));
 AOI221_X2 _32298_ (.A(_09510_),
    .B1(_09362_),
    .B2(_09400_),
    .C1(_09381_),
    .C2(_09542_),
    .ZN(_09816_));
 OAI22_X1 _32299_ (.A1(_09448_),
    .A2(_09469_),
    .B1(_09810_),
    .B2(_09464_),
    .ZN(_09817_));
 NOR2_X1 _32300_ (.A1(_09492_),
    .A2(_09294_),
    .ZN(_09818_));
 AOI22_X1 _32301_ (.A1(_09650_),
    .A2(_09452_),
    .B1(_09817_),
    .B2(_09818_),
    .ZN(_09819_));
 OAI21_X2 _32302_ (.A(_09816_),
    .B1(_09819_),
    .B2(_09335_),
    .ZN(_09820_));
 OAI21_X1 _32303_ (.A(_09384_),
    .B1(_09488_),
    .B2(_09603_),
    .ZN(_09821_));
 NAND2_X1 _32304_ (.A1(_09524_),
    .A2(_09665_),
    .ZN(_09822_));
 AOI21_X1 _32305_ (.A(_09639_),
    .B1(_09821_),
    .B2(_09822_),
    .ZN(_09823_));
 NAND3_X1 _32306_ (.A1(_09660_),
    .A2(_09754_),
    .A3(_09559_),
    .ZN(_09824_));
 NAND3_X1 _32307_ (.A1(_09570_),
    .A2(_09650_),
    .A3(_09330_),
    .ZN(_09825_));
 AOI21_X1 _32308_ (.A(_09630_),
    .B1(_09824_),
    .B2(_09825_),
    .ZN(_09826_));
 NOR3_X1 _32309_ (.A1(_09820_),
    .A2(_09823_),
    .A3(_09826_),
    .ZN(_09827_));
 NOR3_X1 _32310_ (.A1(_09466_),
    .A2(_09454_),
    .A3(_09423_),
    .ZN(_09828_));
 NOR3_X1 _32311_ (.A1(_09390_),
    .A2(_09272_),
    .A3(_09304_),
    .ZN(_09829_));
 NOR3_X1 _32312_ (.A1(_09504_),
    .A2(_09828_),
    .A3(_09829_),
    .ZN(_09830_));
 NAND2_X1 _32313_ (.A1(_09333_),
    .A2(_09641_),
    .ZN(_09831_));
 AOI221_X2 _32314_ (.A(_09830_),
    .B1(_09831_),
    .B2(_09504_),
    .C1(_09230_),
    .C2(_09237_),
    .ZN(_09832_));
 NAND2_X2 _32315_ (.A1(_09579_),
    .A2(_09383_),
    .ZN(_09833_));
 NOR3_X1 _32316_ (.A1(_09650_),
    .A2(_09599_),
    .A3(_09542_),
    .ZN(_09834_));
 NOR3_X2 _32317_ (.A1(_09526_),
    .A2(_09833_),
    .A3(_09834_),
    .ZN(_09835_));
 NOR2_X1 _32318_ (.A1(_09412_),
    .A2(_09343_),
    .ZN(_09836_));
 AOI22_X2 _32319_ (.A1(_09476_),
    .A2(_09626_),
    .B1(_09603_),
    .B2(_09836_),
    .ZN(_09837_));
 OAI22_X2 _32320_ (.A1(_09589_),
    .A2(_09604_),
    .B1(_09837_),
    .B2(_09580_),
    .ZN(_09838_));
 AOI211_X2 _32321_ (.A(_09832_),
    .B(_09835_),
    .C1(_09754_),
    .C2(_09838_),
    .ZN(_09839_));
 OAI21_X1 _32322_ (.A(_09370_),
    .B1(_09612_),
    .B2(_09664_),
    .ZN(_09840_));
 AOI21_X1 _32323_ (.A(_09654_),
    .B1(_09840_),
    .B2(_09790_),
    .ZN(_09841_));
 INV_X1 _32324_ (.A(_09376_),
    .ZN(_09842_));
 OAI221_X2 _32325_ (.A(_09711_),
    .B1(_09841_),
    .B2(_09842_),
    .C1(_09384_),
    .C2(_09712_),
    .ZN(_09843_));
 OAI21_X1 _32326_ (.A(_09613_),
    .B1(_09362_),
    .B2(_09543_),
    .ZN(_09844_));
 OAI21_X1 _32327_ (.A(_09499_),
    .B1(_09542_),
    .B2(_09599_),
    .ZN(_09845_));
 AOI21_X1 _32328_ (.A(_09306_),
    .B1(_09585_),
    .B2(_09673_),
    .ZN(_09846_));
 AOI222_X2 _32329_ (.A1(_09601_),
    .A2(_09552_),
    .B1(_09555_),
    .B2(_09846_),
    .C1(_09372_),
    .C2(_09550_),
    .ZN(_09847_));
 AOI22_X1 _32330_ (.A1(_09505_),
    .A2(_09452_),
    .B1(_09619_),
    .B2(_09650_),
    .ZN(_09848_));
 NAND4_X1 _32331_ (.A1(_09844_),
    .A2(_09845_),
    .A3(_09847_),
    .A4(_09848_),
    .ZN(_09849_));
 NOR2_X1 _32332_ (.A1(_09664_),
    .A2(_09417_),
    .ZN(_09850_));
 OAI21_X1 _32333_ (.A(_09422_),
    .B1(_09592_),
    .B2(_09476_),
    .ZN(_09851_));
 OAI21_X1 _32334_ (.A(_09601_),
    .B1(_09850_),
    .B2(_09851_),
    .ZN(_09852_));
 AOI21_X1 _32335_ (.A(_09630_),
    .B1(_09749_),
    .B2(_09852_),
    .ZN(_09853_));
 NAND2_X1 _32336_ (.A1(_09353_),
    .A2(_09564_),
    .ZN(_09854_));
 OAI33_X1 _32337_ (.A1(_09307_),
    .A2(_09584_),
    .A3(_09810_),
    .B1(_09383_),
    .B2(_09854_),
    .B3(_09469_),
    .ZN(_09855_));
 AND2_X1 _32338_ (.A1(_09660_),
    .A2(_09855_),
    .ZN(_09856_));
 NOR4_X2 _32339_ (.A1(_09843_),
    .A2(_09849_),
    .A3(_09853_),
    .A4(_09856_),
    .ZN(_09857_));
 AND4_X2 _32340_ (.A1(_09815_),
    .A2(_09827_),
    .A3(_09839_),
    .A4(_09857_),
    .ZN(_09858_));
 AND2_X2 _32341_ (.A1(_09808_),
    .A2(_09858_),
    .ZN(_09859_));
 NOR2_X2 _32342_ (.A1(_06707_),
    .A2(_09859_),
    .ZN(_09860_));
 XOR2_X1 _32343_ (.A(_07644_),
    .B(_08999_),
    .Z(_09861_));
 XNOR2_X1 _32344_ (.A(_08806_),
    .B(_09861_),
    .ZN(_09862_));
 MUX2_X1 _32345_ (.A(_07643_),
    .B(_09862_),
    .S(_07242_),
    .Z(_09863_));
 AOI22_X1 _32346_ (.A1(\block_reg[0][26] ),
    .A2(_07806_),
    .B1(_08599_),
    .B2(_09863_),
    .ZN(_09864_));
 INV_X1 _32347_ (.A(_09864_),
    .ZN(_09865_));
 OAI22_X1 _32348_ (.A1(\block_reg[0][26] ),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_09863_),
    .ZN(_09866_));
 MUX2_X1 _32349_ (.A(_09865_),
    .B(_09866_),
    .S(_04678_),
    .Z(_09867_));
 NOR3_X1 _32350_ (.A1(_08177_),
    .A2(_09860_),
    .A3(_09867_),
    .ZN(_09868_));
 AOI21_X1 _32351_ (.A(_09868_),
    .B1(_06705_),
    .B2(_09247_),
    .ZN(_00720_));
 NOR3_X2 _32352_ (.A1(_09413_),
    .A2(_09306_),
    .A3(_09407_),
    .ZN(_09869_));
 NAND2_X1 _32353_ (.A1(_09612_),
    .A2(_09869_),
    .ZN(_09870_));
 NOR3_X2 _32354_ (.A1(_09306_),
    .A2(_09407_),
    .A3(_09343_),
    .ZN(_09871_));
 NOR2_X1 _32355_ (.A1(_09476_),
    .A2(_09671_),
    .ZN(_09872_));
 AOI22_X1 _32356_ (.A1(_09660_),
    .A2(_09871_),
    .B1(_09872_),
    .B2(_09293_),
    .ZN(_09873_));
 OAI21_X2 _32357_ (.A(_09870_),
    .B1(_09873_),
    .B2(_09754_),
    .ZN(_09874_));
 AOI21_X1 _32358_ (.A(_09595_),
    .B1(_09293_),
    .B2(_09335_),
    .ZN(_09875_));
 OAI21_X2 _32359_ (.A(_09625_),
    .B1(_09875_),
    .B2(_09754_),
    .ZN(_09876_));
 AOI22_X4 _32360_ (.A1(_09790_),
    .A2(_09874_),
    .B1(_09876_),
    .B2(_09251_),
    .ZN(_09877_));
 OR2_X1 _32361_ (.A1(_09498_),
    .A2(_09398_),
    .ZN(_09878_));
 NOR4_X1 _32362_ (.A1(_09374_),
    .A2(_09599_),
    .A3(_09542_),
    .A4(_09362_),
    .ZN(_09879_));
 NOR2_X1 _32363_ (.A1(_09878_),
    .A2(_09879_),
    .ZN(_09880_));
 NOR4_X2 _32364_ (.A1(_09272_),
    .A2(_09433_),
    .A3(_09333_),
    .A4(_09426_),
    .ZN(_09881_));
 AOI221_X2 _32365_ (.A(_09881_),
    .B1(_09441_),
    .B2(_09719_),
    .C1(_09374_),
    .C2(_09555_),
    .ZN(_09882_));
 NAND2_X1 _32366_ (.A1(_09539_),
    .A2(_09882_),
    .ZN(_09883_));
 NAND3_X1 _32367_ (.A1(_09651_),
    .A2(_09446_),
    .A3(_09362_),
    .ZN(_09884_));
 NOR3_X1 _32368_ (.A1(_09490_),
    .A2(_09334_),
    .A3(_09526_),
    .ZN(_09885_));
 OAI21_X1 _32369_ (.A(_09885_),
    .B1(_09481_),
    .B2(_09601_),
    .ZN(_09886_));
 NAND3_X1 _32370_ (.A1(_09560_),
    .A2(_09353_),
    .A3(_09372_),
    .ZN(_09887_));
 NAND3_X1 _32371_ (.A1(_09594_),
    .A2(_09650_),
    .A3(_09251_),
    .ZN(_09888_));
 NAND4_X2 _32372_ (.A1(_09884_),
    .A2(_09886_),
    .A3(_09887_),
    .A4(_09888_),
    .ZN(_09889_));
 NOR4_X4 _32373_ (.A1(_09820_),
    .A2(_09880_),
    .A3(_09883_),
    .A4(_09889_),
    .ZN(_09890_));
 AOI22_X2 _32374_ (.A1(_09485_),
    .A2(_09293_),
    .B1(_09769_),
    .B2(_09488_),
    .ZN(_09891_));
 NOR2_X1 _32375_ (.A1(_09492_),
    .A2(_09337_),
    .ZN(_09892_));
 NOR2_X1 _32376_ (.A1(_09476_),
    .A2(_09504_),
    .ZN(_09893_));
 AOI22_X2 _32377_ (.A1(_09550_),
    .A2(_09892_),
    .B1(_09893_),
    .B2(_09374_),
    .ZN(_09894_));
 OAI22_X2 _32378_ (.A1(_09709_),
    .A2(_09891_),
    .B1(_09894_),
    .B2(_09833_),
    .ZN(_09895_));
 NOR3_X1 _32379_ (.A1(_09579_),
    .A2(_09443_),
    .A3(_09408_),
    .ZN(_09896_));
 OAI21_X1 _32380_ (.A(_09535_),
    .B1(_09573_),
    .B2(_09572_),
    .ZN(_09897_));
 AOI22_X1 _32381_ (.A1(_09580_),
    .A2(_09871_),
    .B1(_09896_),
    .B2(_09897_),
    .ZN(_09898_));
 NOR2_X1 _32382_ (.A1(_09380_),
    .A2(_09898_),
    .ZN(_09899_));
 NOR2_X1 _32383_ (.A1(_09476_),
    .A2(_09592_),
    .ZN(_09900_));
 OAI21_X1 _32384_ (.A(_09900_),
    .B1(_09641_),
    .B2(_09374_),
    .ZN(_09901_));
 AOI21_X1 _32385_ (.A(_09657_),
    .B1(_09892_),
    .B2(_09376_),
    .ZN(_09902_));
 AOI21_X2 _32386_ (.A(_09580_),
    .B1(_09901_),
    .B2(_09902_),
    .ZN(_09903_));
 NOR3_X2 _32387_ (.A1(_09895_),
    .A2(_09899_),
    .A3(_09903_),
    .ZN(_09904_));
 AND2_X1 _32388_ (.A1(_09609_),
    .A2(_09614_),
    .ZN(_09905_));
 AOI221_X1 _32389_ (.A(_09589_),
    .B1(_09666_),
    .B2(_09854_),
    .C1(_09379_),
    .C2(_09378_),
    .ZN(_09906_));
 NAND3_X1 _32390_ (.A1(_09506_),
    .A2(_09723_),
    .A3(_09449_),
    .ZN(_09907_));
 OR3_X1 _32391_ (.A1(_09390_),
    .A2(_09448_),
    .A3(_09573_),
    .ZN(_09908_));
 NAND3_X1 _32392_ (.A1(_09415_),
    .A2(_09460_),
    .A3(_09448_),
    .ZN(_09909_));
 AOI21_X1 _32393_ (.A(_09907_),
    .B1(_09908_),
    .B2(_09909_),
    .ZN(_09910_));
 OR2_X1 _32394_ (.A1(_09406_),
    .A2(_09433_),
    .ZN(_09911_));
 NOR3_X1 _32395_ (.A1(_09415_),
    .A2(_09911_),
    .A3(_09370_),
    .ZN(_09912_));
 NAND2_X1 _32396_ (.A1(_09415_),
    .A2(_09501_),
    .ZN(_09913_));
 OAI21_X1 _32397_ (.A(_09572_),
    .B1(_09913_),
    .B2(_09822_),
    .ZN(_09914_));
 NAND3_X1 _32398_ (.A1(_09472_),
    .A2(_09353_),
    .A3(_09564_),
    .ZN(_09915_));
 NAND3_X1 _32399_ (.A1(_09336_),
    .A2(_09665_),
    .A3(_09347_),
    .ZN(_09916_));
 AOI21_X1 _32400_ (.A(_09345_),
    .B1(_09915_),
    .B2(_09916_),
    .ZN(_09917_));
 OAI33_X1 _32401_ (.A1(_09383_),
    .A2(_09906_),
    .A3(_09910_),
    .B1(_09912_),
    .B2(_09914_),
    .B3(_09917_),
    .ZN(_09918_));
 AOI22_X2 _32402_ (.A1(_09378_),
    .A2(_09379_),
    .B1(_09258_),
    .B2(_09459_),
    .ZN(_09919_));
 AOI22_X1 _32403_ (.A1(_09348_),
    .A2(_09623_),
    .B1(_09340_),
    .B2(_09341_),
    .ZN(_09920_));
 NOR4_X2 _32404_ (.A1(_09266_),
    .A2(_09721_),
    .A3(_09320_),
    .A4(_09328_),
    .ZN(_09921_));
 OAI211_X2 _32405_ (.A(_09524_),
    .B(_09919_),
    .C1(_09920_),
    .C2(_09921_),
    .ZN(_09922_));
 NAND3_X1 _32406_ (.A1(_09524_),
    .A2(_09665_),
    .A3(_09582_),
    .ZN(_09923_));
 AOI21_X1 _32407_ (.A(_09427_),
    .B1(_09922_),
    .B2(_09923_),
    .ZN(_09924_));
 OAI33_X1 _32408_ (.A1(_09594_),
    .A2(_09354_),
    .A3(_09589_),
    .B1(_09526_),
    .B2(_09911_),
    .B3(_09415_),
    .ZN(_09925_));
 AOI21_X2 _32409_ (.A(_09924_),
    .B1(_09925_),
    .B2(_09335_),
    .ZN(_09926_));
 AOI22_X2 _32410_ (.A1(_09401_),
    .A2(_09400_),
    .B1(_09381_),
    .B2(_09484_),
    .ZN(_09927_));
 OAI211_X2 _32411_ (.A(_09473_),
    .B(_09543_),
    .C1(_09836_),
    .C2(_09487_),
    .ZN(_09928_));
 NOR3_X1 _32412_ (.A1(_09364_),
    .A2(_09469_),
    .A3(_09291_),
    .ZN(_09929_));
 NOR4_X1 _32413_ (.A1(_09490_),
    .A2(_09361_),
    .A3(_09305_),
    .A4(_09422_),
    .ZN(_09930_));
 OAI21_X1 _32414_ (.A(_09492_),
    .B1(_09929_),
    .B2(_09930_),
    .ZN(_09931_));
 AND3_X1 _32415_ (.A1(_09927_),
    .A2(_09928_),
    .A3(_09931_),
    .ZN(_09932_));
 AND4_X1 _32416_ (.A1(_09905_),
    .A2(_09918_),
    .A3(_09926_),
    .A4(_09932_),
    .ZN(_09933_));
 NAND4_X4 _32417_ (.A1(_09877_),
    .A2(_09890_),
    .A3(_09904_),
    .A4(_09933_),
    .ZN(_09934_));
 OAI33_X1 _32418_ (.A1(_09364_),
    .A2(_09589_),
    .A3(_09408_),
    .B1(_09345_),
    .B2(_09424_),
    .B3(_09464_),
    .ZN(_09935_));
 AOI22_X2 _32419_ (.A1(_09626_),
    .A2(_09400_),
    .B1(_09935_),
    .B2(_09582_),
    .ZN(_09936_));
 OAI21_X1 _32420_ (.A(_09612_),
    .B1(_09485_),
    .B2(_09560_),
    .ZN(_09937_));
 NOR2_X1 _32421_ (.A1(_09610_),
    .A2(_09364_),
    .ZN(_09938_));
 AOI21_X1 _32422_ (.A(_09772_),
    .B1(_09937_),
    .B2(_09938_),
    .ZN(_09939_));
 AOI22_X2 _32423_ (.A1(_09594_),
    .A2(_09550_),
    .B1(_09422_),
    .B2(_09543_),
    .ZN(_09940_));
 OAI221_X2 _32424_ (.A(_09936_),
    .B1(_09939_),
    .B2(_09709_),
    .C1(_09345_),
    .C2(_09940_),
    .ZN(_09941_));
 AND2_X1 _32425_ (.A1(_09651_),
    .A2(_09591_),
    .ZN(_09942_));
 NAND3_X1 _32426_ (.A1(_09506_),
    .A2(_09722_),
    .A3(_09330_),
    .ZN(_09943_));
 OR3_X1 _32427_ (.A1(_09490_),
    .A2(_09439_),
    .A3(_09444_),
    .ZN(_09944_));
 NAND3_X1 _32428_ (.A1(_09490_),
    .A2(_09460_),
    .A3(_09347_),
    .ZN(_09945_));
 AOI21_X1 _32429_ (.A(_09943_),
    .B1(_09944_),
    .B2(_09945_),
    .ZN(_09946_));
 OR3_X1 _32430_ (.A1(_09748_),
    .A2(_09942_),
    .A3(_09946_),
    .ZN(_09947_));
 OR3_X4 _32431_ (.A1(_09718_),
    .A2(_09941_),
    .A3(_09947_),
    .ZN(_09948_));
 NOR2_X4 _32432_ (.A1(_09934_),
    .A2(_09948_),
    .ZN(_09949_));
 NOR2_X4 _32433_ (.A1(_06707_),
    .A2(_09949_),
    .ZN(_09950_));
 XNOR2_X1 _32434_ (.A(_07643_),
    .B(_07794_),
    .ZN(_09951_));
 XNOR2_X1 _32435_ (.A(_08892_),
    .B(_09951_),
    .ZN(_09952_));
 XNOR2_X1 _32436_ (.A(_07283_),
    .B(_08166_),
    .ZN(_09953_));
 XNOR2_X1 _32437_ (.A(_09952_),
    .B(_09953_),
    .ZN(_09954_));
 MUX2_X1 _32438_ (.A(_07795_),
    .B(_09954_),
    .S(_07242_),
    .Z(_09955_));
 AOI22_X1 _32439_ (.A1(\block_reg[0][27] ),
    .A2(_07806_),
    .B1(_08599_),
    .B2(_09955_),
    .ZN(_09956_));
 INV_X1 _32440_ (.A(_09956_),
    .ZN(_09957_));
 OAI22_X1 _32441_ (.A1(\block_reg[0][27] ),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_09955_),
    .ZN(_09958_));
 MUX2_X1 _32442_ (.A(_09957_),
    .B(_09958_),
    .S(_04803_),
    .Z(_09959_));
 NOR3_X1 _32443_ (.A1(_08906_),
    .A2(_09950_),
    .A3(_09959_),
    .ZN(_09960_));
 INV_X1 _32444_ (.A(_07795_),
    .ZN(_09961_));
 AOI21_X1 _32445_ (.A(_09960_),
    .B1(_06705_),
    .B2(_09961_),
    .ZN(_00721_));
 NAND2_X1 _32446_ (.A1(_09769_),
    .A2(_09828_),
    .ZN(_09962_));
 NAND2_X1 _32447_ (.A1(_09754_),
    .A2(_09599_),
    .ZN(_09963_));
 OAI21_X1 _32448_ (.A(_09962_),
    .B1(_09963_),
    .B2(_09630_),
    .ZN(_09964_));
 AOI22_X2 _32449_ (.A1(_09524_),
    .A2(_09624_),
    .B1(_09353_),
    .B2(_09347_),
    .ZN(_09965_));
 AOI21_X1 _32450_ (.A(_09334_),
    .B1(_09353_),
    .B2(_09564_),
    .ZN(_09966_));
 AOI21_X1 _32451_ (.A(_09337_),
    .B1(_09965_),
    .B2(_09966_),
    .ZN(_09967_));
 NAND2_X1 _32452_ (.A1(_09417_),
    .A2(_09965_),
    .ZN(_09968_));
 OAI221_X1 _32453_ (.A(_09580_),
    .B1(_09550_),
    .B2(_09967_),
    .C1(_09968_),
    .C2(_09603_),
    .ZN(_09969_));
 NAND3_X1 _32454_ (.A1(_09671_),
    .A2(_09353_),
    .A3(_09564_),
    .ZN(_09970_));
 OAI21_X1 _32455_ (.A(_09970_),
    .B1(_09965_),
    .B2(_09335_),
    .ZN(_09971_));
 AOI21_X1 _32456_ (.A(_09293_),
    .B1(_09971_),
    .B2(_09338_),
    .ZN(_09972_));
 OAI21_X1 _32457_ (.A(_09969_),
    .B1(_09972_),
    .B2(_09630_),
    .ZN(_09973_));
 MUX2_X2 _32458_ (.A(_09964_),
    .B(_09973_),
    .S(_09570_),
    .Z(_09974_));
 NOR2_X1 _32459_ (.A1(_09504_),
    .A2(_09709_),
    .ZN(_09975_));
 OAI33_X1 _32460_ (.A1(_09443_),
    .A2(_09573_),
    .A3(_09305_),
    .B1(_09343_),
    .B2(_09423_),
    .B3(_09291_),
    .ZN(_09976_));
 AOI222_X2 _32461_ (.A1(_09542_),
    .A2(_09452_),
    .B1(_09975_),
    .B2(_09976_),
    .C1(_09381_),
    .C2(_09603_),
    .ZN(_09977_));
 AOI21_X1 _32462_ (.A(_09626_),
    .B1(_09559_),
    .B2(_09579_),
    .ZN(_09978_));
 AOI22_X2 _32463_ (.A1(_09599_),
    .A2(_09552_),
    .B1(_09869_),
    .B2(_09621_),
    .ZN(_09979_));
 OAI221_X2 _32464_ (.A(_09977_),
    .B1(_09978_),
    .B2(_09418_),
    .C1(_09979_),
    .C2(_09422_),
    .ZN(_09980_));
 OAI22_X1 _32465_ (.A1(_09592_),
    .A2(_09709_),
    .B1(_09427_),
    .B2(_09671_),
    .ZN(_09981_));
 OAI33_X1 _32466_ (.A1(_09364_),
    .A2(_09596_),
    .A3(_09651_),
    .B1(_09408_),
    .B2(_09573_),
    .B3(_09574_),
    .ZN(_09982_));
 AOI22_X1 _32467_ (.A1(_09650_),
    .A2(_09981_),
    .B1(_09982_),
    .B2(_09541_),
    .ZN(_09983_));
 NOR3_X1 _32468_ (.A1(_09583_),
    .A2(_09295_),
    .A3(_09427_),
    .ZN(_09984_));
 NOR4_X1 _32469_ (.A1(_09492_),
    .A2(_09491_),
    .A3(_09295_),
    .A4(_09306_),
    .ZN(_09985_));
 OAI21_X1 _32470_ (.A(_09754_),
    .B1(_09984_),
    .B2(_09985_),
    .ZN(_09986_));
 NAND2_X1 _32471_ (.A1(_09983_),
    .A2(_09986_),
    .ZN(_09987_));
 NOR3_X2 _32472_ (.A1(_09800_),
    .A2(_09980_),
    .A3(_09987_),
    .ZN(_09988_));
 NAND3_X2 _32473_ (.A1(_09927_),
    .A2(_09928_),
    .A3(_09931_),
    .ZN(_09989_));
 NOR4_X2 _32474_ (.A1(_09506_),
    .A2(_09464_),
    .A3(_09424_),
    .A4(_09651_),
    .ZN(_09990_));
 AOI21_X2 _32475_ (.A(_09990_),
    .B1(_09900_),
    .B2(_09543_),
    .ZN(_09991_));
 NOR3_X1 _32476_ (.A1(_09413_),
    .A2(_09504_),
    .A3(_09596_),
    .ZN(_09992_));
 OAI21_X1 _32477_ (.A(_09380_),
    .B1(_09370_),
    .B2(_09448_),
    .ZN(_09993_));
 AOI21_X2 _32478_ (.A(_09992_),
    .B1(_09993_),
    .B2(_09560_),
    .ZN(_09994_));
 NAND2_X1 _32479_ (.A1(_09621_),
    .A2(_09624_),
    .ZN(_09995_));
 OAI22_X4 _32480_ (.A1(_09621_),
    .A2(_09991_),
    .B1(_09994_),
    .B2(_09995_),
    .ZN(_09996_));
 NAND2_X1 _32481_ (.A1(_09374_),
    .A2(_09502_),
    .ZN(_09997_));
 AOI22_X2 _32482_ (.A1(_09293_),
    .A2(_09499_),
    .B1(_09555_),
    .B2(_09362_),
    .ZN(_09998_));
 NAND2_X2 _32483_ (.A1(_09997_),
    .A2(_09998_),
    .ZN(_09999_));
 NOR4_X4 _32484_ (.A1(_09752_),
    .A2(_09989_),
    .A3(_09996_),
    .A4(_09999_),
    .ZN(_10000_));
 OAI221_X2 _32485_ (.A(_09468_),
    .B1(_09489_),
    .B2(_09790_),
    .C1(_09475_),
    .C2(_09660_),
    .ZN(_10001_));
 NAND2_X1 _32486_ (.A1(_09790_),
    .A2(_09651_),
    .ZN(_10002_));
 NOR3_X1 _32487_ (.A1(_09664_),
    .A2(_09583_),
    .A3(_09673_),
    .ZN(_10003_));
 AOI21_X1 _32488_ (.A(_10003_),
    .B1(_09601_),
    .B2(_09664_),
    .ZN(_10004_));
 AOI22_X2 _32489_ (.A1(_09650_),
    .A2(_09501_),
    .B1(_09362_),
    .B2(_09594_),
    .ZN(_10005_));
 OAI22_X2 _32490_ (.A1(_10002_),
    .A2(_10004_),
    .B1(_10005_),
    .B2(_09741_),
    .ZN(_10006_));
 NOR2_X2 _32491_ (.A1(_10001_),
    .A2(_10006_),
    .ZN(_10007_));
 NAND4_X4 _32492_ (.A1(_09670_),
    .A2(_09988_),
    .A3(_10000_),
    .A4(_10007_),
    .ZN(_10008_));
 NOR2_X4 _32493_ (.A1(_09974_),
    .A2(_10008_),
    .ZN(_10009_));
 NOR2_X4 _32494_ (.A1(_06707_),
    .A2(_10009_),
    .ZN(_10010_));
 XNOR2_X1 _32495_ (.A(_08166_),
    .B(_09127_),
    .ZN(_10011_));
 XNOR2_X1 _32496_ (.A(_07897_),
    .B(_07796_),
    .ZN(_10012_));
 XNOR2_X1 _32497_ (.A(_10011_),
    .B(_10012_),
    .ZN(_10013_));
 NAND2_X1 _32498_ (.A1(_08039_),
    .A2(_10013_),
    .ZN(_10014_));
 OAI21_X1 _32499_ (.A(_10014_),
    .B1(_08048_),
    .B2(_00330_),
    .ZN(_10015_));
 OAI22_X1 _32500_ (.A1(\block_reg[0][28] ),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_10015_),
    .ZN(_10016_));
 NOR2_X1 _32501_ (.A1(_04913_),
    .A2(_10016_),
    .ZN(_10017_));
 AOI22_X1 _32502_ (.A1(\block_reg[0][28] ),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_10015_),
    .ZN(_10018_));
 AOI21_X1 _32503_ (.A(_10017_),
    .B1(_10018_),
    .B2(_04913_),
    .ZN(_10019_));
 NOR3_X1 _32504_ (.A1(_08906_),
    .A2(_10010_),
    .A3(_10019_),
    .ZN(_10020_));
 INV_X1 _32505_ (.A(\core.enc_block.block_w0_reg[28] ),
    .ZN(_10021_));
 AOI21_X1 _32506_ (.A(_10020_),
    .B1(_06705_),
    .B2(_10021_),
    .ZN(_00722_));
 INV_X1 _32507_ (.A(_08041_),
    .ZN(_10022_));
 NOR3_X1 _32508_ (.A1(_09790_),
    .A2(_09673_),
    .A3(_09307_),
    .ZN(_10023_));
 OAI21_X1 _32509_ (.A(_09570_),
    .B1(_09829_),
    .B2(_10023_),
    .ZN(_10024_));
 NOR2_X1 _32510_ (.A1(_09535_),
    .A2(_09536_),
    .ZN(_10025_));
 XNOR2_X1 _32511_ (.A(_09439_),
    .B(_09335_),
    .ZN(_10026_));
 NAND3_X1 _32512_ (.A1(_10025_),
    .A2(_09552_),
    .A3(_10026_),
    .ZN(_10027_));
 AOI21_X1 _32513_ (.A(_09754_),
    .B1(_10024_),
    .B2(_10027_),
    .ZN(_10028_));
 NOR2_X1 _32514_ (.A1(_09580_),
    .A2(_09384_),
    .ZN(_10029_));
 NOR4_X2 _32515_ (.A1(_09476_),
    .A2(_09504_),
    .A3(_09515_),
    .A4(_09424_),
    .ZN(_10030_));
 OAI21_X1 _32516_ (.A(_09485_),
    .B1(_09330_),
    .B2(_09476_),
    .ZN(_10031_));
 NOR3_X2 _32517_ (.A1(_09386_),
    .A2(_09360_),
    .A3(_09290_),
    .ZN(_10032_));
 AOI22_X1 _32518_ (.A1(_10029_),
    .A2(_10030_),
    .B1(_10031_),
    .B2(_10032_),
    .ZN(_10033_));
 NOR3_X2 _32519_ (.A1(_09584_),
    .A2(_09596_),
    .A3(_09334_),
    .ZN(_10034_));
 AOI22_X2 _32520_ (.A1(_09702_),
    .A2(_10034_),
    .B1(_09850_),
    .B2(_09601_),
    .ZN(_10035_));
 NAND2_X1 _32521_ (.A1(_10025_),
    .A2(_09538_),
    .ZN(_10036_));
 NAND2_X1 _32522_ (.A1(_09570_),
    .A2(_09335_),
    .ZN(_10037_));
 OAI221_X1 _32523_ (.A(_10033_),
    .B1(_10035_),
    .B2(_09630_),
    .C1(_10036_),
    .C2(_10037_),
    .ZN(_10038_));
 NOR4_X1 _32524_ (.A1(_09594_),
    .A2(_09583_),
    .A3(_09295_),
    .A4(_09427_),
    .ZN(_10039_));
 NOR4_X1 _32525_ (.A1(_09594_),
    .A2(_09596_),
    .A3(_09585_),
    .A4(_09589_),
    .ZN(_10040_));
 OAI21_X1 _32526_ (.A(_09335_),
    .B1(_10039_),
    .B2(_10040_),
    .ZN(_10041_));
 NOR3_X1 _32527_ (.A1(_09660_),
    .A2(_09673_),
    .A3(_09586_),
    .ZN(_10042_));
 OAI21_X1 _32528_ (.A(_09521_),
    .B1(_09809_),
    .B2(_10042_),
    .ZN(_10043_));
 AOI222_X2 _32529_ (.A1(_09376_),
    .A2(_09502_),
    .B1(_09613_),
    .B2(_09626_),
    .C1(_09381_),
    .C2(_09374_),
    .ZN(_10044_));
 NOR4_X1 _32530_ (.A1(_09583_),
    .A2(_09295_),
    .A3(_09709_),
    .A4(_09612_),
    .ZN(_10045_));
 NOR4_X1 _32531_ (.A1(_09584_),
    .A2(_09586_),
    .A3(_09592_),
    .A4(_09709_),
    .ZN(_10046_));
 NOR4_X1 _32532_ (.A1(_09307_),
    .A2(_09585_),
    .A3(_09370_),
    .A4(_09371_),
    .ZN(_10047_));
 NOR4_X1 _32533_ (.A1(_09491_),
    .A2(_09585_),
    .A3(_09370_),
    .A4(_09408_),
    .ZN(_10048_));
 NOR4_X1 _32534_ (.A1(_10045_),
    .A2(_10046_),
    .A3(_10047_),
    .A4(_10048_),
    .ZN(_10049_));
 NAND4_X1 _32535_ (.A1(_10041_),
    .A2(_10043_),
    .A3(_10044_),
    .A4(_10049_),
    .ZN(_10050_));
 NAND2_X1 _32536_ (.A1(_09524_),
    .A2(_09624_),
    .ZN(_10051_));
 OR2_X1 _32537_ (.A1(_09498_),
    .A2(_09427_),
    .ZN(_10052_));
 MUX2_X1 _32538_ (.A(_09402_),
    .B(_09345_),
    .S(_09610_),
    .Z(_10053_));
 NAND3_X1 _32539_ (.A1(_09560_),
    .A2(_09665_),
    .A3(_09330_),
    .ZN(_10054_));
 OAI222_X2 _32540_ (.A1(_10051_),
    .A2(_09878_),
    .B1(_10052_),
    .B2(_09625_),
    .C1(_10053_),
    .C2(_10054_),
    .ZN(_10055_));
 OR4_X1 _32541_ (.A1(_09924_),
    .A2(_09942_),
    .A3(_09946_),
    .A4(_10055_),
    .ZN(_10056_));
 NOR4_X1 _32542_ (.A1(_10028_),
    .A2(_10038_),
    .A3(_10050_),
    .A4(_10056_),
    .ZN(_10057_));
 AND2_X1 _32543_ (.A1(_09983_),
    .A2(_09986_),
    .ZN(_10058_));
 AOI22_X1 _32544_ (.A1(_09347_),
    .A2(_09671_),
    .B1(_09564_),
    .B2(_09582_),
    .ZN(_10059_));
 NOR3_X1 _32545_ (.A1(_09660_),
    .A2(_09584_),
    .A3(_10059_),
    .ZN(_10060_));
 NAND4_X1 _32546_ (.A1(_09524_),
    .A2(_09353_),
    .A3(_09592_),
    .A4(_09422_),
    .ZN(_10061_));
 OAI211_X2 _32547_ (.A(_09524_),
    .B(_09635_),
    .C1(_09417_),
    .C2(_09582_),
    .ZN(_10062_));
 AOI21_X1 _32548_ (.A(_09664_),
    .B1(_10061_),
    .B2(_10062_),
    .ZN(_10063_));
 OAI21_X1 _32549_ (.A(_09630_),
    .B1(_10060_),
    .B2(_10063_),
    .ZN(_10064_));
 NOR2_X1 _32550_ (.A1(_09384_),
    .A2(_09668_),
    .ZN(_10065_));
 NAND2_X1 _32551_ (.A1(_09338_),
    .A2(_09911_),
    .ZN(_10066_));
 OAI221_X1 _32552_ (.A(_09446_),
    .B1(_09772_),
    .B2(_09338_),
    .C1(_10065_),
    .C2(_10066_),
    .ZN(_10067_));
 AND4_X1 _32553_ (.A1(_09815_),
    .A2(_10058_),
    .A3(_10064_),
    .A4(_10067_),
    .ZN(_10068_));
 NAND2_X1 _32554_ (.A1(_09430_),
    .A2(_09442_),
    .ZN(_10069_));
 AOI22_X2 _32555_ (.A1(_09637_),
    .A2(_09251_),
    .B1(_09500_),
    .B2(_09487_),
    .ZN(_10070_));
 AOI21_X1 _32556_ (.A(_10030_),
    .B1(_09650_),
    .B2(_09664_),
    .ZN(_10071_));
 OAI22_X2 _32557_ (.A1(_09338_),
    .A2(_10070_),
    .B1(_10071_),
    .B2(_09833_),
    .ZN(_10072_));
 NOR4_X2 _32558_ (.A1(_10069_),
    .A2(_09727_),
    .A3(_09748_),
    .A4(_10072_),
    .ZN(_10073_));
 NAND3_X2 _32559_ (.A1(_10057_),
    .A2(_10068_),
    .A3(_10073_),
    .ZN(_10074_));
 OR2_X4 _32560_ (.A1(_09569_),
    .A2(_10074_),
    .ZN(_10075_));
 NAND2_X2 _32561_ (.A1(_07260_),
    .A2(_10075_),
    .ZN(_10076_));
 XNOR2_X1 _32562_ (.A(_08043_),
    .B(_07896_),
    .ZN(_10077_));
 OR2_X1 _32563_ (.A1(_09173_),
    .A2(_10077_),
    .ZN(_10078_));
 NAND2_X1 _32564_ (.A1(_09173_),
    .A2(_10077_),
    .ZN(_10079_));
 NAND3_X1 _32565_ (.A1(_08722_),
    .A2(_10078_),
    .A3(_10079_),
    .ZN(_10080_));
 OAI21_X2 _32566_ (.A(_10080_),
    .B1(_08048_),
    .B2(_00333_),
    .ZN(_10081_));
 NAND2_X1 _32567_ (.A1(_07808_),
    .A2(_10081_),
    .ZN(_10082_));
 INV_X1 _32568_ (.A(\block_reg[0][29] ),
    .ZN(_10083_));
 OAI21_X1 _32569_ (.A(_10082_),
    .B1(_07248_),
    .B2(_10083_),
    .ZN(_10084_));
 OAI22_X1 _32570_ (.A1(\block_reg[0][29] ),
    .A2(_07251_),
    .B1(_07254_),
    .B2(_10081_),
    .ZN(_10085_));
 MUX2_X1 _32571_ (.A(_10084_),
    .B(_10085_),
    .S(_04288_),
    .Z(_10086_));
 NOR2_X1 _32572_ (.A1(_07224_),
    .A2(_10086_),
    .ZN(_10087_));
 AOI22_X1 _32573_ (.A1(_10022_),
    .A2(_08177_),
    .B1(_10076_),
    .B2(_10087_),
    .ZN(_00723_));
 BUF_X2 _32574_ (.A(\core.enc_block.block_w0_reg[2] ),
    .Z(_10088_));
 INV_X1 _32575_ (.A(_10088_),
    .ZN(_10089_));
 NOR4_X2 _32576_ (.A1(_06922_),
    .A2(_06853_),
    .A3(_08911_),
    .A4(_07087_),
    .ZN(_10090_));
 NOR2_X2 _32577_ (.A1(_06974_),
    .A2(_07102_),
    .ZN(_10091_));
 AOI221_X2 _32578_ (.A(_10090_),
    .B1(_07030_),
    .B2(_07083_),
    .C1(_07146_),
    .C2(_10091_),
    .ZN(_10092_));
 NAND2_X1 _32579_ (.A1(_07020_),
    .A2(_08934_),
    .ZN(_10093_));
 OAI221_X2 _32580_ (.A(_10092_),
    .B1(_07209_),
    .B2(_10093_),
    .C1(_07203_),
    .C2(_07204_),
    .ZN(_10094_));
 NAND4_X1 _32581_ (.A1(_07067_),
    .A2(_07046_),
    .A3(_07159_),
    .A4(_08968_),
    .ZN(_10095_));
 NOR2_X1 _32582_ (.A1(_06922_),
    .A2(_07051_),
    .ZN(_10096_));
 AOI22_X2 _32583_ (.A1(_06947_),
    .A2(_06906_),
    .B1(_10096_),
    .B2(_07146_),
    .ZN(_10097_));
 AOI222_X2 _32584_ (.A1(_06991_),
    .A2(_07048_),
    .B1(_07082_),
    .B2(_06985_),
    .C1(_07151_),
    .C2(_06989_),
    .ZN(_10098_));
 NAND3_X2 _32585_ (.A1(_10095_),
    .A2(_10097_),
    .A3(_10098_),
    .ZN(_10099_));
 NOR2_X2 _32586_ (.A1(_06955_),
    .A2(_06962_),
    .ZN(_10100_));
 NOR2_X1 _32587_ (.A1(_07011_),
    .A2(_07050_),
    .ZN(_10101_));
 OAI21_X1 _32588_ (.A(_10100_),
    .B1(_10101_),
    .B2(_06906_),
    .ZN(_10102_));
 NOR3_X1 _32589_ (.A1(_07099_),
    .A2(_07053_),
    .A3(_07202_),
    .ZN(_10103_));
 NOR3_X1 _32590_ (.A1(_07067_),
    .A2(_07131_),
    .A3(_07099_),
    .ZN(_10104_));
 OAI21_X1 _32591_ (.A(_06964_),
    .B1(_10103_),
    .B2(_10104_),
    .ZN(_10105_));
 NOR3_X1 _32592_ (.A1(_07068_),
    .A2(_07092_),
    .A3(_07078_),
    .ZN(_10106_));
 NOR3_X1 _32593_ (.A1(_07058_),
    .A2(_07080_),
    .A3(_07107_),
    .ZN(_10107_));
 OAI21_X1 _32594_ (.A(_06957_),
    .B1(_10106_),
    .B2(_10107_),
    .ZN(_10108_));
 OAI22_X1 _32595_ (.A1(_07028_),
    .A2(_07046_),
    .B1(_07102_),
    .B2(_07093_),
    .ZN(_10109_));
 AOI22_X1 _32596_ (.A1(_07146_),
    .A2(_08942_),
    .B1(_10109_),
    .B2(_07083_),
    .ZN(_10110_));
 NAND4_X1 _32597_ (.A1(_10102_),
    .A2(_10105_),
    .A3(_10108_),
    .A4(_10110_),
    .ZN(_10111_));
 NOR4_X1 _32598_ (.A1(_07085_),
    .A2(_07086_),
    .A3(_07099_),
    .A4(_07080_),
    .ZN(_10112_));
 NOR4_X1 _32599_ (.A1(_07112_),
    .A2(_07068_),
    .A3(_07078_),
    .A4(_07080_),
    .ZN(_10113_));
 OAI21_X1 _32600_ (.A(_07165_),
    .B1(_10112_),
    .B2(_10113_),
    .ZN(_10114_));
 NAND3_X1 _32601_ (.A1(_08941_),
    .A2(_08944_),
    .A3(_10114_),
    .ZN(_10115_));
 OR4_X2 _32602_ (.A1(_10094_),
    .A2(_10099_),
    .A3(_10111_),
    .A4(_10115_),
    .ZN(_10116_));
 NOR4_X2 _32603_ (.A1(_07091_),
    .A2(_06885_),
    .A3(_06943_),
    .A4(_06944_),
    .ZN(_10117_));
 NOR4_X1 _32604_ (.A1(_06921_),
    .A2(_06902_),
    .A3(_06914_),
    .A4(_06968_),
    .ZN(_10118_));
 OR2_X1 _32605_ (.A1(_10117_),
    .A2(_10118_),
    .ZN(_10119_));
 NAND2_X1 _32606_ (.A1(_06731_),
    .A2(_06874_),
    .ZN(_10120_));
 OR2_X2 _32607_ (.A1(_06904_),
    .A2(_06885_),
    .ZN(_10121_));
 AOI21_X2 _32608_ (.A(_10120_),
    .B1(_10121_),
    .B2(_06900_),
    .ZN(_10122_));
 OR3_X1 _32609_ (.A1(_06899_),
    .A2(_06910_),
    .A3(_08927_),
    .ZN(_10123_));
 NAND4_X1 _32610_ (.A1(_07104_),
    .A2(_07128_),
    .A3(_07129_),
    .A4(_07119_),
    .ZN(_10124_));
 OAI21_X1 _32611_ (.A(_10124_),
    .B1(_10121_),
    .B2(_07120_),
    .ZN(_10125_));
 AOI221_X2 _32612_ (.A(_10119_),
    .B1(_10122_),
    .B2(_10123_),
    .C1(_07155_),
    .C2(_10125_),
    .ZN(_10126_));
 NOR2_X1 _32613_ (.A1(_07208_),
    .A2(_07051_),
    .ZN(_10127_));
 NAND3_X1 _32614_ (.A1(_07129_),
    .A2(_07122_),
    .A3(_07059_),
    .ZN(_10128_));
 AOI21_X1 _32615_ (.A(_07062_),
    .B1(_08925_),
    .B2(_10128_),
    .ZN(_10129_));
 OAI21_X2 _32616_ (.A(_07155_),
    .B1(_10127_),
    .B2(_10129_),
    .ZN(_10130_));
 AOI21_X2 _32617_ (.A(_07112_),
    .B1(_08939_),
    .B2(_07017_),
    .ZN(_10131_));
 AOI22_X4 _32618_ (.A1(_08926_),
    .A2(_07083_),
    .B1(_10131_),
    .B2(_06999_),
    .ZN(_10132_));
 OAI211_X4 _32619_ (.A(_10126_),
    .B(_10130_),
    .C1(_10132_),
    .C2(_07144_),
    .ZN(_10133_));
 NAND2_X1 _32620_ (.A1(_07130_),
    .A2(_07184_),
    .ZN(_10134_));
 AOI221_X2 _32621_ (.A(_06870_),
    .B1(_06845_),
    .B2(_06787_),
    .C1(_06858_),
    .C2(_07109_),
    .ZN(_10135_));
 OAI33_X1 _32622_ (.A1(_07058_),
    .A2(_07165_),
    .A3(_10134_),
    .B1(_10135_),
    .B2(_07204_),
    .B3(_07106_),
    .ZN(_10136_));
 NAND2_X1 _32623_ (.A1(_07085_),
    .A2(_10136_),
    .ZN(_10137_));
 AOI22_X2 _32624_ (.A1(_07062_),
    .A2(_07204_),
    .B1(_10121_),
    .B2(_07200_),
    .ZN(_10138_));
 OAI221_X2 _32625_ (.A(_07060_),
    .B1(_07045_),
    .B2(_10138_),
    .C1(_06995_),
    .C2(_07058_),
    .ZN(_10139_));
 OAI21_X2 _32626_ (.A(_10137_),
    .B1(_10139_),
    .B2(_07085_),
    .ZN(_10140_));
 NOR4_X1 _32627_ (.A1(_07076_),
    .A2(_07137_),
    .A3(_07092_),
    .A4(_07107_),
    .ZN(_10141_));
 OAI21_X1 _32628_ (.A(_07058_),
    .B1(_07141_),
    .B2(_10141_),
    .ZN(_10142_));
 NAND2_X1 _32629_ (.A1(_07055_),
    .A2(_07147_),
    .ZN(_10143_));
 NOR3_X1 _32630_ (.A1(_07137_),
    .A2(_07011_),
    .A3(_07028_),
    .ZN(_10144_));
 OAI221_X2 _32631_ (.A(_07129_),
    .B1(_06947_),
    .B2(_10144_),
    .C1(_06836_),
    .C2(_06834_),
    .ZN(_10145_));
 AOI22_X2 _32632_ (.A1(_07045_),
    .A2(_07152_),
    .B1(_08942_),
    .B2(_06906_),
    .ZN(_10146_));
 NAND4_X2 _32633_ (.A1(_10142_),
    .A2(_10143_),
    .A3(_10145_),
    .A4(_10146_),
    .ZN(_10147_));
 NOR3_X1 _32634_ (.A1(_06971_),
    .A2(_07025_),
    .A3(_07093_),
    .ZN(_10148_));
 NAND4_X1 _32635_ (.A1(_06814_),
    .A2(_06767_),
    .A3(_06744_),
    .A4(_06881_),
    .ZN(_10149_));
 OAI21_X1 _32636_ (.A(_06891_),
    .B1(_07120_),
    .B2(_10149_),
    .ZN(_10150_));
 NOR2_X1 _32637_ (.A1(_07105_),
    .A2(_07011_),
    .ZN(_10151_));
 AOI21_X1 _32638_ (.A(_10148_),
    .B1(_10150_),
    .B2(_10151_),
    .ZN(_10152_));
 AND2_X1 _32639_ (.A1(_06932_),
    .A2(_10124_),
    .ZN(_10153_));
 NOR2_X1 _32640_ (.A1(_07005_),
    .A2(_08943_),
    .ZN(_10154_));
 OAI33_X1 _32641_ (.A1(_07028_),
    .A2(_10152_),
    .A3(_10153_),
    .B1(_10154_),
    .B2(_07074_),
    .B3(_07102_),
    .ZN(_10155_));
 OR3_X2 _32642_ (.A1(_06901_),
    .A2(_10147_),
    .A3(_10155_),
    .ZN(_10156_));
 OR4_X4 _32643_ (.A1(_10116_),
    .A2(_10133_),
    .A3(_10140_),
    .A4(_10156_),
    .ZN(_10157_));
 NOR2_X1 _32644_ (.A1(_06922_),
    .A2(_10134_),
    .ZN(_10158_));
 NAND3_X2 _32645_ (.A1(_07120_),
    .A2(_07130_),
    .A3(_07184_),
    .ZN(_10159_));
 NOR2_X1 _32646_ (.A1(_07058_),
    .A2(_10159_),
    .ZN(_10160_));
 NOR2_X1 _32647_ (.A1(_07069_),
    .A2(_07187_),
    .ZN(_10161_));
 OAI21_X1 _32648_ (.A(_07067_),
    .B1(_10160_),
    .B2(_10161_),
    .ZN(_10162_));
 AOI221_X2 _32649_ (.A(_07058_),
    .B1(_07005_),
    .B2(_07202_),
    .C1(_07201_),
    .C2(_07178_),
    .ZN(_10163_));
 OAI22_X2 _32650_ (.A1(_07187_),
    .A2(_07144_),
    .B1(_10159_),
    .B2(_07067_),
    .ZN(_10164_));
 AOI221_X2 _32651_ (.A(_10164_),
    .B1(_06906_),
    .B2(_07144_),
    .C1(_06787_),
    .C2(_06845_),
    .ZN(_10165_));
 OAI21_X2 _32652_ (.A(_10162_),
    .B1(_10163_),
    .B2(_10165_),
    .ZN(_10166_));
 MUX2_X2 _32653_ (.A(_10158_),
    .B(_10166_),
    .S(_07106_),
    .Z(_10167_));
 OAI21_X4 _32654_ (.A(_07662_),
    .B1(_10157_),
    .B2(_10167_),
    .ZN(_10168_));
 XNOR2_X1 _32655_ (.A(_07274_),
    .B(_08999_),
    .ZN(_10169_));
 XNOR2_X1 _32656_ (.A(_07647_),
    .B(_10169_),
    .ZN(_10170_));
 NAND2_X1 _32657_ (.A1(_07801_),
    .A2(_10170_),
    .ZN(_10171_));
 BUF_X4 _32658_ (.A(_08722_),
    .Z(_10172_));
 OAI21_X2 _32659_ (.A(_10171_),
    .B1(_10172_),
    .B2(_00367_),
    .ZN(_10173_));
 OAI221_X2 _32660_ (.A(_04698_),
    .B1(_09223_),
    .B2(_10173_),
    .C1(_09221_),
    .C2(\block_reg[0][2] ),
    .ZN(_10174_));
 AOI22_X1 _32661_ (.A1(\block_reg[0][2] ),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_10173_),
    .ZN(_10175_));
 OAI21_X1 _32662_ (.A(_10175_),
    .B1(_04697_),
    .B2(_04685_),
    .ZN(_10176_));
 AOI21_X2 _32663_ (.A(_06704_),
    .B1(_10174_),
    .B2(_10176_),
    .ZN(_10177_));
 AOI22_X1 _32664_ (.A1(_10089_),
    .A2(_08177_),
    .B1(_10168_),
    .B2(_10177_),
    .ZN(_00724_));
 INV_X1 _32665_ (.A(_09705_),
    .ZN(_10178_));
 OAI21_X4 _32666_ (.A(_10178_),
    .B1(_09496_),
    .B2(_09568_),
    .ZN(_10179_));
 MUX2_X1 _32667_ (.A(_09250_),
    .B(_09446_),
    .S(_09610_),
    .Z(_10180_));
 NOR3_X1 _32668_ (.A1(_09439_),
    .A2(_09364_),
    .A3(_09612_),
    .ZN(_10181_));
 AOI222_X2 _32669_ (.A1(_09626_),
    .A2(_09499_),
    .B1(_09502_),
    .B2(_09401_),
    .C1(_10180_),
    .C2(_10181_),
    .ZN(_10182_));
 NOR3_X1 _32670_ (.A1(_09307_),
    .A2(_09383_),
    .A3(_09585_),
    .ZN(_10183_));
 OAI21_X1 _32671_ (.A(_09802_),
    .B1(_10183_),
    .B2(_09550_),
    .ZN(_10184_));
 NOR4_X1 _32672_ (.A1(_09394_),
    .A2(_09396_),
    .A3(_09296_),
    .A4(_09298_),
    .ZN(_10185_));
 AOI22_X2 _32673_ (.A1(_09239_),
    .A2(_09249_),
    .B1(_09274_),
    .B2(_09281_),
    .ZN(_10186_));
 MUX2_X2 _32674_ (.A(_10185_),
    .B(_10186_),
    .S(_09610_),
    .Z(_10187_));
 NOR3_X2 _32675_ (.A1(_09664_),
    .A2(_09584_),
    .A3(_09422_),
    .ZN(_10188_));
 OAI21_X2 _32676_ (.A(_09535_),
    .B1(_09573_),
    .B2(_09671_),
    .ZN(_10189_));
 NOR4_X4 _32677_ (.A1(_09337_),
    .A2(_09443_),
    .A3(_09306_),
    .A4(_09709_),
    .ZN(_10190_));
 AOI22_X4 _32678_ (.A1(_10187_),
    .A2(_10188_),
    .B1(_10189_),
    .B2(_10190_),
    .ZN(_10191_));
 AOI222_X2 _32679_ (.A1(_09405_),
    .A2(_09499_),
    .B1(_09641_),
    .B2(_09403_),
    .C1(_09613_),
    .C2(_09376_),
    .ZN(_10192_));
 NAND4_X2 _32680_ (.A1(_10182_),
    .A2(_10184_),
    .A3(_10191_),
    .A4(_10192_),
    .ZN(_10193_));
 NOR3_X2 _32681_ (.A1(_09653_),
    .A2(_09941_),
    .A3(_10193_),
    .ZN(_10194_));
 NAND2_X1 _32682_ (.A1(_09251_),
    .A2(_09603_),
    .ZN(_10195_));
 NAND3_X1 _32683_ (.A1(_09621_),
    .A2(_09374_),
    .A3(_09627_),
    .ZN(_10196_));
 NAND4_X2 _32684_ (.A1(_09544_),
    .A2(_09547_),
    .A3(_10195_),
    .A4(_10196_),
    .ZN(_10197_));
 NOR4_X4 _32685_ (.A1(_09640_),
    .A2(_09805_),
    .A3(_09999_),
    .A4(_10197_),
    .ZN(_10198_));
 NAND2_X1 _32686_ (.A1(_09790_),
    .A2(_09626_),
    .ZN(_10199_));
 MUX2_X1 _32687_ (.A(_09354_),
    .B(_09625_),
    .S(_09660_),
    .Z(_10200_));
 OAI221_X2 _32688_ (.A(_09754_),
    .B1(_10199_),
    .B2(_09570_),
    .C1(_10200_),
    .C2(_09790_),
    .ZN(_10201_));
 NOR2_X1 _32689_ (.A1(_09293_),
    .A2(_09869_),
    .ZN(_10202_));
 OAI221_X2 _32690_ (.A(_09338_),
    .B1(_09427_),
    .B2(_09720_),
    .C1(_10202_),
    .C2(_09790_),
    .ZN(_10203_));
 NAND3_X2 _32691_ (.A1(_09384_),
    .A2(_10201_),
    .A3(_10203_),
    .ZN(_10204_));
 NOR4_X2 _32692_ (.A1(_09433_),
    .A2(_09392_),
    .A3(_09402_),
    .A4(_09422_),
    .ZN(_10205_));
 AOI221_X2 _32693_ (.A(_10205_),
    .B1(_10032_),
    .B2(_09329_),
    .C1(_09549_),
    .C2(_09401_),
    .ZN(_10206_));
 AOI21_X1 _32694_ (.A(_09488_),
    .B1(_09405_),
    .B2(_09504_),
    .ZN(_10207_));
 NAND2_X1 _32695_ (.A1(_09572_),
    .A2(_09446_),
    .ZN(_10208_));
 AOI22_X1 _32696_ (.A1(_09601_),
    .A2(_09410_),
    .B1(_09362_),
    .B2(_09471_),
    .ZN(_10209_));
 OAI221_X2 _32697_ (.A(_10206_),
    .B1(_10207_),
    .B2(_10208_),
    .C1(_10209_),
    .C2(_09664_),
    .ZN(_10210_));
 NOR3_X1 _32698_ (.A1(_09415_),
    .A2(_09535_),
    .A3(_09515_),
    .ZN(_10211_));
 NOR2_X1 _32699_ (.A1(_09610_),
    .A2(_09573_),
    .ZN(_10212_));
 AOI21_X1 _32700_ (.A(_10211_),
    .B1(_10186_),
    .B2(_10212_),
    .ZN(_10213_));
 NOR4_X1 _32701_ (.A1(_09412_),
    .A2(_09390_),
    .A3(_09439_),
    .A4(_09342_),
    .ZN(_10214_));
 AOI21_X1 _32702_ (.A(_10214_),
    .B1(_09439_),
    .B2(_09413_),
    .ZN(_10215_));
 OAI33_X1 _32703_ (.A1(_09443_),
    .A2(_09383_),
    .A3(_10213_),
    .B1(_10215_),
    .B2(_09536_),
    .B3(_09573_),
    .ZN(_10216_));
 OAI21_X1 _32704_ (.A(_09702_),
    .B1(_10034_),
    .B2(_09601_),
    .ZN(_10217_));
 OAI21_X1 _32705_ (.A(_10217_),
    .B1(_09831_),
    .B2(_09380_),
    .ZN(_10218_));
 AOI221_X2 _32706_ (.A(_10210_),
    .B1(_10216_),
    .B2(_09338_),
    .C1(_10218_),
    .C2(_09790_),
    .ZN(_10219_));
 NAND4_X4 _32707_ (.A1(_10194_),
    .A2(_10198_),
    .A3(_10204_),
    .A4(_10219_),
    .ZN(_10220_));
 NOR2_X4 _32708_ (.A1(_10179_),
    .A2(_10220_),
    .ZN(_10221_));
 NOR2_X4 _32709_ (.A1(_06707_),
    .A2(_10221_),
    .ZN(_10222_));
 CLKBUF_X3 _32710_ (.A(_07901_),
    .Z(_10223_));
 XOR2_X2 _32711_ (.A(_07329_),
    .B(_08041_),
    .Z(_10224_));
 XNOR2_X1 _32712_ (.A(_08106_),
    .B(_08110_),
    .ZN(_10225_));
 XNOR2_X2 _32713_ (.A(_10224_),
    .B(_10225_),
    .ZN(_10226_));
 XNOR2_X1 _32714_ (.A(_08227_),
    .B(_10226_),
    .ZN(_10227_));
 NOR2_X1 _32715_ (.A1(_10223_),
    .A2(_10227_),
    .ZN(_10228_));
 AOI21_X2 _32716_ (.A(_10228_),
    .B1(_07902_),
    .B2(_00336_),
    .ZN(_10229_));
 OAI22_X1 _32717_ (.A1(\block_reg[0][30] ),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_10229_),
    .ZN(_10230_));
 NAND2_X1 _32718_ (.A1(_07808_),
    .A2(_10229_),
    .ZN(_10231_));
 CLKBUF_X3 _32719_ (.A(_07247_),
    .Z(_10232_));
 OAI21_X1 _32720_ (.A(_10231_),
    .B1(_10232_),
    .B2(_05194_),
    .ZN(_10233_));
 MUX2_X1 _32721_ (.A(_10230_),
    .B(_10233_),
    .S(_04310_),
    .Z(_10234_));
 NOR3_X2 _32722_ (.A1(_08906_),
    .A2(_10222_),
    .A3(_10234_),
    .ZN(_10235_));
 INV_X1 _32723_ (.A(_08107_),
    .ZN(_10236_));
 AOI21_X1 _32724_ (.A(_10235_),
    .B1(_06705_),
    .B2(_10236_),
    .ZN(_00725_));
 NAND2_X1 _32725_ (.A1(_09374_),
    .A2(_09384_),
    .ZN(_10237_));
 OAI33_X1 _32726_ (.A1(_09560_),
    .A2(_09443_),
    .A3(_09444_),
    .B1(_09335_),
    .B2(_09295_),
    .B3(_09583_),
    .ZN(_10238_));
 OAI21_X2 _32727_ (.A(_09251_),
    .B1(_09976_),
    .B2(_10238_),
    .ZN(_10239_));
 OAI21_X2 _32728_ (.A(_09338_),
    .B1(_10237_),
    .B2(_10239_),
    .ZN(_10240_));
 NAND2_X1 _32729_ (.A1(_09446_),
    .A2(_09871_),
    .ZN(_10241_));
 OAI21_X1 _32730_ (.A(_09543_),
    .B1(_09346_),
    .B2(_09654_),
    .ZN(_10242_));
 NAND3_X2 _32731_ (.A1(_10239_),
    .A2(_10241_),
    .A3(_10242_),
    .ZN(_10243_));
 OAI33_X1 _32732_ (.A1(_09535_),
    .A2(_09574_),
    .A3(_09583_),
    .B1(_09295_),
    .B2(_09307_),
    .B3(_09621_),
    .ZN(_10244_));
 AOI22_X4 _32733_ (.A1(_09473_),
    .A2(_09405_),
    .B1(_10244_),
    .B2(_09754_),
    .ZN(_10245_));
 OAI22_X4 _32734_ (.A1(_09745_),
    .A2(_09605_),
    .B1(_10245_),
    .B2(_09570_),
    .ZN(_10246_));
 AOI22_X4 _32735_ (.A1(_10240_),
    .A2(_10243_),
    .B1(_10246_),
    .B2(_09384_),
    .ZN(_10247_));
 AOI21_X1 _32736_ (.A(_09990_),
    .B1(_09293_),
    .B2(_09702_),
    .ZN(_10248_));
 OAI22_X2 _32737_ (.A1(_09370_),
    .A2(_09746_),
    .B1(_10248_),
    .B2(_09630_),
    .ZN(_10249_));
 AOI21_X2 _32738_ (.A(_09980_),
    .B1(_10249_),
    .B2(_09833_),
    .ZN(_10250_));
 NAND2_X1 _32739_ (.A1(_09447_),
    .A2(_09462_),
    .ZN(_10251_));
 NOR4_X4 _32740_ (.A1(_10251_),
    .A2(_09758_),
    .A3(_09768_),
    .A4(_10210_),
    .ZN(_10252_));
 NAND3_X4 _32741_ (.A1(_10247_),
    .A2(_10250_),
    .A3(_10252_),
    .ZN(_10253_));
 NOR2_X1 _32742_ (.A1(_09832_),
    .A2(_09835_),
    .ZN(_10254_));
 AND2_X1 _32743_ (.A1(_10064_),
    .A2(_10067_),
    .ZN(_10255_));
 AOI21_X1 _32744_ (.A(_09651_),
    .B1(_09330_),
    .B2(_09570_),
    .ZN(_10256_));
 OAI33_X1 _32745_ (.A1(_09295_),
    .A2(_09485_),
    .A3(_09586_),
    .B1(_10256_),
    .B2(_09583_),
    .B3(_09673_),
    .ZN(_10257_));
 AOI21_X2 _32746_ (.A(_09606_),
    .B1(_10257_),
    .B2(_09630_),
    .ZN(_10258_));
 NAND4_X4 _32747_ (.A1(_10254_),
    .A2(_09926_),
    .A3(_10255_),
    .A4(_10258_),
    .ZN(_10259_));
 NOR2_X4 _32748_ (.A1(_10253_),
    .A2(_10259_),
    .ZN(_10260_));
 NOR2_X4 _32749_ (.A1(_06707_),
    .A2(_10260_),
    .ZN(_10261_));
 XNOR2_X1 _32750_ (.A(_07792_),
    .B(_08108_),
    .ZN(_10262_));
 XNOR2_X1 _32751_ (.A(_08165_),
    .B(_10262_),
    .ZN(_10263_));
 NAND2_X1 _32752_ (.A1(_08896_),
    .A2(_10263_),
    .ZN(_10264_));
 BUF_X4 _32753_ (.A(_08038_),
    .Z(_10265_));
 OAI21_X1 _32754_ (.A(_10264_),
    .B1(_10265_),
    .B2(_00339_),
    .ZN(_10266_));
 AOI22_X1 _32755_ (.A1(\block_reg[0][31] ),
    .A2(_07806_),
    .B1(_08599_),
    .B2(_10266_),
    .ZN(_10267_));
 INV_X1 _32756_ (.A(_10267_),
    .ZN(_10268_));
 CLKBUF_X3 _32757_ (.A(_07253_),
    .Z(_10269_));
 OAI22_X1 _32758_ (.A1(\block_reg[0][31] ),
    .A2(_08607_),
    .B1(_10269_),
    .B2(_10266_),
    .ZN(_10270_));
 MUX2_X1 _32759_ (.A(_10268_),
    .B(_10270_),
    .S(_04348_),
    .Z(_10271_));
 NOR3_X1 _32760_ (.A1(_08906_),
    .A2(_10261_),
    .A3(_10271_),
    .ZN(_10272_));
 INV_X1 _32761_ (.A(_07235_),
    .ZN(_10273_));
 AOI21_X1 _32762_ (.A(_10272_),
    .B1(_06705_),
    .B2(_10273_),
    .ZN(_00726_));
 CLKBUF_X2 _32763_ (.A(\core.enc_block.block_w0_reg[3] ),
    .Z(_10274_));
 INV_X1 _32764_ (.A(_10274_),
    .ZN(_10275_));
 NAND2_X1 _32765_ (.A1(_06853_),
    .A2(_07128_),
    .ZN(_10276_));
 NAND2_X1 _32766_ (.A1(_06731_),
    .A2(_07011_),
    .ZN(_10277_));
 MUX2_X1 _32767_ (.A(_08939_),
    .B(_07017_),
    .S(_06913_),
    .Z(_10278_));
 OAI33_X1 _32768_ (.A1(_07050_),
    .A2(_07102_),
    .A3(_10276_),
    .B1(_10277_),
    .B2(_10278_),
    .B3(_07097_),
    .ZN(_10279_));
 OAI33_X1 _32769_ (.A1(_08911_),
    .A2(_07087_),
    .A3(_07017_),
    .B1(_10121_),
    .B2(_07186_),
    .B3(_06899_),
    .ZN(_10280_));
 MUX2_X1 _32770_ (.A(_10279_),
    .B(_10280_),
    .S(_07059_),
    .Z(_10281_));
 NOR4_X2 _32771_ (.A1(_07077_),
    .A2(_07165_),
    .A3(_07052_),
    .A4(_07074_),
    .ZN(_10282_));
 AOI22_X4 _32772_ (.A1(_06947_),
    .A2(_07045_),
    .B1(_10282_),
    .B2(_07162_),
    .ZN(_10283_));
 XNOR2_X1 _32773_ (.A(_06900_),
    .B(_07120_),
    .ZN(_10284_));
 AOI21_X1 _32774_ (.A(_08908_),
    .B1(_10284_),
    .B2(_06957_),
    .ZN(_10285_));
 NAND2_X1 _32775_ (.A1(_07129_),
    .A2(_07184_),
    .ZN(_10286_));
 OAI21_X1 _32776_ (.A(_10283_),
    .B1(_10285_),
    .B2(_10286_),
    .ZN(_10287_));
 NOR4_X2 _32777_ (.A1(_07097_),
    .A2(_07028_),
    .A3(_06955_),
    .A4(_07052_),
    .ZN(_10288_));
 AOI21_X1 _32778_ (.A(_10288_),
    .B1(_07151_),
    .B2(_07083_),
    .ZN(_10289_));
 AOI22_X1 _32779_ (.A1(_06991_),
    .A2(_06947_),
    .B1(_07047_),
    .B2(_07005_),
    .ZN(_10290_));
 NOR4_X4 _32780_ (.A1(_07091_),
    .A2(_06856_),
    .A3(_06943_),
    .A4(_06968_),
    .ZN(_10291_));
 OAI22_X4 _32781_ (.A1(_07138_),
    .A2(_07083_),
    .B1(_07048_),
    .B2(_10291_),
    .ZN(_10292_));
 NAND3_X1 _32782_ (.A1(_10289_),
    .A2(_10290_),
    .A3(_10292_),
    .ZN(_10293_));
 OR4_X2 _32783_ (.A1(_06854_),
    .A2(_10281_),
    .A3(_10287_),
    .A4(_10293_),
    .ZN(_10294_));
 NAND3_X1 _32784_ (.A1(_07067_),
    .A2(_07137_),
    .A3(_07045_),
    .ZN(_10295_));
 NAND2_X1 _32785_ (.A1(_07093_),
    .A2(_07148_),
    .ZN(_10296_));
 AOI21_X1 _32786_ (.A(_07058_),
    .B1(_10295_),
    .B2(_10296_),
    .ZN(_10297_));
 OR2_X1 _32787_ (.A1(_07097_),
    .A2(_07140_),
    .ZN(_10298_));
 OAI33_X1 _32788_ (.A1(_07120_),
    .A2(_10298_),
    .A3(_07017_),
    .B1(_10134_),
    .B2(_07020_),
    .B3(_06900_),
    .ZN(_10299_));
 AND2_X1 _32789_ (.A1(_07112_),
    .A2(_10299_),
    .ZN(_10300_));
 NOR3_X1 _32790_ (.A1(_06922_),
    .A2(_06880_),
    .A3(_07087_),
    .ZN(_10301_));
 AOI21_X1 _32791_ (.A(_07119_),
    .B1(_06971_),
    .B2(_07061_),
    .ZN(_10302_));
 NOR3_X1 _32792_ (.A1(_07104_),
    .A2(_07011_),
    .A3(_06928_),
    .ZN(_10303_));
 OAI21_X1 _32793_ (.A(_10301_),
    .B1(_10302_),
    .B2(_10303_),
    .ZN(_10304_));
 MUX2_X1 _32794_ (.A(_06928_),
    .B(_07001_),
    .S(_07131_),
    .Z(_10305_));
 NAND4_X1 _32795_ (.A1(_07168_),
    .A2(_06971_),
    .A3(_07130_),
    .A4(_10305_),
    .ZN(_10306_));
 OAI21_X1 _32796_ (.A(_06829_),
    .B1(_07048_),
    .B2(_07152_),
    .ZN(_10307_));
 NAND4_X1 _32797_ (.A1(_10146_),
    .A2(_10304_),
    .A3(_10306_),
    .A4(_10307_),
    .ZN(_10308_));
 NOR2_X4 _32798_ (.A1(_06928_),
    .A2(_06962_),
    .ZN(_10309_));
 AOI22_X1 _32799_ (.A1(_06833_),
    .A2(_07117_),
    .B1(_10309_),
    .B2(_08943_),
    .ZN(_10310_));
 NOR2_X1 _32800_ (.A1(_07106_),
    .A2(_10310_),
    .ZN(_10311_));
 OR4_X2 _32801_ (.A1(_10297_),
    .A2(_10300_),
    .A3(_10308_),
    .A4(_10311_),
    .ZN(_10312_));
 OAI22_X4 _32802_ (.A1(_07035_),
    .A2(_07091_),
    .B1(_06932_),
    .B2(_06971_),
    .ZN(_10313_));
 NOR2_X2 _32803_ (.A1(_06891_),
    .A2(_07046_),
    .ZN(_10314_));
 OAI33_X1 _32804_ (.A1(_07035_),
    .A2(_07025_),
    .A3(_07091_),
    .B1(_06856_),
    .B2(_07140_),
    .B3(_06874_),
    .ZN(_10315_));
 AOI22_X4 _32805_ (.A1(_10313_),
    .A2(_10314_),
    .B1(_10315_),
    .B2(_07059_),
    .ZN(_10316_));
 OAI21_X1 _32806_ (.A(_07105_),
    .B1(_07077_),
    .B2(_07070_),
    .ZN(_10317_));
 AOI21_X2 _32807_ (.A(_07178_),
    .B1(_10317_),
    .B2(_07059_),
    .ZN(_10318_));
 OAI21_X2 _32808_ (.A(_06833_),
    .B1(_07023_),
    .B2(_07051_),
    .ZN(_10319_));
 OAI22_X4 _32809_ (.A1(_06922_),
    .A2(_10316_),
    .B1(_10318_),
    .B2(_10319_),
    .ZN(_10320_));
 AND2_X1 _32810_ (.A1(_07137_),
    .A2(_07177_),
    .ZN(_10321_));
 NAND2_X1 _32811_ (.A1(_07168_),
    .A2(_07055_),
    .ZN(_10322_));
 NAND2_X2 _32812_ (.A1(_07051_),
    .A2(_07093_),
    .ZN(_10323_));
 AOI22_X2 _32813_ (.A1(_08926_),
    .A2(_06973_),
    .B1(_06999_),
    .B2(_06964_),
    .ZN(_10324_));
 NOR4_X1 _32814_ (.A1(_06795_),
    .A2(_06902_),
    .A3(_06914_),
    .A4(_06872_),
    .ZN(_10325_));
 AOI21_X1 _32815_ (.A(_10325_),
    .B1(_06989_),
    .B2(_07057_),
    .ZN(_10326_));
 OAI222_X2 _32816_ (.A1(_10322_),
    .A2(_10323_),
    .B1(_10324_),
    .B2(_08938_),
    .C1(_10326_),
    .C2(_06877_),
    .ZN(_10327_));
 OR4_X2 _32817_ (.A1(_07173_),
    .A2(_10117_),
    .A3(_10321_),
    .A4(_10327_),
    .ZN(_10328_));
 NOR4_X4 _32818_ (.A1(_10294_),
    .A2(_10312_),
    .A3(_10320_),
    .A4(_10328_),
    .ZN(_10329_));
 OAI21_X2 _32819_ (.A(_10130_),
    .B1(_10132_),
    .B2(_07144_),
    .ZN(_10330_));
 NAND2_X1 _32820_ (.A1(_06928_),
    .A2(_06857_),
    .ZN(_10331_));
 AOI21_X1 _32821_ (.A(_07039_),
    .B1(_06906_),
    .B2(_06928_),
    .ZN(_10332_));
 MUX2_X1 _32822_ (.A(_10331_),
    .B(_10332_),
    .S(_07104_),
    .Z(_10333_));
 NOR2_X1 _32823_ (.A1(_07076_),
    .A2(_07159_),
    .ZN(_10334_));
 NAND2_X1 _32824_ (.A1(_07005_),
    .A2(_10323_),
    .ZN(_10335_));
 AOI221_X2 _32825_ (.A(_07069_),
    .B1(_10333_),
    .B2(_10334_),
    .C1(_10335_),
    .C2(_07085_),
    .ZN(_10336_));
 NOR4_X1 _32826_ (.A1(_07106_),
    .A2(_07092_),
    .A3(_07107_),
    .A4(_07201_),
    .ZN(_10337_));
 NOR3_X1 _32827_ (.A1(_07092_),
    .A2(_07099_),
    .A3(_06877_),
    .ZN(_10338_));
 OAI21_X1 _32828_ (.A(_07058_),
    .B1(_10337_),
    .B2(_10338_),
    .ZN(_10339_));
 NOR2_X1 _32829_ (.A1(_07137_),
    .A2(_07004_),
    .ZN(_10340_));
 NOR3_X1 _32830_ (.A1(_07099_),
    .A2(_07144_),
    .A3(_07080_),
    .ZN(_10341_));
 OAI21_X1 _32831_ (.A(_10340_),
    .B1(_10341_),
    .B2(_07159_),
    .ZN(_10342_));
 NOR4_X2 _32832_ (.A1(_07112_),
    .A2(_07137_),
    .A3(_07011_),
    .A4(_07098_),
    .ZN(_10343_));
 AND2_X1 _32833_ (.A1(_07131_),
    .A2(_10135_),
    .ZN(_10344_));
 OAI221_X2 _32834_ (.A(_06845_),
    .B1(_06860_),
    .B2(_06870_),
    .C1(_06887_),
    .C2(_06783_),
    .ZN(_10345_));
 NOR2_X1 _32835_ (.A1(_07131_),
    .A2(_10345_),
    .ZN(_10346_));
 OAI21_X2 _32836_ (.A(_10343_),
    .B1(_10344_),
    .B2(_10346_),
    .ZN(_10347_));
 NOR3_X1 _32837_ (.A1(_07137_),
    .A2(_07099_),
    .A3(_07080_),
    .ZN(_10348_));
 OAI21_X2 _32838_ (.A(_07162_),
    .B1(_07096_),
    .B2(_10348_),
    .ZN(_10349_));
 NAND4_X4 _32839_ (.A1(_10339_),
    .A2(_10342_),
    .A3(_10347_),
    .A4(_10349_),
    .ZN(_10350_));
 NOR4_X4 _32840_ (.A1(_08955_),
    .A2(_10330_),
    .A3(_10336_),
    .A4(_10350_),
    .ZN(_10351_));
 AND2_X2 _32841_ (.A1(_10329_),
    .A2(_10351_),
    .ZN(_10352_));
 OR2_X2 _32842_ (.A1(_06706_),
    .A2(_10352_),
    .ZN(_10353_));
 CLKBUF_X3 _32843_ (.A(_08038_),
    .Z(_10354_));
 XNOR2_X1 _32844_ (.A(_07791_),
    .B(_07795_),
    .ZN(_10355_));
 XNOR2_X1 _32845_ (.A(_07235_),
    .B(_10355_),
    .ZN(_10356_));
 XOR2_X1 _32846_ (.A(_00313_),
    .B(_07648_),
    .Z(_10357_));
 XNOR2_X1 _32847_ (.A(_09951_),
    .B(_10357_),
    .ZN(_10358_));
 XNOR2_X1 _32848_ (.A(_10356_),
    .B(_10358_),
    .ZN(_10359_));
 NAND2_X1 _32849_ (.A1(_10354_),
    .A2(_10359_),
    .ZN(_10360_));
 OAI21_X2 _32850_ (.A(_10360_),
    .B1(_09217_),
    .B2(_00370_),
    .ZN(_10361_));
 OAI221_X2 _32851_ (.A(_04832_),
    .B1(_09223_),
    .B2(_10361_),
    .C1(_09221_),
    .C2(\block_reg[0][3] ),
    .ZN(_10362_));
 NAND2_X1 _32852_ (.A1(_07908_),
    .A2(_10361_),
    .ZN(_10363_));
 INV_X1 _32853_ (.A(\block_reg[0][3] ),
    .ZN(_10364_));
 OAI21_X1 _32854_ (.A(_10363_),
    .B1(_07787_),
    .B2(_10364_),
    .ZN(_10365_));
 OR2_X1 _32855_ (.A1(_04832_),
    .A2(_10365_),
    .ZN(_10366_));
 AOI21_X2 _32856_ (.A(_06703_),
    .B1(_10362_),
    .B2(_10366_),
    .ZN(_10367_));
 AOI22_X1 _32857_ (.A1(_10275_),
    .A2(_08177_),
    .B1(_10353_),
    .B2(_10367_),
    .ZN(_00727_));
 BUF_X2 _32858_ (.A(\core.enc_block.block_w0_reg[4] ),
    .Z(_10368_));
 INV_X1 _32859_ (.A(_10368_),
    .ZN(_10369_));
 AOI21_X2 _32860_ (.A(_07153_),
    .B1(_08942_),
    .B2(_07055_),
    .ZN(_10370_));
 NOR4_X2 _32861_ (.A1(_06902_),
    .A2(_06856_),
    .A3(_06962_),
    .A4(_07001_),
    .ZN(_10371_));
 OAI22_X2 _32862_ (.A1(_06944_),
    .A2(_07004_),
    .B1(_07093_),
    .B2(_06943_),
    .ZN(_10372_));
 AOI221_X2 _32863_ (.A(_10371_),
    .B1(_07151_),
    .B2(_07023_),
    .C1(_06991_),
    .C2(_10372_),
    .ZN(_10373_));
 NAND4_X2 _32864_ (.A1(_07150_),
    .A2(_08936_),
    .A3(_10370_),
    .A4(_10373_),
    .ZN(_10374_));
 AOI22_X4 _32865_ (.A1(_07155_),
    .A2(_08927_),
    .B1(_10309_),
    .B2(_07146_),
    .ZN(_10375_));
 NOR3_X2 _32866_ (.A1(_06900_),
    .A2(_07090_),
    .A3(_07053_),
    .ZN(_10376_));
 AOI21_X2 _32867_ (.A(_10376_),
    .B1(_06964_),
    .B2(_08943_),
    .ZN(_10377_));
 OAI22_X4 _32868_ (.A1(_07062_),
    .A2(_10375_),
    .B1(_10377_),
    .B2(_07067_),
    .ZN(_10378_));
 NOR4_X4 _32869_ (.A1(_07003_),
    .A2(_07009_),
    .A3(_10374_),
    .A4(_10378_),
    .ZN(_10379_));
 OAI21_X1 _32870_ (.A(_08911_),
    .B1(_07053_),
    .B2(_07061_),
    .ZN(_10380_));
 NAND2_X1 _32871_ (.A1(_07126_),
    .A2(_10380_),
    .ZN(_10381_));
 AOI22_X2 _32872_ (.A1(_06744_),
    .A2(_07123_),
    .B1(_06923_),
    .B2(_06924_),
    .ZN(_10382_));
 MUX2_X1 _32873_ (.A(_08921_),
    .B(_10382_),
    .S(_06971_),
    .Z(_10383_));
 NOR3_X1 _32874_ (.A1(_07104_),
    .A2(_06880_),
    .A3(_07035_),
    .ZN(_10384_));
 AOI21_X1 _32875_ (.A(_08991_),
    .B1(_10383_),
    .B2(_10384_),
    .ZN(_10385_));
 AOI221_X2 _32876_ (.A(_07102_),
    .B1(_07204_),
    .B2(_07074_),
    .C1(_10381_),
    .C2(_10385_),
    .ZN(_10386_));
 OR2_X1 _32877_ (.A1(_08921_),
    .A2(_10382_),
    .ZN(_10387_));
 NOR4_X4 _32878_ (.A1(_06853_),
    .A2(_07035_),
    .A3(_07091_),
    .A4(_07028_),
    .ZN(_10388_));
 AOI22_X4 _32879_ (.A1(_06974_),
    .A2(_08962_),
    .B1(_10387_),
    .B2(_10388_),
    .ZN(_10389_));
 NAND3_X1 _32880_ (.A1(_07155_),
    .A2(_06906_),
    .A3(_10323_),
    .ZN(_10390_));
 NAND2_X1 _32881_ (.A1(_10389_),
    .A2(_10390_),
    .ZN(_10391_));
 AOI22_X1 _32882_ (.A1(_07178_),
    .A2(_07147_),
    .B1(_10340_),
    .B2(_07146_),
    .ZN(_10392_));
 AOI22_X2 _32883_ (.A1(_07005_),
    .A2(_06945_),
    .B1(_08908_),
    .B2(_07138_),
    .ZN(_10393_));
 NOR2_X1 _32884_ (.A1(_07086_),
    .A2(_07046_),
    .ZN(_10394_));
 NOR3_X1 _32885_ (.A1(_07076_),
    .A2(_07080_),
    .A3(_07107_),
    .ZN(_10395_));
 OAI21_X1 _32886_ (.A(_10394_),
    .B1(_10395_),
    .B2(_08956_),
    .ZN(_10396_));
 NAND3_X2 _32887_ (.A1(_10392_),
    .A2(_10393_),
    .A3(_10396_),
    .ZN(_10397_));
 NOR4_X4 _32888_ (.A1(_10099_),
    .A2(_10386_),
    .A3(_10391_),
    .A4(_10397_),
    .ZN(_10398_));
 AOI21_X1 _32889_ (.A(_07063_),
    .B1(_07050_),
    .B2(_07099_),
    .ZN(_10399_));
 AOI22_X1 _32890_ (.A1(_07062_),
    .A2(_07117_),
    .B1(_10399_),
    .B2(_07144_),
    .ZN(_10400_));
 OAI22_X2 _32891_ (.A1(_07017_),
    .A2(_10159_),
    .B1(_10400_),
    .B2(_07069_),
    .ZN(_10401_));
 AOI21_X2 _32892_ (.A(_07103_),
    .B1(_10401_),
    .B2(_07085_),
    .ZN(_10402_));
 AOI221_X2 _32893_ (.A(_10288_),
    .B1(_08923_),
    .B2(_07005_),
    .C1(_07138_),
    .C2(_07082_),
    .ZN(_10403_));
 AOI21_X1 _32894_ (.A(_07144_),
    .B1(_08943_),
    .B2(_07172_),
    .ZN(_10404_));
 NOR2_X1 _32895_ (.A1(_07066_),
    .A2(_06853_),
    .ZN(_10405_));
 AOI221_X2 _32896_ (.A(_07059_),
    .B1(_06847_),
    .B2(_06910_),
    .C1(_10405_),
    .C2(_06991_),
    .ZN(_10406_));
 OAI21_X2 _32897_ (.A(_10403_),
    .B1(_10404_),
    .B2(_10406_),
    .ZN(_10407_));
 NOR3_X1 _32898_ (.A1(_07068_),
    .A2(_07092_),
    .A3(_07107_),
    .ZN(_10408_));
 OAI21_X1 _32899_ (.A(_10405_),
    .B1(_10408_),
    .B2(_08943_),
    .ZN(_10409_));
 OAI221_X2 _32900_ (.A(_06809_),
    .B1(_07178_),
    .B2(_07083_),
    .C1(_06728_),
    .C2(_06712_),
    .ZN(_10410_));
 AOI21_X1 _32901_ (.A(_07144_),
    .B1(_10409_),
    .B2(_10410_),
    .ZN(_10411_));
 NOR3_X2 _32902_ (.A1(_10350_),
    .A2(_10407_),
    .A3(_10411_),
    .ZN(_10412_));
 NAND4_X4 _32903_ (.A1(_10379_),
    .A2(_10398_),
    .A3(_10402_),
    .A4(_10412_),
    .ZN(_10413_));
 NAND2_X2 _32904_ (.A1(_07662_),
    .A2(_10413_),
    .ZN(_10414_));
 XNOR2_X1 _32905_ (.A(_00314_),
    .B(_07790_),
    .ZN(_10415_));
 XNOR2_X1 _32906_ (.A(_07896_),
    .B(_10415_),
    .ZN(_10416_));
 XNOR2_X1 _32907_ (.A(_10356_),
    .B(_10416_),
    .ZN(_10417_));
 NAND2_X1 _32908_ (.A1(_08039_),
    .A2(_10417_),
    .ZN(_10418_));
 OAI21_X1 _32909_ (.A(_10418_),
    .B1(_08048_),
    .B2(_00350_),
    .ZN(_10419_));
 OAI22_X1 _32910_ (.A1(\block_reg[0][4] ),
    .A2(_07251_),
    .B1(_08608_),
    .B2(_10419_),
    .ZN(_10420_));
 NAND2_X1 _32911_ (.A1(_07229_),
    .A2(_10419_),
    .ZN(_10421_));
 OAI21_X1 _32912_ (.A(_10421_),
    .B1(_07248_),
    .B2(_06632_),
    .ZN(_10422_));
 MUX2_X1 _32913_ (.A(_10420_),
    .B(_10422_),
    .S(_04936_),
    .Z(_10423_));
 NOR2_X1 _32914_ (.A1(_07224_),
    .A2(_10423_),
    .ZN(_10424_));
 AOI22_X1 _32915_ (.A1(_10369_),
    .A2(_08177_),
    .B1(_10414_),
    .B2(_10424_),
    .ZN(_00728_));
 CLKBUF_X2 _32916_ (.A(\core.enc_block.block_w0_reg[5] ),
    .Z(_10425_));
 INV_X1 _32917_ (.A(_10425_),
    .ZN(_10426_));
 OAI33_X1 _32918_ (.A1(_07050_),
    .A2(_07120_),
    .A3(_07079_),
    .B1(_07070_),
    .B2(_07093_),
    .B3(_07077_),
    .ZN(_10427_));
 NOR2_X1 _32919_ (.A1(_07066_),
    .A2(_06974_),
    .ZN(_10428_));
 AOI22_X1 _32920_ (.A1(_07067_),
    .A2(_10427_),
    .B1(_10428_),
    .B2(_07055_),
    .ZN(_10429_));
 OR2_X1 _32921_ (.A1(_07069_),
    .A2(_10429_),
    .ZN(_10430_));
 AND2_X1 _32922_ (.A1(_10126_),
    .A2(_10430_),
    .ZN(_10431_));
 AOI22_X4 _32923_ (.A1(_07062_),
    .A2(_07146_),
    .B1(_07074_),
    .B2(_08952_),
    .ZN(_10432_));
 NOR3_X2 _32924_ (.A1(_07138_),
    .A2(_07046_),
    .A3(_06906_),
    .ZN(_10433_));
 OAI21_X2 _32925_ (.A(_07155_),
    .B1(_07083_),
    .B2(_07020_),
    .ZN(_10434_));
 OAI22_X4 _32926_ (.A1(_06922_),
    .A2(_10432_),
    .B1(_10433_),
    .B2(_10434_),
    .ZN(_10435_));
 NAND4_X2 _32927_ (.A1(_08930_),
    .A2(_08933_),
    .A3(_10389_),
    .A4(_10390_),
    .ZN(_10436_));
 NOR3_X1 _32928_ (.A1(_07092_),
    .A2(_07087_),
    .A3(_07051_),
    .ZN(_10437_));
 NOR3_X1 _32929_ (.A1(_07063_),
    .A2(_07087_),
    .A3(_07165_),
    .ZN(_10438_));
 OAI21_X2 _32930_ (.A(_06847_),
    .B1(_10437_),
    .B2(_10438_),
    .ZN(_10439_));
 NOR4_X4 _32931_ (.A1(_06894_),
    .A2(_06874_),
    .A3(_06876_),
    .A4(_07052_),
    .ZN(_10440_));
 NOR4_X2 _32932_ (.A1(_06731_),
    .A2(_07104_),
    .A3(_07077_),
    .A4(_07070_),
    .ZN(_10441_));
 OAI21_X2 _32933_ (.A(_07086_),
    .B1(_10440_),
    .B2(_10441_),
    .ZN(_10442_));
 NAND4_X4 _32934_ (.A1(_06948_),
    .A2(_10283_),
    .A3(_10439_),
    .A4(_10442_),
    .ZN(_10443_));
 NOR3_X1 _32935_ (.A1(_07131_),
    .A2(_06914_),
    .A3(_06951_),
    .ZN(_10444_));
 AOI221_X2 _32936_ (.A(_10444_),
    .B1(_07082_),
    .B2(_07146_),
    .C1(_08943_),
    .C2(_08923_),
    .ZN(_10445_));
 OAI21_X1 _32937_ (.A(_10345_),
    .B1(_10135_),
    .B2(_06731_),
    .ZN(_10446_));
 AOI22_X2 _32938_ (.A1(_08943_),
    .A2(_10309_),
    .B1(_10446_),
    .B2(_06857_),
    .ZN(_10447_));
 OAI211_X2 _32939_ (.A(_10098_),
    .B(_10445_),
    .C1(_10447_),
    .C2(_07062_),
    .ZN(_10448_));
 NOR4_X4 _32940_ (.A1(_10435_),
    .A2(_10436_),
    .A3(_10443_),
    .A4(_10448_),
    .ZN(_10449_));
 NOR4_X1 _32941_ (.A1(_06894_),
    .A2(_07057_),
    .A3(_07097_),
    .A4(_07140_),
    .ZN(_10450_));
 NOR4_X1 _32942_ (.A1(_08911_),
    .A2(_06928_),
    .A3(_07077_),
    .A4(_06962_),
    .ZN(_10451_));
 OAI21_X1 _32943_ (.A(_07061_),
    .B1(_10450_),
    .B2(_10451_),
    .ZN(_10452_));
 AOI22_X2 _32944_ (.A1(_07055_),
    .A2(_08942_),
    .B1(_10100_),
    .B2(_07159_),
    .ZN(_10453_));
 NOR4_X1 _32945_ (.A1(_07091_),
    .A2(_06885_),
    .A3(_07164_),
    .A4(_07001_),
    .ZN(_10454_));
 AOI211_X2 _32946_ (.A(_06855_),
    .B(_06914_),
    .C1(_06955_),
    .C2(_06968_),
    .ZN(_10455_));
 OAI21_X2 _32947_ (.A(_07168_),
    .B1(_10454_),
    .B2(_10455_),
    .ZN(_10456_));
 NAND4_X1 _32948_ (.A1(_10292_),
    .A2(_10452_),
    .A3(_10453_),
    .A4(_10456_),
    .ZN(_10457_));
 AOI22_X2 _32949_ (.A1(_06809_),
    .A2(_07159_),
    .B1(_07023_),
    .B2(_07200_),
    .ZN(_10458_));
 AND2_X1 _32950_ (.A1(_06894_),
    .A2(_08989_),
    .ZN(_10459_));
 AOI22_X2 _32951_ (.A1(_07076_),
    .A2(_08973_),
    .B1(_10459_),
    .B2(_06910_),
    .ZN(_10460_));
 AOI21_X1 _32952_ (.A(_06969_),
    .B1(_06996_),
    .B2(_07066_),
    .ZN(_10461_));
 OAI222_X2 _32953_ (.A1(_08938_),
    .A2(_10458_),
    .B1(_10460_),
    .B2(_07059_),
    .C1(_07086_),
    .C2(_10461_),
    .ZN(_10462_));
 AOI21_X2 _32954_ (.A(_07086_),
    .B1(_07006_),
    .B2(_07085_),
    .ZN(_10463_));
 NOR2_X1 _32955_ (.A1(_07105_),
    .A2(_06926_),
    .ZN(_10464_));
 AOI221_X2 _32956_ (.A(_07156_),
    .B1(_06819_),
    .B2(_06872_),
    .C1(_06799_),
    .C2(_06953_),
    .ZN(_10465_));
 OAI221_X2 _32957_ (.A(_07112_),
    .B1(_06974_),
    .B2(_10298_),
    .C1(_10464_),
    .C2(_10465_),
    .ZN(_10466_));
 AOI211_X2 _32958_ (.A(_10457_),
    .B(_10462_),
    .C1(_10463_),
    .C2(_10466_),
    .ZN(_10467_));
 NAND3_X2 _32959_ (.A1(_10431_),
    .A2(_10449_),
    .A3(_10467_),
    .ZN(_10468_));
 NOR3_X4 _32960_ (.A1(_07044_),
    .A2(_07073_),
    .A3(_10468_),
    .ZN(_10469_));
 OR2_X2 _32961_ (.A1(_06707_),
    .A2(_10469_),
    .ZN(_10470_));
 XNOR2_X1 _32962_ (.A(_08042_),
    .B(_09173_),
    .ZN(_10471_));
 XNOR2_X1 _32963_ (.A(_10021_),
    .B(_10471_),
    .ZN(_10472_));
 NAND2_X1 _32964_ (.A1(_08039_),
    .A2(_10472_),
    .ZN(_10473_));
 OAI21_X2 _32965_ (.A(_10473_),
    .B1(_08048_),
    .B2(_00353_),
    .ZN(_10474_));
 NAND2_X1 _32966_ (.A1(_07808_),
    .A2(_10474_),
    .ZN(_10475_));
 CLKBUF_X3 _32967_ (.A(_07247_),
    .Z(_10476_));
 INV_X1 _32968_ (.A(\block_reg[0][5] ),
    .ZN(_10477_));
 OAI21_X1 _32969_ (.A(_10475_),
    .B1(_10476_),
    .B2(_10477_),
    .ZN(_10478_));
 OAI22_X1 _32970_ (.A1(\block_reg[0][5] ),
    .A2(_07251_),
    .B1(_07254_),
    .B2(_10474_),
    .ZN(_10479_));
 MUX2_X1 _32971_ (.A(_10478_),
    .B(_10479_),
    .S(_04364_),
    .Z(_10480_));
 NOR2_X1 _32972_ (.A1(_07224_),
    .A2(_10480_),
    .ZN(_10481_));
 AOI22_X1 _32973_ (.A1(_10426_),
    .A2(_08177_),
    .B1(_10470_),
    .B2(_10481_),
    .ZN(_00729_));
 BUF_X2 _32974_ (.A(\core.enc_block.block_w0_reg[6] ),
    .Z(_10482_));
 INV_X1 _32975_ (.A(_10482_),
    .ZN(_10483_));
 NAND2_X1 _32976_ (.A1(_10466_),
    .A2(_10463_),
    .ZN(_10484_));
 OAI21_X1 _32977_ (.A(_07106_),
    .B1(_07178_),
    .B2(_07156_),
    .ZN(_10485_));
 AOI21_X2 _32978_ (.A(_07102_),
    .B1(_10485_),
    .B2(_08970_),
    .ZN(_10486_));
 NAND3_X1 _32979_ (.A1(_07168_),
    .A2(_06829_),
    .A3(_10323_),
    .ZN(_10487_));
 AOI21_X1 _32980_ (.A(_10118_),
    .B1(_07045_),
    .B2(_06947_),
    .ZN(_10488_));
 AOI22_X2 _32981_ (.A1(_07159_),
    .A2(_07030_),
    .B1(_07047_),
    .B2(_07083_),
    .ZN(_10489_));
 NAND4_X2 _32982_ (.A1(_06956_),
    .A2(_10487_),
    .A3(_10488_),
    .A4(_10489_),
    .ZN(_10490_));
 AOI22_X2 _32983_ (.A1(_07202_),
    .A2(_06999_),
    .B1(_07117_),
    .B2(_07112_),
    .ZN(_10491_));
 NAND4_X1 _32984_ (.A1(_06880_),
    .A2(_07130_),
    .A3(_07074_),
    .A4(_06896_),
    .ZN(_10492_));
 OAI22_X2 _32985_ (.A1(_07017_),
    .A2(_10491_),
    .B1(_10492_),
    .B2(_07069_),
    .ZN(_10493_));
 NOR3_X4 _32986_ (.A1(_10486_),
    .A2(_10490_),
    .A3(_10493_),
    .ZN(_10494_));
 NAND2_X1 _32987_ (.A1(_07086_),
    .A2(_07060_),
    .ZN(_10495_));
 AOI21_X2 _32988_ (.A(_10440_),
    .B1(_06957_),
    .B2(_06991_),
    .ZN(_10496_));
 OAI22_X4 _32989_ (.A1(_07180_),
    .A2(_07181_),
    .B1(_10495_),
    .B2(_10496_),
    .ZN(_10497_));
 NAND2_X1 _32990_ (.A1(_10370_),
    .A2(_10373_),
    .ZN(_10498_));
 OAI21_X1 _32991_ (.A(_06944_),
    .B1(_06974_),
    .B2(_07131_),
    .ZN(_10499_));
 NOR4_X2 _32992_ (.A1(_06971_),
    .A2(_06891_),
    .A3(_06932_),
    .A4(_06951_),
    .ZN(_10500_));
 AOI222_X2 _32993_ (.A1(_06947_),
    .A2(_07159_),
    .B1(_10499_),
    .B2(_10500_),
    .C1(_10100_),
    .C2(_06829_),
    .ZN(_10501_));
 NOR2_X1 _32994_ (.A1(_07061_),
    .A2(_08962_),
    .ZN(_10502_));
 AOI21_X2 _32995_ (.A(_07105_),
    .B1(_06833_),
    .B2(_07055_),
    .ZN(_10503_));
 OAI21_X2 _32996_ (.A(_10501_),
    .B1(_10502_),
    .B2(_10503_),
    .ZN(_10504_));
 NOR4_X4 _32997_ (.A1(_10497_),
    .A2(_10320_),
    .A3(_10498_),
    .A4(_10504_),
    .ZN(_10505_));
 AND2_X1 _32998_ (.A1(_07131_),
    .A2(_07200_),
    .ZN(_10506_));
 AND3_X1 _32999_ (.A1(_06852_),
    .A2(_06880_),
    .A3(_10345_),
    .ZN(_10507_));
 OAI21_X1 _33000_ (.A(_07011_),
    .B1(_10506_),
    .B2(_10507_),
    .ZN(_10508_));
 NAND2_X1 _33001_ (.A1(_08926_),
    .A2(_07184_),
    .ZN(_10509_));
 AOI221_X2 _33002_ (.A(_07077_),
    .B1(_10508_),
    .B2(_10509_),
    .C1(_06844_),
    .C2(_06842_),
    .ZN(_10510_));
 NOR3_X2 _33003_ (.A1(_07098_),
    .A2(_07119_),
    .A3(_07070_),
    .ZN(_10511_));
 NOR3_X1 _33004_ (.A1(_07087_),
    .A2(_07070_),
    .A3(_08938_),
    .ZN(_10512_));
 OAI21_X1 _33005_ (.A(_07086_),
    .B1(_10511_),
    .B2(_10512_),
    .ZN(_10513_));
 NAND4_X1 _33006_ (.A1(_06787_),
    .A2(_06845_),
    .A3(_06923_),
    .A4(_06924_),
    .ZN(_10514_));
 OAI33_X1 _33007_ (.A1(_06900_),
    .A2(_07079_),
    .A3(_06885_),
    .B1(_07070_),
    .B2(_10514_),
    .B3(_07097_),
    .ZN(_10515_));
 AOI21_X1 _33008_ (.A(_08956_),
    .B1(_10515_),
    .B2(_07066_),
    .ZN(_10516_));
 AOI21_X2 _33009_ (.A(_07106_),
    .B1(_10513_),
    .B2(_10516_),
    .ZN(_10517_));
 NOR2_X1 _33010_ (.A1(_07105_),
    .A2(_07028_),
    .ZN(_10518_));
 OAI22_X2 _33011_ (.A1(_07090_),
    .A2(_07091_),
    .B1(_07097_),
    .B2(_08911_),
    .ZN(_10519_));
 AOI22_X2 _33012_ (.A1(_07117_),
    .A2(_07172_),
    .B1(_10518_),
    .B2(_10519_),
    .ZN(_10520_));
 OAI33_X1 _33013_ (.A1(_06853_),
    .A2(_07090_),
    .A3(_07140_),
    .B1(_07052_),
    .B2(_06932_),
    .B3(_07025_),
    .ZN(_10521_));
 AOI22_X2 _33014_ (.A1(_06929_),
    .A2(_06957_),
    .B1(_07110_),
    .B2(_10521_),
    .ZN(_10522_));
 OAI21_X2 _33015_ (.A(_10520_),
    .B1(_10522_),
    .B2(_07086_),
    .ZN(_10523_));
 NOR4_X4 _33016_ (.A1(_10155_),
    .A2(_10510_),
    .A3(_10517_),
    .A4(_10523_),
    .ZN(_10524_));
 NAND4_X4 _33017_ (.A1(_10484_),
    .A2(_10494_),
    .A3(_10505_),
    .A4(_10524_),
    .ZN(_10525_));
 NOR3_X4 _33018_ (.A1(_07044_),
    .A2(_08916_),
    .A3(_10525_),
    .ZN(_10526_));
 OR2_X2 _33019_ (.A1(_06706_),
    .A2(_10526_),
    .ZN(_10527_));
 XOR2_X1 _33020_ (.A(_08109_),
    .B(_10224_),
    .Z(_10528_));
 NAND2_X1 _33021_ (.A1(_08039_),
    .A2(_10528_),
    .ZN(_10529_));
 OAI21_X2 _33022_ (.A(_10529_),
    .B1(_08048_),
    .B2(_00356_),
    .ZN(_10530_));
 NAND2_X1 _33023_ (.A1(_07808_),
    .A2(_10530_),
    .ZN(_10531_));
 INV_X1 _33024_ (.A(\block_reg[0][6] ),
    .ZN(_10532_));
 OAI21_X1 _33025_ (.A(_10531_),
    .B1(_10476_),
    .B2(_10532_),
    .ZN(_10533_));
 OAI22_X1 _33026_ (.A1(\block_reg[0][6] ),
    .A2(_07251_),
    .B1(_07254_),
    .B2(_10530_),
    .ZN(_10534_));
 MUX2_X1 _33027_ (.A(_10533_),
    .B(_10534_),
    .S(_04588_),
    .Z(_10535_));
 NOR2_X1 _33028_ (.A1(_07224_),
    .A2(_10535_),
    .ZN(_10536_));
 AOI22_X1 _33029_ (.A1(_10483_),
    .A2(_08177_),
    .B1(_10527_),
    .B2(_10536_),
    .ZN(_00730_));
 BUF_X4 _33030_ (.A(\core.enc_block.block_w0_reg[7] ),
    .Z(_10537_));
 INV_X1 _33031_ (.A(_10537_),
    .ZN(_10538_));
 AND2_X1 _33032_ (.A1(_08972_),
    .A2(_08985_),
    .ZN(_10539_));
 NAND4_X2 _33033_ (.A1(_07038_),
    .A2(_10292_),
    .A3(_10453_),
    .A4(_10456_),
    .ZN(_10540_));
 AOI22_X2 _33034_ (.A1(_07155_),
    .A2(_07178_),
    .B1(_10309_),
    .B2(_07138_),
    .ZN(_10541_));
 NAND3_X1 _33035_ (.A1(_07060_),
    .A2(_06847_),
    .A3(_07023_),
    .ZN(_10542_));
 AOI21_X2 _33036_ (.A(_07106_),
    .B1(_10541_),
    .B2(_10542_),
    .ZN(_10543_));
 NOR4_X4 _33037_ (.A1(_10147_),
    .A2(_10327_),
    .A3(_10540_),
    .A4(_10543_),
    .ZN(_10544_));
 OAI33_X1 _33038_ (.A1(_08943_),
    .A2(_07178_),
    .A3(_07045_),
    .B1(_10511_),
    .B2(_06849_),
    .B3(_06851_),
    .ZN(_10545_));
 OAI22_X2 _33039_ (.A1(_07208_),
    .A2(_07102_),
    .B1(_10545_),
    .B2(_07004_),
    .ZN(_10546_));
 AOI21_X2 _33040_ (.A(_10407_),
    .B1(_10546_),
    .B2(_06974_),
    .ZN(_10547_));
 OAI211_X2 _33041_ (.A(_07095_),
    .B(_10501_),
    .C1(_10502_),
    .C2(_10503_),
    .ZN(_10548_));
 NOR3_X1 _33042_ (.A1(_07061_),
    .A2(_07063_),
    .A3(_07050_),
    .ZN(_10549_));
 NOR4_X1 _33043_ (.A1(_07112_),
    .A2(_07105_),
    .A3(_08911_),
    .A4(_07078_),
    .ZN(_10550_));
 OAI21_X1 _33044_ (.A(_07183_),
    .B1(_10549_),
    .B2(_10550_),
    .ZN(_10551_));
 OAI221_X2 _33045_ (.A(_07137_),
    .B1(_07063_),
    .B2(_07050_),
    .C1(_07107_),
    .C2(_07053_),
    .ZN(_10552_));
 AOI21_X1 _33046_ (.A(_07063_),
    .B1(_07099_),
    .B2(_07078_),
    .ZN(_10553_));
 OAI211_X2 _33047_ (.A(_07162_),
    .B(_10552_),
    .C1(_10553_),
    .C2(_07106_),
    .ZN(_10554_));
 NAND4_X2 _33048_ (.A1(_07167_),
    .A2(_07169_),
    .A3(_10551_),
    .A4(_10554_),
    .ZN(_10555_));
 NAND2_X1 _33049_ (.A1(_07085_),
    .A2(_07060_),
    .ZN(_10556_));
 MUX2_X1 _33050_ (.A(_07208_),
    .B(_08970_),
    .S(_08968_),
    .Z(_10557_));
 AOI21_X1 _33051_ (.A(_10376_),
    .B1(_08943_),
    .B2(_07068_),
    .ZN(_10558_));
 OAI22_X2 _33052_ (.A1(_10556_),
    .A2(_10557_),
    .B1(_10558_),
    .B2(_10120_),
    .ZN(_10559_));
 AOI222_X2 _33053_ (.A1(_06847_),
    .A2(_07071_),
    .B1(_07147_),
    .B2(_06906_),
    .C1(_10091_),
    .C2(_07138_),
    .ZN(_10560_));
 AND3_X1 _33054_ (.A1(_07122_),
    .A2(_07126_),
    .A3(_07201_),
    .ZN(_10561_));
 AOI21_X1 _33055_ (.A(_10561_),
    .B1(_07138_),
    .B2(_07085_),
    .ZN(_10562_));
 OAI21_X2 _33056_ (.A(_10560_),
    .B1(_10562_),
    .B2(_08968_),
    .ZN(_10563_));
 NOR4_X4 _33057_ (.A1(_10548_),
    .A2(_10555_),
    .A3(_10559_),
    .A4(_10563_),
    .ZN(_10564_));
 NAND4_X4 _33058_ (.A1(_10539_),
    .A2(_10544_),
    .A3(_10547_),
    .A4(_10564_),
    .ZN(_10565_));
 NAND2_X2 _33059_ (.A1(_07662_),
    .A2(_10565_),
    .ZN(_10566_));
 XNOR2_X1 _33060_ (.A(_07338_),
    .B(_08107_),
    .ZN(_10567_));
 XNOR2_X1 _33061_ (.A(_08167_),
    .B(_10567_),
    .ZN(_10568_));
 NAND2_X1 _33062_ (.A1(_08039_),
    .A2(_10568_),
    .ZN(_10569_));
 OAI21_X2 _33063_ (.A(_10569_),
    .B1(_08048_),
    .B2(_06742_),
    .ZN(_10570_));
 NAND2_X1 _33064_ (.A1(_07808_),
    .A2(_10570_),
    .ZN(_10571_));
 INV_X1 _33065_ (.A(\block_reg[0][7] ),
    .ZN(_10572_));
 OAI21_X1 _33066_ (.A(_10571_),
    .B1(_10476_),
    .B2(_10572_),
    .ZN(_10573_));
 OAI22_X1 _33067_ (.A1(\block_reg[0][7] ),
    .A2(_07251_),
    .B1(_07254_),
    .B2(_10570_),
    .ZN(_10574_));
 MUX2_X1 _33068_ (.A(_10573_),
    .B(_10574_),
    .S(_04722_),
    .Z(_10575_));
 NOR2_X1 _33069_ (.A1(_07224_),
    .A2(_10575_),
    .ZN(_10576_));
 AOI22_X1 _33070_ (.A1(_10538_),
    .A2(_08177_),
    .B1(_10566_),
    .B2(_10576_),
    .ZN(_00731_));
 OAI21_X1 _33071_ (.A(_07417_),
    .B1(_07695_),
    .B2(_07437_),
    .ZN(_10577_));
 NAND2_X1 _33072_ (.A1(_07425_),
    .A2(_07769_),
    .ZN(_10578_));
 NOR3_X1 _33073_ (.A1(_07531_),
    .A2(_07984_),
    .A3(_07621_),
    .ZN(_10579_));
 AOI221_X2 _33074_ (.A(_07432_),
    .B1(_07407_),
    .B2(_07472_),
    .C1(_10578_),
    .C2(_10579_),
    .ZN(_10580_));
 NOR3_X1 _33075_ (.A1(_07408_),
    .A2(_07451_),
    .A3(_07694_),
    .ZN(_10581_));
 OAI21_X1 _33076_ (.A(_07457_),
    .B1(_07544_),
    .B2(_10581_),
    .ZN(_10582_));
 AOI21_X2 _33077_ (.A(_10577_),
    .B1(_10580_),
    .B2(_10582_),
    .ZN(_10583_));
 NAND2_X1 _33078_ (.A1(_07457_),
    .A2(_07404_),
    .ZN(_10584_));
 OAI21_X1 _33079_ (.A(_07408_),
    .B1(_07404_),
    .B2(_07884_),
    .ZN(_10585_));
 AOI21_X2 _33080_ (.A(_07388_),
    .B1(_10584_),
    .B2(_10585_),
    .ZN(_10586_));
 AOI22_X4 _33081_ (.A1(_07426_),
    .A2(_07513_),
    .B1(_07493_),
    .B2(_07818_),
    .ZN(_10587_));
 NOR3_X1 _33082_ (.A1(_07571_),
    .A2(_07451_),
    .A3(_07458_),
    .ZN(_10588_));
 OAI21_X1 _33083_ (.A(_07764_),
    .B1(_07987_),
    .B2(_10588_),
    .ZN(_10589_));
 AOI22_X1 _33084_ (.A1(_07362_),
    .A2(_07607_),
    .B1(_07703_),
    .B2(_07507_),
    .ZN(_10590_));
 NAND3_X1 _33085_ (.A1(_10587_),
    .A2(_10589_),
    .A3(_10590_),
    .ZN(_10591_));
 NOR4_X4 _33086_ (.A1(_07920_),
    .A2(_10583_),
    .A3(_10586_),
    .A4(_10591_),
    .ZN(_10592_));
 OAI21_X2 _33087_ (.A(_07684_),
    .B1(_07689_),
    .B2(_07427_),
    .ZN(_10593_));
 OAI221_X1 _33088_ (.A(_07391_),
    .B1(_07742_),
    .B2(_07621_),
    .C1(_07526_),
    .C2(_07524_),
    .ZN(_10594_));
 NAND2_X1 _33089_ (.A1(_07532_),
    .A2(_07476_),
    .ZN(_10595_));
 NAND4_X1 _33090_ (.A1(_07530_),
    .A2(_07829_),
    .A3(_10594_),
    .A4(_10595_),
    .ZN(_10596_));
 AOI22_X2 _33091_ (.A1(_07390_),
    .A2(_07482_),
    .B1(_07704_),
    .B2(_07368_),
    .ZN(_10597_));
 NAND3_X2 _33092_ (.A1(_08072_),
    .A2(_10596_),
    .A3(_10597_),
    .ZN(_10598_));
 AOI22_X4 _33093_ (.A1(_07474_),
    .A2(_07623_),
    .B1(_07688_),
    .B2(_07481_),
    .ZN(_10599_));
 AOI211_X2 _33094_ (.A(_07535_),
    .B(_07346_),
    .C1(_07531_),
    .C2(_07396_),
    .ZN(_10600_));
 NOR4_X2 _33095_ (.A1(_07397_),
    .A2(_07523_),
    .A3(_07454_),
    .A4(_07526_),
    .ZN(_10601_));
 NOR3_X2 _33096_ (.A1(_07544_),
    .A2(_10600_),
    .A3(_10601_),
    .ZN(_10602_));
 INV_X1 _33097_ (.A(_07379_),
    .ZN(_10603_));
 OAI22_X4 _33098_ (.A1(_07427_),
    .A2(_10599_),
    .B1(_10602_),
    .B2(_10603_),
    .ZN(_10604_));
 NOR4_X4 _33099_ (.A1(_07640_),
    .A2(_10593_),
    .A3(_10598_),
    .A4(_10604_),
    .ZN(_10605_));
 OAI221_X1 _33100_ (.A(_07436_),
    .B1(_07393_),
    .B2(_07458_),
    .C1(_07715_),
    .C2(_07682_),
    .ZN(_10606_));
 OAI221_X1 _33101_ (.A(_07432_),
    .B1(_07441_),
    .B2(_07392_),
    .C1(_07694_),
    .C2(_07476_),
    .ZN(_10607_));
 NAND3_X1 _33102_ (.A1(_07417_),
    .A2(_10606_),
    .A3(_10607_),
    .ZN(_10608_));
 OAI21_X1 _33103_ (.A(_07749_),
    .B1(_07710_),
    .B2(_07443_),
    .ZN(_10609_));
 AOI21_X2 _33104_ (.A(_07399_),
    .B1(_10608_),
    .B2(_10609_),
    .ZN(_10610_));
 NOR4_X4 _33105_ (.A1(_07821_),
    .A2(_07827_),
    .A3(_08133_),
    .A4(_10610_),
    .ZN(_10611_));
 NAND3_X4 _33106_ (.A1(_10592_),
    .A2(_10605_),
    .A3(_10611_),
    .ZN(_10612_));
 NOR3_X4 _33107_ (.A1(_07974_),
    .A2(_07982_),
    .A3(_10612_),
    .ZN(_10613_));
 OR2_X2 _33108_ (.A1(_06706_),
    .A2(_10613_),
    .ZN(_10614_));
 XNOR2_X1 _33109_ (.A(_07238_),
    .B(_00315_),
    .ZN(_10615_));
 XNOR2_X1 _33110_ (.A(_08998_),
    .B(_10615_),
    .ZN(_10616_));
 XNOR2_X1 _33111_ (.A(_07234_),
    .B(_10616_),
    .ZN(_10617_));
 MUX2_X1 _33112_ (.A(_07237_),
    .B(_10617_),
    .S(_09131_),
    .Z(_10618_));
 AOI22_X1 _33113_ (.A1(\block_reg[0][8] ),
    .A2(_09125_),
    .B1(_09126_),
    .B2(_10618_),
    .ZN(_10619_));
 OAI22_X1 _33114_ (.A1(\block_reg[0][8] ),
    .A2(_07904_),
    .B1(_09007_),
    .B2(_10618_),
    .ZN(_10620_));
 INV_X1 _33115_ (.A(_10620_),
    .ZN(_10621_));
 MUX2_X1 _33116_ (.A(_10619_),
    .B(_10621_),
    .S(_04326_),
    .Z(_10622_));
 NAND2_X1 _33117_ (.A1(_10614_),
    .A2(_10622_),
    .ZN(_10623_));
 CLKBUF_X3 _33118_ (.A(\core.enc_block.block_w0_reg[8] ),
    .Z(_10624_));
 MUX2_X1 _33119_ (.A(_10623_),
    .B(_10624_),
    .S(_08906_),
    .Z(_00732_));
 AND3_X1 _33120_ (.A1(_07484_),
    .A2(_07489_),
    .A3(_07616_),
    .ZN(_10625_));
 AOI21_X1 _33121_ (.A(_07445_),
    .B1(_10625_),
    .B2(_07447_),
    .ZN(_10626_));
 AOI21_X1 _33122_ (.A(_07975_),
    .B1(_07688_),
    .B2(_07507_),
    .ZN(_10627_));
 OAI221_X2 _33123_ (.A(_10587_),
    .B1(_10626_),
    .B2(_07663_),
    .C1(_10627_),
    .C2(_07447_),
    .ZN(_10628_));
 OAI21_X1 _33124_ (.A(_07487_),
    .B1(_07513_),
    .B2(_07547_),
    .ZN(_10629_));
 NAND3_X1 _33125_ (.A1(_07439_),
    .A2(_07362_),
    .A3(_10629_),
    .ZN(_10630_));
 AOI21_X1 _33126_ (.A(_07950_),
    .B1(_07853_),
    .B2(_07547_),
    .ZN(_10631_));
 OAI21_X2 _33127_ (.A(_10630_),
    .B1(_10631_),
    .B2(_07517_),
    .ZN(_10632_));
 AOI21_X1 _33128_ (.A(_07755_),
    .B1(_07545_),
    .B2(_07463_),
    .ZN(_10633_));
 NOR4_X1 _33129_ (.A1(_07532_),
    .A2(_07742_),
    .A3(_07522_),
    .A4(_07670_),
    .ZN(_10634_));
 NOR3_X1 _33130_ (.A1(_07439_),
    .A2(_07536_),
    .A3(_07621_),
    .ZN(_10635_));
 NOR3_X1 _33131_ (.A1(_07449_),
    .A2(_07530_),
    .A3(_07524_),
    .ZN(_10636_));
 OAI21_X1 _33132_ (.A(_10634_),
    .B1(_10635_),
    .B2(_10636_),
    .ZN(_10637_));
 NOR2_X1 _33133_ (.A1(_07532_),
    .A2(_07418_),
    .ZN(_10638_));
 OAI21_X1 _33134_ (.A(_07829_),
    .B1(_10638_),
    .B2(_07552_),
    .ZN(_10639_));
 NAND2_X1 _33135_ (.A1(_07532_),
    .A2(_07758_),
    .ZN(_10640_));
 XNOR2_X1 _33136_ (.A(_07448_),
    .B(_07535_),
    .ZN(_10641_));
 OR4_X1 _33137_ (.A1(_07522_),
    .A2(_10640_),
    .A3(_07670_),
    .A4(_10641_),
    .ZN(_10642_));
 NAND4_X2 _33138_ (.A1(_10633_),
    .A2(_10637_),
    .A3(_10639_),
    .A4(_10642_),
    .ZN(_10643_));
 NOR4_X2 _33139_ (.A1(_07595_),
    .A2(_07532_),
    .A3(_07621_),
    .A4(_07497_),
    .ZN(_10644_));
 AOI22_X2 _33140_ (.A1(_07596_),
    .A2(_07604_),
    .B1(_07977_),
    .B2(_10644_),
    .ZN(_10645_));
 NOR3_X1 _33141_ (.A1(_07543_),
    .A2(_07452_),
    .A3(_07499_),
    .ZN(_10646_));
 MUX2_X1 _33142_ (.A(_07758_),
    .B(_07848_),
    .S(_07536_),
    .Z(_10647_));
 AOI22_X2 _33143_ (.A1(_10641_),
    .A2(_10646_),
    .B1(_10647_),
    .B2(_07704_),
    .ZN(_10648_));
 OAI21_X2 _33144_ (.A(_10645_),
    .B1(_10648_),
    .B2(_07391_),
    .ZN(_10649_));
 NOR4_X4 _33145_ (.A1(_10628_),
    .A2(_10632_),
    .A3(_10643_),
    .A4(_10649_),
    .ZN(_10650_));
 NAND2_X1 _33146_ (.A1(_07777_),
    .A2(_07545_),
    .ZN(_10651_));
 AOI21_X1 _33147_ (.A(_07444_),
    .B1(_07976_),
    .B2(_10651_),
    .ZN(_10652_));
 NOR3_X2 _33148_ (.A1(_08157_),
    .A2(_08161_),
    .A3(_10652_),
    .ZN(_10653_));
 AOI22_X1 _33149_ (.A1(_07829_),
    .A2(_07545_),
    .B1(_07594_),
    .B2(_07868_),
    .ZN(_10654_));
 NAND2_X1 _33150_ (.A1(_07869_),
    .A2(_07870_),
    .ZN(_10655_));
 NAND2_X1 _33151_ (.A1(_10654_),
    .A2(_10655_),
    .ZN(_10656_));
 NOR4_X1 _33152_ (.A1(_07449_),
    .A2(_07455_),
    .A3(_07585_),
    .A4(_07582_),
    .ZN(_10657_));
 AOI21_X1 _33153_ (.A(_10657_),
    .B1(_07859_),
    .B2(_07369_),
    .ZN(_10658_));
 AOI21_X1 _33154_ (.A(_07447_),
    .B1(_07696_),
    .B2(_10658_),
    .ZN(_10659_));
 OAI21_X1 _33155_ (.A(_07707_),
    .B1(_07347_),
    .B2(_07443_),
    .ZN(_10660_));
 NAND2_X1 _33156_ (.A1(_07440_),
    .A2(_07443_),
    .ZN(_10661_));
 AOI21_X1 _33157_ (.A(_07543_),
    .B1(_10660_),
    .B2(_10661_),
    .ZN(_10662_));
 OAI33_X1 _33158_ (.A1(_07547_),
    .A2(_07586_),
    .A3(_07682_),
    .B1(_07474_),
    .B2(_07585_),
    .B3(_07455_),
    .ZN(_10663_));
 NAND2_X1 _33159_ (.A1(_07569_),
    .A2(_10663_),
    .ZN(_10664_));
 NAND4_X2 _33160_ (.A1(_07501_),
    .A2(_07673_),
    .A3(_07928_),
    .A4(_10664_),
    .ZN(_10665_));
 NOR4_X2 _33161_ (.A1(_10656_),
    .A2(_10659_),
    .A3(_10662_),
    .A4(_10665_),
    .ZN(_10666_));
 NOR2_X1 _33162_ (.A1(_07993_),
    .A2(_08084_),
    .ZN(_10667_));
 NAND4_X4 _33163_ (.A1(_10650_),
    .A2(_10653_),
    .A3(_10666_),
    .A4(_10667_),
    .ZN(_10668_));
 NOR2_X4 _33164_ (.A1(_07974_),
    .A2(_10668_),
    .ZN(_10669_));
 NOR2_X4 _33165_ (.A1(_06707_),
    .A2(_10669_),
    .ZN(_10670_));
 INV_X1 _33166_ (.A(_07645_),
    .ZN(_10671_));
 XNOR2_X1 _33167_ (.A(_10671_),
    .B(_08600_),
    .ZN(_10672_));
 XNOR2_X1 _33168_ (.A(_09001_),
    .B(_10672_),
    .ZN(_10673_));
 NAND2_X1 _33169_ (.A1(_08896_),
    .A2(_10673_),
    .ZN(_10674_));
 OAI21_X1 _33170_ (.A(_10674_),
    .B1(_10265_),
    .B2(_00312_),
    .ZN(_10675_));
 AOI22_X1 _33171_ (.A1(\block_reg[0][9] ),
    .A2(_07806_),
    .B1(_08599_),
    .B2(_10675_),
    .ZN(_10676_));
 INV_X1 _33172_ (.A(_10676_),
    .ZN(_10677_));
 CLKBUF_X3 _33173_ (.A(_07247_),
    .Z(_10678_));
 OAI22_X1 _33174_ (.A1(\block_reg[0][9] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_10675_),
    .ZN(_10679_));
 MUX2_X1 _33175_ (.A(_10677_),
    .B(_10679_),
    .S(_04563_),
    .Z(_10680_));
 NOR3_X2 _33176_ (.A1(_08906_),
    .A2(_10670_),
    .A3(_10680_),
    .ZN(_10681_));
 BUF_X2 _33177_ (.A(\core.enc_block.block_w0_reg[9] ),
    .Z(_10682_));
 INV_X1 _33178_ (.A(_10682_),
    .ZN(_10683_));
 AOI21_X1 _33179_ (.A(_10681_),
    .B1(_06705_),
    .B2(_10683_),
    .ZN(_00733_));
 AOI21_X4 _33180_ (.A(_06692_),
    .B1(_06698_),
    .B2(_06718_),
    .ZN(_10684_));
 BUF_X4 _33181_ (.A(_10684_),
    .Z(_10685_));
 CLKBUF_X3 _33182_ (.A(_10685_),
    .Z(_10686_));
 XNOR2_X2 _33183_ (.A(_09253_),
    .B(_09323_),
    .ZN(_10687_));
 XNOR2_X2 _33184_ (.A(_08178_),
    .B(\core.enc_block.block_w3_reg[8] ),
    .ZN(_10688_));
 XNOR2_X1 _33185_ (.A(_10687_),
    .B(_10688_),
    .ZN(_10689_));
 XNOR2_X1 _33186_ (.A(_10537_),
    .B(_10689_),
    .ZN(_10690_));
 NAND2_X1 _33187_ (.A1(_09217_),
    .A2(_10690_),
    .ZN(_10691_));
 OAI21_X2 _33188_ (.A(_10691_),
    .B1(_10172_),
    .B2(_06867_),
    .ZN(_10692_));
 OAI22_X1 _33189_ (.A1(\block_reg[1][0] ),
    .A2(_07905_),
    .B1(_08889_),
    .B2(_10692_),
    .ZN(_10693_));
 OR2_X1 _33190_ (.A1(_16490_),
    .A2(_10693_),
    .ZN(_10694_));
 CLKBUF_X3 _33191_ (.A(_09125_),
    .Z(_10695_));
 CLKBUF_X3 _33192_ (.A(_09126_),
    .Z(_10696_));
 AOI22_X1 _33193_ (.A1(\block_reg[1][0] ),
    .A2(_10695_),
    .B1(_10696_),
    .B2(_10692_),
    .ZN(_10697_));
 NAND2_X1 _33194_ (.A1(_16490_),
    .A2(_10697_),
    .ZN(_10698_));
 AOI21_X2 _33195_ (.A(_10685_),
    .B1(_10694_),
    .B2(_10698_),
    .ZN(_10699_));
 AOI22_X1 _33196_ (.A1(_06864_),
    .A2(_10686_),
    .B1(_10699_),
    .B2(_07223_),
    .ZN(_00734_));
 BUF_X4 _33197_ (.A(_07788_),
    .Z(_10700_));
 XNOR2_X1 _33198_ (.A(_08199_),
    .B(\core.enc_block.block_w0_reg[1] ),
    .ZN(_10701_));
 XNOR2_X1 _33199_ (.A(_09240_),
    .B(_10701_),
    .ZN(_10702_));
 XOR2_X1 _33200_ (.A(_07296_),
    .B(_10088_),
    .Z(_10703_));
 XNOR2_X1 _33201_ (.A(_10702_),
    .B(_10703_),
    .ZN(_10704_));
 NOR2_X1 _33202_ (.A1(_07902_),
    .A2(_10704_),
    .ZN(_10705_));
 AOI21_X4 _33203_ (.A(_10705_),
    .B1(_07902_),
    .B2(_00400_),
    .ZN(_10706_));
 BUF_X4 _33204_ (.A(_08888_),
    .Z(_10707_));
 OAI221_X2 _33205_ (.A(_05157_),
    .B1(_10700_),
    .B2(_10706_),
    .C1(_10707_),
    .C2(\block_reg[1][10] ),
    .ZN(_10708_));
 NAND2_X1 _33206_ (.A1(_00240_),
    .A2(_16549_),
    .ZN(_10709_));
 OAI21_X2 _33207_ (.A(_10709_),
    .B1(_05156_),
    .B2(_16549_),
    .ZN(_10710_));
 AOI22_X1 _33208_ (.A1(\block_reg[1][10] ),
    .A2(_10695_),
    .B1(_10696_),
    .B2(_10706_),
    .ZN(_10711_));
 NAND2_X1 _33209_ (.A1(_10710_),
    .A2(_10711_),
    .ZN(_10712_));
 AOI21_X2 _33210_ (.A(_10685_),
    .B1(_10708_),
    .B2(_10712_),
    .ZN(_10713_));
 AOI22_X1 _33211_ (.A1(_07277_),
    .A2(_10686_),
    .B1(_10713_),
    .B2(_07642_),
    .ZN(_00735_));
 CLKBUF_X3 _33212_ (.A(_10685_),
    .Z(_10714_));
 CLKBUF_X3 _33213_ (.A(_10684_),
    .Z(_10715_));
 CLKBUF_X3 _33214_ (.A(_07228_),
    .Z(_10716_));
 CLKBUF_X3 _33215_ (.A(_08038_),
    .Z(_10717_));
 XNOR2_X1 _33216_ (.A(_10537_),
    .B(_10088_),
    .ZN(_10718_));
 XNOR2_X1 _33217_ (.A(_09233_),
    .B(_08207_),
    .ZN(_10719_));
 XNOR2_X2 _33218_ (.A(_10718_),
    .B(_10719_),
    .ZN(_10720_));
 CLKBUF_X3 _33219_ (.A(\core.enc_block.block_w3_reg[10] ),
    .Z(_10721_));
 BUF_X4 _33220_ (.A(\core.enc_block.block_w3_reg[15] ),
    .Z(_10722_));
 XNOR2_X1 _33221_ (.A(_10274_),
    .B(_10722_),
    .ZN(_10723_));
 XNOR2_X1 _33222_ (.A(_10721_),
    .B(_10723_),
    .ZN(_10724_));
 XNOR2_X1 _33223_ (.A(_10720_),
    .B(_10724_),
    .ZN(_10725_));
 NAND2_X1 _33224_ (.A1(_10717_),
    .A2(_10725_),
    .ZN(_10726_));
 OAI21_X2 _33225_ (.A(_10726_),
    .B1(_07789_),
    .B2(_00403_),
    .ZN(_10727_));
 NAND2_X1 _33226_ (.A1(_10716_),
    .A2(_10727_),
    .ZN(_10728_));
 CLKBUF_X3 _33227_ (.A(_07247_),
    .Z(_10729_));
 INV_X1 _33228_ (.A(\block_reg[1][11] ),
    .ZN(_10730_));
 OAI21_X1 _33229_ (.A(_10728_),
    .B1(_10729_),
    .B2(_10730_),
    .ZN(_10731_));
 OAI22_X1 _33230_ (.A1(\block_reg[1][11] ),
    .A2(_10476_),
    .B1(_07788_),
    .B2(_10727_),
    .ZN(_10732_));
 MUX2_X1 _33231_ (.A(_10731_),
    .B(_10732_),
    .S(_05384_),
    .Z(_10733_));
 NOR2_X1 _33232_ (.A1(_10715_),
    .A2(_10733_),
    .ZN(_10734_));
 AOI22_X1 _33233_ (.A1(_07286_),
    .A2(_10714_),
    .B1(_10734_),
    .B2(_07786_),
    .ZN(_00736_));
 NOR2_X1 _33234_ (.A1(_07321_),
    .A2(_07231_),
    .ZN(_10735_));
 XNOR2_X1 _33235_ (.A(_10537_),
    .B(_10274_),
    .ZN(_10736_));
 XNOR2_X1 _33236_ (.A(_09285_),
    .B(_08218_),
    .ZN(_10737_));
 XNOR2_X2 _33237_ (.A(_10736_),
    .B(_10737_),
    .ZN(_10738_));
 BUF_X2 _33238_ (.A(\core.enc_block.block_w3_reg[11] ),
    .Z(_10739_));
 XNOR2_X2 _33239_ (.A(_10722_),
    .B(_10739_),
    .ZN(_10740_));
 XNOR2_X1 _33240_ (.A(_10368_),
    .B(_10740_),
    .ZN(_10741_));
 XNOR2_X2 _33241_ (.A(_10738_),
    .B(_10741_),
    .ZN(_10742_));
 AOI21_X4 _33242_ (.A(_10735_),
    .B1(_10742_),
    .B2(_07232_),
    .ZN(_10743_));
 AOI221_X2 _33243_ (.A(_05536_),
    .B1(_07228_),
    .B2(_10743_),
    .C1(_07805_),
    .C2(_06437_),
    .ZN(_10744_));
 NOR2_X1 _33244_ (.A1(_07788_),
    .A2(_10743_),
    .ZN(_10745_));
 AOI21_X1 _33245_ (.A(_10745_),
    .B1(_10695_),
    .B2(\block_reg[1][12] ),
    .ZN(_10746_));
 AOI21_X2 _33246_ (.A(_10744_),
    .B1(_10746_),
    .B2(_05536_),
    .ZN(_10747_));
 NOR2_X1 _33247_ (.A1(_10715_),
    .A2(_10747_),
    .ZN(_10748_));
 AOI22_X1 _33248_ (.A1(_07320_),
    .A2(_10714_),
    .B1(_10748_),
    .B2(_07892_),
    .ZN(_00737_));
 CLKBUF_X3 _33249_ (.A(_10684_),
    .Z(_10749_));
 INV_X1 _33250_ (.A(\block_reg[1][13] ),
    .ZN(_10750_));
 XNOR2_X2 _33251_ (.A(_09277_),
    .B(_08225_),
    .ZN(_10751_));
 XNOR2_X1 _33252_ (.A(_10368_),
    .B(_10751_),
    .ZN(_10752_));
 XNOR2_X1 _33253_ (.A(_07321_),
    .B(_10425_),
    .ZN(_10753_));
 XNOR2_X1 _33254_ (.A(_10752_),
    .B(_10753_),
    .ZN(_10754_));
 MUX2_X1 _33255_ (.A(_00386_),
    .B(_10754_),
    .S(_08809_),
    .Z(_10755_));
 OAI22_X1 _33256_ (.A1(_10750_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_10755_),
    .ZN(_10756_));
 NOR2_X1 _33257_ (.A1(_17061_),
    .A2(_10756_),
    .ZN(_10757_));
 AOI22_X1 _33258_ (.A1(_10750_),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_10755_),
    .ZN(_10758_));
 AOI21_X1 _33259_ (.A(_10757_),
    .B1(_10758_),
    .B2(_17061_),
    .ZN(_10759_));
 NOR2_X1 _33260_ (.A1(_10749_),
    .A2(_10759_),
    .ZN(_10760_));
 AOI22_X1 _33261_ (.A1(_07309_),
    .A2(_10714_),
    .B1(_10760_),
    .B2(_08037_),
    .ZN(_00738_));
 INV_X1 _33262_ (.A(\block_reg[1][14] ),
    .ZN(_10761_));
 XNOR2_X2 _33263_ (.A(_09260_),
    .B(_08243_),
    .ZN(_10762_));
 XNOR2_X2 _33264_ (.A(_10425_),
    .B(_10762_),
    .ZN(_10763_));
 XNOR2_X1 _33265_ (.A(_00386_),
    .B(_10482_),
    .ZN(_10764_));
 XNOR2_X1 _33266_ (.A(_10763_),
    .B(_10764_),
    .ZN(_10765_));
 MUX2_X1 _33267_ (.A(_00389_),
    .B(_10765_),
    .S(_08809_),
    .Z(_10766_));
 OAI22_X1 _33268_ (.A1(_10761_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_10766_),
    .ZN(_10767_));
 NOR2_X1 _33269_ (.A1(_03595_),
    .A2(_10767_),
    .ZN(_10768_));
 AOI22_X1 _33270_ (.A1(_10761_),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_10766_),
    .ZN(_10769_));
 AOI21_X2 _33271_ (.A(_10768_),
    .B1(_10769_),
    .B2(_03595_),
    .ZN(_10770_));
 NOR2_X1 _33272_ (.A1(_10749_),
    .A2(_10770_),
    .ZN(_10771_));
 AOI22_X1 _33273_ (.A1(_07332_),
    .A2(_10714_),
    .B1(_10771_),
    .B2(_08102_),
    .ZN(_00739_));
 INV_X1 _33274_ (.A(\block_reg[1][15] ),
    .ZN(_10772_));
 XNOR2_X2 _33275_ (.A(_09253_),
    .B(_08236_),
    .ZN(_10773_));
 XNOR2_X2 _33276_ (.A(_10482_),
    .B(_10773_),
    .ZN(_10774_));
 XNOR2_X1 _33277_ (.A(_00389_),
    .B(_10537_),
    .ZN(_10775_));
 XNOR2_X1 _33278_ (.A(_10774_),
    .B(_10775_),
    .ZN(_10776_));
 MUX2_X1 _33279_ (.A(_00392_),
    .B(_10776_),
    .S(_08809_),
    .Z(_10777_));
 OAI22_X1 _33280_ (.A1(_10772_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_10777_),
    .ZN(_10778_));
 NOR2_X1 _33281_ (.A1(_05114_),
    .A2(_10778_),
    .ZN(_10779_));
 AOI22_X1 _33282_ (.A1(_10772_),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_10777_),
    .ZN(_10780_));
 AOI21_X2 _33283_ (.A(_10779_),
    .B1(_10780_),
    .B2(_05114_),
    .ZN(_10781_));
 NOR2_X1 _33284_ (.A1(_10749_),
    .A2(_10781_),
    .ZN(_10782_));
 AOI22_X1 _33285_ (.A1(_07341_),
    .A2(_10714_),
    .B1(_10782_),
    .B2(_08164_),
    .ZN(_00740_));
 BUF_X4 _33286_ (.A(_10684_),
    .Z(_10783_));
 XNOR2_X2 _33287_ (.A(\core.enc_block.block_w3_reg[8] ),
    .B(_10722_),
    .ZN(_10784_));
 XOR2_X1 _33288_ (.A(_06867_),
    .B(_08236_),
    .Z(_10785_));
 XNOR2_X1 _33289_ (.A(_10784_),
    .B(_10785_),
    .ZN(_10786_));
 XNOR2_X1 _33290_ (.A(_09323_),
    .B(_10786_),
    .ZN(_10787_));
 MUX2_X1 _33291_ (.A(_08178_),
    .B(_10787_),
    .S(_07242_),
    .Z(_10788_));
 AOI22_X1 _33292_ (.A1(\block_reg[1][16] ),
    .A2(_07806_),
    .B1(_08599_),
    .B2(_10788_),
    .ZN(_10789_));
 INV_X1 _33293_ (.A(_10789_),
    .ZN(_10790_));
 OAI22_X1 _33294_ (.A1(\block_reg[1][16] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_10788_),
    .ZN(_10791_));
 MUX2_X1 _33295_ (.A(_10790_),
    .B(_10791_),
    .S(_17138_),
    .Z(_10792_));
 NOR3_X1 _33296_ (.A1(_08598_),
    .A2(_10783_),
    .A3(_10792_),
    .ZN(_10793_));
 AOI21_X1 _33297_ (.A(_10793_),
    .B1(_10686_),
    .B2(_08180_),
    .ZN(_00741_));
 CLKBUF_X3 _33298_ (.A(_07247_),
    .Z(_10794_));
 CLKBUF_X3 _33299_ (.A(_07253_),
    .Z(_10795_));
 BUF_X2 _33300_ (.A(\core.enc_block.block_w3_reg[9] ),
    .Z(_10796_));
 XOR2_X2 _33301_ (.A(_08178_),
    .B(_10796_),
    .Z(_10797_));
 XNOR2_X1 _33302_ (.A(_00363_),
    .B(_08236_),
    .ZN(_10798_));
 XNOR2_X2 _33303_ (.A(_10797_),
    .B(_10798_),
    .ZN(_10799_));
 XNOR2_X1 _33304_ (.A(_09312_),
    .B(_10784_),
    .ZN(_10800_));
 XNOR2_X2 _33305_ (.A(_10799_),
    .B(_10800_),
    .ZN(_10801_));
 MUX2_X2 _33306_ (.A(_08185_),
    .B(_10801_),
    .S(_07232_),
    .Z(_10802_));
 OAI22_X1 _33307_ (.A1(\block_reg[1][17] ),
    .A2(_10794_),
    .B1(_10795_),
    .B2(_10802_),
    .ZN(_10803_));
 NAND2_X1 _33308_ (.A1(_07908_),
    .A2(_10802_),
    .ZN(_10804_));
 OAI21_X1 _33309_ (.A(_10804_),
    .B1(_07787_),
    .B2(_06197_),
    .ZN(_10805_));
 MUX2_X1 _33310_ (.A(_10803_),
    .B(_10805_),
    .S(_03615_),
    .Z(_10806_));
 NOR2_X1 _33311_ (.A1(_10749_),
    .A2(_10806_),
    .ZN(_10807_));
 AOI22_X1 _33312_ (.A1(_08188_),
    .A2(_10714_),
    .B1(_10807_),
    .B2(_08716_),
    .ZN(_00742_));
 XOR2_X2 _33313_ (.A(_00366_),
    .B(_08185_),
    .Z(_10808_));
 XNOR2_X1 _33314_ (.A(_10721_),
    .B(_10796_),
    .ZN(_10809_));
 XNOR2_X1 _33315_ (.A(_10808_),
    .B(_10809_),
    .ZN(_10810_));
 XNOR2_X1 _33316_ (.A(_09240_),
    .B(_10810_),
    .ZN(_10811_));
 MUX2_X2 _33317_ (.A(_08199_),
    .B(_10811_),
    .S(_09131_),
    .Z(_10812_));
 AOI22_X1 _33318_ (.A1(\block_reg[1][18] ),
    .A2(_09125_),
    .B1(_09126_),
    .B2(_10812_),
    .ZN(_10813_));
 OAI22_X1 _33319_ (.A1(\block_reg[1][18] ),
    .A2(_07904_),
    .B1(_09007_),
    .B2(_10812_),
    .ZN(_10814_));
 INV_X1 _33320_ (.A(_10814_),
    .ZN(_10815_));
 MUX2_X1 _33321_ (.A(_10813_),
    .B(_10815_),
    .S(_05175_),
    .Z(_10816_));
 NAND2_X1 _33322_ (.A1(_08804_),
    .A2(_10816_),
    .ZN(_10817_));
 MUX2_X1 _33323_ (.A(_10817_),
    .B(_07644_),
    .S(_10783_),
    .Z(_00743_));
 XNOR2_X1 _33324_ (.A(_08236_),
    .B(_10740_),
    .ZN(_10818_));
 XNOR2_X1 _33325_ (.A(_00369_),
    .B(_08199_),
    .ZN(_10819_));
 XOR2_X1 _33326_ (.A(_09233_),
    .B(_10721_),
    .Z(_10820_));
 XNOR2_X1 _33327_ (.A(_10819_),
    .B(_10820_),
    .ZN(_10821_));
 XNOR2_X1 _33328_ (.A(_10818_),
    .B(_10821_),
    .ZN(_10822_));
 MUX2_X2 _33329_ (.A(_08207_),
    .B(_10822_),
    .S(_10265_),
    .Z(_10823_));
 OAI22_X1 _33330_ (.A1(\block_reg[1][19] ),
    .A2(_07905_),
    .B1(_08889_),
    .B2(_10823_),
    .ZN(_10824_));
 OR2_X1 _33331_ (.A1(_05405_),
    .A2(_10824_),
    .ZN(_10825_));
 AOI22_X1 _33332_ (.A1(\block_reg[1][19] ),
    .A2(_10695_),
    .B1(_10696_),
    .B2(_10823_),
    .ZN(_10826_));
 NAND2_X1 _33333_ (.A1(_05405_),
    .A2(_10826_),
    .ZN(_10827_));
 AOI21_X1 _33334_ (.A(_10685_),
    .B1(_10825_),
    .B2(_10827_),
    .ZN(_10828_));
 AOI22_X1 _33335_ (.A1(_08209_),
    .A2(_10714_),
    .B1(_10828_),
    .B2(_08887_),
    .ZN(_00744_));
 INV_X1 _33336_ (.A(\block_reg[1][1] ),
    .ZN(_10829_));
 XOR2_X2 _33337_ (.A(_10537_),
    .B(\core.enc_block.block_w0_reg[0] ),
    .Z(_10830_));
 XOR2_X1 _33338_ (.A(_09312_),
    .B(_08185_),
    .Z(_10831_));
 XNOR2_X1 _33339_ (.A(_10830_),
    .B(_10831_),
    .ZN(_10832_));
 XNOR2_X1 _33340_ (.A(_07296_),
    .B(_10687_),
    .ZN(_10833_));
 XNOR2_X1 _33341_ (.A(_10832_),
    .B(_10833_),
    .ZN(_10834_));
 MUX2_X2 _33342_ (.A(_00363_),
    .B(_10834_),
    .S(_08809_),
    .Z(_10835_));
 OAI22_X1 _33343_ (.A1(_10829_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_10835_),
    .ZN(_10836_));
 NOR2_X1 _33344_ (.A1(_03520_),
    .A2(_10836_),
    .ZN(_10837_));
 AOI22_X1 _33345_ (.A1(_10829_),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_10835_),
    .ZN(_10838_));
 AOI21_X2 _33346_ (.A(_10837_),
    .B1(_10838_),
    .B2(_03520_),
    .ZN(_10839_));
 NOR2_X1 _33347_ (.A1(_10749_),
    .A2(_10839_),
    .ZN(_10840_));
 AOI22_X1 _33348_ (.A1(_06803_),
    .A2(_10714_),
    .B1(_10840_),
    .B2(_08997_),
    .ZN(_00745_));
 CLKBUF_X2 _33349_ (.A(\core.enc_block.block_w3_reg[12] ),
    .Z(_10841_));
 XNOR2_X1 _33350_ (.A(_08207_),
    .B(_10841_),
    .ZN(_10842_));
 XNOR2_X1 _33351_ (.A(_00349_),
    .B(_00311_),
    .ZN(_10843_));
 XNOR2_X1 _33352_ (.A(_10842_),
    .B(_10843_),
    .ZN(_10844_));
 XNOR2_X1 _33353_ (.A(_10818_),
    .B(_10844_),
    .ZN(_10845_));
 MUX2_X1 _33354_ (.A(_08218_),
    .B(_10845_),
    .S(_08722_),
    .Z(_10846_));
 OAI221_X2 _33355_ (.A(_05523_),
    .B1(_10700_),
    .B2(_10846_),
    .C1(_10707_),
    .C2(\block_reg[1][20] ),
    .ZN(_10847_));
 NAND2_X1 _33356_ (.A1(_08901_),
    .A2(_10846_),
    .ZN(_10848_));
 INV_X1 _33357_ (.A(\block_reg[1][20] ),
    .ZN(_10849_));
 OAI21_X1 _33358_ (.A(_10848_),
    .B1(_08888_),
    .B2(_10849_),
    .ZN(_10850_));
 OR2_X1 _33359_ (.A1(_05523_),
    .A2(_10850_),
    .ZN(_10851_));
 AOI21_X2 _33360_ (.A(_10685_),
    .B1(_10847_),
    .B2(_10851_),
    .ZN(_10852_));
 AOI22_X1 _33361_ (.A1(_08220_),
    .A2(_10714_),
    .B1(_10852_),
    .B2(_09059_),
    .ZN(_00746_));
 XOR2_X2 _33362_ (.A(_00352_),
    .B(_08218_),
    .Z(_10853_));
 CLKBUF_X3 _33363_ (.A(\core.enc_block.block_w3_reg[13] ),
    .Z(_10854_));
 XNOR2_X1 _33364_ (.A(_10854_),
    .B(_10841_),
    .ZN(_10855_));
 XNOR2_X1 _33365_ (.A(_10853_),
    .B(_10855_),
    .ZN(_10856_));
 XNOR2_X1 _33366_ (.A(_09277_),
    .B(_10856_),
    .ZN(_10857_));
 MUX2_X1 _33367_ (.A(_08225_),
    .B(_10857_),
    .S(_08896_),
    .Z(_10858_));
 AOI22_X1 _33368_ (.A1(\block_reg[1][21] ),
    .A2(_09005_),
    .B1(_09211_),
    .B2(_10858_),
    .ZN(_10859_));
 NAND2_X1 _33369_ (.A1(_16942_),
    .A2(_10859_),
    .ZN(_10860_));
 OAI22_X1 _33370_ (.A1(\block_reg[1][21] ),
    .A2(_09221_),
    .B1(_09223_),
    .B2(_10858_),
    .ZN(_10861_));
 OAI21_X2 _33371_ (.A(_10860_),
    .B1(_10861_),
    .B2(_16942_),
    .ZN(_10862_));
 NAND2_X1 _33372_ (.A1(_09124_),
    .A2(_10862_),
    .ZN(_10863_));
 MUX2_X1 _33373_ (.A(_10863_),
    .B(_08040_),
    .S(_10783_),
    .Z(_00747_));
 INV_X1 _33374_ (.A(_09260_),
    .ZN(_10864_));
 BUF_X2 _33375_ (.A(\core.enc_block.block_w3_reg[14] ),
    .Z(_10865_));
 XNOR2_X1 _33376_ (.A(_00355_),
    .B(_10865_),
    .ZN(_10866_));
 XNOR2_X2 _33377_ (.A(_08225_),
    .B(_10854_),
    .ZN(_10867_));
 XNOR2_X1 _33378_ (.A(_10866_),
    .B(_10867_),
    .ZN(_10868_));
 XNOR2_X1 _33379_ (.A(_10864_),
    .B(_10868_),
    .ZN(_10869_));
 MUX2_X1 _33380_ (.A(_08243_),
    .B(_10869_),
    .S(_07651_),
    .Z(_10870_));
 OAI22_X1 _33381_ (.A1(\block_reg[1][22] ),
    .A2(_08104_),
    .B1(_09222_),
    .B2(_10870_),
    .ZN(_10871_));
 NOR2_X1 _33382_ (.A1(_16977_),
    .A2(_10871_),
    .ZN(_10872_));
 AOI22_X2 _33383_ (.A1(\block_reg[1][22] ),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_10870_),
    .ZN(_10873_));
 AOI21_X2 _33384_ (.A(_10872_),
    .B1(_10873_),
    .B2(_16977_),
    .ZN(_10874_));
 NOR3_X1 _33385_ (.A1(_09172_),
    .A2(_10783_),
    .A3(_10874_),
    .ZN(_10875_));
 AOI21_X1 _33386_ (.A(_10875_),
    .B1(_10686_),
    .B2(_08245_),
    .ZN(_00748_));
 XOR2_X2 _33387_ (.A(_00358_),
    .B(_10722_),
    .Z(_10876_));
 XNOR2_X1 _33388_ (.A(_08243_),
    .B(_10865_),
    .ZN(_10877_));
 XNOR2_X1 _33389_ (.A(_10876_),
    .B(_10877_),
    .ZN(_10878_));
 XNOR2_X1 _33390_ (.A(_09253_),
    .B(_10878_),
    .ZN(_10879_));
 MUX2_X1 _33391_ (.A(_08236_),
    .B(_10879_),
    .S(_08038_),
    .Z(_10880_));
 AOI22_X1 _33392_ (.A1(\block_reg[1][23] ),
    .A2(_09125_),
    .B1(_09126_),
    .B2(_10880_),
    .ZN(_10881_));
 OAI22_X1 _33393_ (.A1(\block_reg[1][23] ),
    .A2(_07904_),
    .B1(_09007_),
    .B2(_10880_),
    .ZN(_10882_));
 INV_X1 _33394_ (.A(_10882_),
    .ZN(_10883_));
 MUX2_X1 _33395_ (.A(_10881_),
    .B(_10883_),
    .S(_03626_),
    .Z(_10884_));
 NAND2_X1 _33396_ (.A1(_09210_),
    .A2(_10884_),
    .ZN(_10885_));
 MUX2_X1 _33397_ (.A(_10885_),
    .B(_08165_),
    .S(_10783_),
    .Z(_00749_));
 NOR2_X1 _33398_ (.A1(_09323_),
    .A2(_08896_),
    .ZN(_10886_));
 XNOR2_X2 _33399_ (.A(_10688_),
    .B(_10773_),
    .ZN(_10887_));
 XNOR2_X2 _33400_ (.A(_06867_),
    .B(_10887_),
    .ZN(_10888_));
 AOI21_X4 _33401_ (.A(_10886_),
    .B1(_10888_),
    .B2(_07789_),
    .ZN(_10889_));
 OAI22_X1 _33402_ (.A1(\block_reg[1][24] ),
    .A2(_10794_),
    .B1(_10795_),
    .B2(_10889_),
    .ZN(_10890_));
 CLKBUF_X3 _33403_ (.A(_07228_),
    .Z(_10891_));
 NAND2_X1 _33404_ (.A1(_10891_),
    .A2(_10889_),
    .ZN(_10892_));
 OAI21_X1 _33405_ (.A(_10892_),
    .B1(_07787_),
    .B2(_05959_),
    .ZN(_10893_));
 MUX2_X1 _33406_ (.A(_10890_),
    .B(_10893_),
    .S(_17096_),
    .Z(_10894_));
 NOR2_X1 _33407_ (.A1(_10749_),
    .A2(_10894_),
    .ZN(_10895_));
 AOI22_X1 _33408_ (.A1(_09324_),
    .A2(_10714_),
    .B1(_10895_),
    .B2(_09682_),
    .ZN(_00750_));
 XNOR2_X1 _33409_ (.A(_08185_),
    .B(_10687_),
    .ZN(_10896_));
 XNOR2_X2 _33410_ (.A(_10799_),
    .B(_10896_),
    .ZN(_10897_));
 MUX2_X1 _33411_ (.A(_09312_),
    .B(_10897_),
    .S(_08722_),
    .Z(_10898_));
 OAI221_X2 _33412_ (.A(_03555_),
    .B1(_10700_),
    .B2(_10898_),
    .C1(_10707_),
    .C2(\block_reg[1][25] ),
    .ZN(_10899_));
 NAND2_X1 _33413_ (.A1(_09211_),
    .A2(_10898_),
    .ZN(_10900_));
 INV_X1 _33414_ (.A(\block_reg[1][25] ),
    .ZN(_10901_));
 OAI21_X1 _33415_ (.A(_10900_),
    .B1(_08888_),
    .B2(_10901_),
    .ZN(_10902_));
 OR2_X1 _33416_ (.A1(_03555_),
    .A2(_10902_),
    .ZN(_10903_));
 AOI21_X2 _33417_ (.A(_10684_),
    .B1(_10899_),
    .B2(_10903_),
    .ZN(_10904_));
 AOI22_X1 _33418_ (.A1(_09313_),
    .A2(_10715_),
    .B1(_10904_),
    .B2(_09778_),
    .ZN(_00751_));
 CLKBUF_X3 _33419_ (.A(_07805_),
    .Z(_10905_));
 XNOR2_X2 _33420_ (.A(_09312_),
    .B(_10721_),
    .ZN(_10906_));
 XNOR2_X1 _33421_ (.A(_10808_),
    .B(_10906_),
    .ZN(_10907_));
 XNOR2_X1 _33422_ (.A(_08199_),
    .B(_10907_),
    .ZN(_10908_));
 MUX2_X1 _33423_ (.A(_09240_),
    .B(_10908_),
    .S(_09131_),
    .Z(_10909_));
 AOI22_X1 _33424_ (.A1(\block_reg[1][26] ),
    .A2(_10905_),
    .B1(_08599_),
    .B2(_10909_),
    .ZN(_10910_));
 INV_X1 _33425_ (.A(_10910_),
    .ZN(_10911_));
 OAI22_X1 _33426_ (.A1(\block_reg[1][26] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_10909_),
    .ZN(_10912_));
 MUX2_X1 _33427_ (.A(_10911_),
    .B(_10912_),
    .S(_05137_),
    .Z(_10913_));
 NOR3_X1 _33428_ (.A1(_09860_),
    .A2(_10783_),
    .A3(_10913_),
    .ZN(_10914_));
 INV_X1 _33429_ (.A(_09240_),
    .ZN(_10915_));
 AOI21_X1 _33430_ (.A(_10914_),
    .B1(_10686_),
    .B2(_10915_),
    .ZN(_00752_));
 XNOR2_X1 _33431_ (.A(_10773_),
    .B(_10819_),
    .ZN(_10916_));
 XNOR2_X1 _33432_ (.A(_08207_),
    .B(_10739_),
    .ZN(_10917_));
 XNOR2_X1 _33433_ (.A(_10915_),
    .B(_10917_),
    .ZN(_10918_));
 XNOR2_X1 _33434_ (.A(_10916_),
    .B(_10918_),
    .ZN(_10919_));
 MUX2_X1 _33435_ (.A(_09233_),
    .B(_10919_),
    .S(_09131_),
    .Z(_10920_));
 AOI22_X1 _33436_ (.A1(\block_reg[1][27] ),
    .A2(_10905_),
    .B1(_08599_),
    .B2(_10920_),
    .ZN(_10921_));
 INV_X1 _33437_ (.A(_10921_),
    .ZN(_10922_));
 OAI22_X1 _33438_ (.A1(\block_reg[1][27] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_10920_),
    .ZN(_10923_));
 MUX2_X1 _33439_ (.A(_10922_),
    .B(_10923_),
    .S(_05361_),
    .Z(_10924_));
 NOR3_X1 _33440_ (.A1(_09950_),
    .A2(_10783_),
    .A3(_10924_),
    .ZN(_10925_));
 AOI21_X1 _33441_ (.A(_10925_),
    .B1(_10686_),
    .B2(_09234_),
    .ZN(_00753_));
 XOR2_X1 _33442_ (.A(_10773_),
    .B(_10842_),
    .Z(_10926_));
 XNOR2_X1 _33443_ (.A(_08218_),
    .B(_10368_),
    .ZN(_10927_));
 XNOR2_X1 _33444_ (.A(_09234_),
    .B(_10927_),
    .ZN(_10928_));
 XNOR2_X1 _33445_ (.A(_10926_),
    .B(_10928_),
    .ZN(_10929_));
 NAND2_X1 _33446_ (.A1(_08809_),
    .A2(_10929_),
    .ZN(_10930_));
 OAI21_X2 _33447_ (.A(_10930_),
    .B1(_10265_),
    .B2(_00311_),
    .ZN(_10931_));
 AOI22_X1 _33448_ (.A1(\block_reg[1][28] ),
    .A2(_10905_),
    .B1(_08599_),
    .B2(_10931_),
    .ZN(_10932_));
 INV_X1 _33449_ (.A(_10932_),
    .ZN(_10933_));
 OAI22_X1 _33450_ (.A1(\block_reg[1][28] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_10931_),
    .ZN(_10934_));
 MUX2_X1 _33451_ (.A(_10933_),
    .B(_10934_),
    .S(_05509_),
    .Z(_10935_));
 NOR3_X1 _33452_ (.A1(_10010_),
    .A2(_10685_),
    .A3(_10935_),
    .ZN(_10936_));
 AOI21_X1 _33453_ (.A(_10936_),
    .B1(_10686_),
    .B2(_09286_),
    .ZN(_00754_));
 NOR2_X1 _33454_ (.A1(_09277_),
    .A2(_08896_),
    .ZN(_10937_));
 XNOR2_X1 _33455_ (.A(_10853_),
    .B(_10867_),
    .ZN(_10938_));
 XNOR2_X2 _33456_ (.A(_09286_),
    .B(_10938_),
    .ZN(_10939_));
 AOI21_X4 _33457_ (.A(_10937_),
    .B1(_10939_),
    .B2(_07789_),
    .ZN(_10940_));
 OAI22_X1 _33458_ (.A1(\block_reg[1][29] ),
    .A2(_10794_),
    .B1(_10795_),
    .B2(_10940_),
    .ZN(_10941_));
 NAND2_X1 _33459_ (.A1(_10891_),
    .A2(_10940_),
    .ZN(_10942_));
 OAI21_X1 _33460_ (.A(_10942_),
    .B1(_07787_),
    .B2(_06014_),
    .ZN(_10943_));
 MUX2_X1 _33461_ (.A(_10941_),
    .B(_10943_),
    .S(_17078_),
    .Z(_10944_));
 NOR2_X1 _33462_ (.A1(_10749_),
    .A2(_10944_),
    .ZN(_10945_));
 AOI22_X1 _33463_ (.A1(_09278_),
    .A2(_10715_),
    .B1(_10945_),
    .B2(_10076_),
    .ZN(_00755_));
 XNOR2_X1 _33464_ (.A(_10702_),
    .B(_10906_),
    .ZN(_10946_));
 NAND2_X1 _33465_ (.A1(_10354_),
    .A2(_10946_),
    .ZN(_10947_));
 BUF_X4 _33466_ (.A(_07651_),
    .Z(_10948_));
 OAI21_X2 _33467_ (.A(_10947_),
    .B1(_10948_),
    .B2(_00366_),
    .ZN(_10949_));
 OAI22_X1 _33468_ (.A1(\block_reg[1][2] ),
    .A2(_10794_),
    .B1(_10795_),
    .B2(_10949_),
    .ZN(_10950_));
 NAND2_X1 _33469_ (.A1(_10891_),
    .A2(_10949_),
    .ZN(_10951_));
 INV_X1 _33470_ (.A(\block_reg[1][2] ),
    .ZN(_10952_));
 OAI21_X1 _33471_ (.A(_10951_),
    .B1(_07787_),
    .B2(_10952_),
    .ZN(_10953_));
 MUX2_X1 _33472_ (.A(_10950_),
    .B(_10953_),
    .S(_05033_),
    .Z(_10954_));
 NOR2_X1 _33473_ (.A1(_10749_),
    .A2(_10954_),
    .ZN(_10955_));
 AOI22_X1 _33474_ (.A1(_06791_),
    .A2(_10715_),
    .B1(_10955_),
    .B2(_10168_),
    .ZN(_00756_));
 CLKBUF_X3 _33475_ (.A(_07227_),
    .Z(_10956_));
 INV_X1 _33476_ (.A(_08243_),
    .ZN(_10957_));
 XNOR2_X1 _33477_ (.A(_10751_),
    .B(_10866_),
    .ZN(_10958_));
 XNOR2_X1 _33478_ (.A(_10957_),
    .B(_10958_),
    .ZN(_10959_));
 MUX2_X1 _33479_ (.A(_09260_),
    .B(_10959_),
    .S(_09131_),
    .Z(_10960_));
 AOI22_X1 _33480_ (.A1(\block_reg[1][30] ),
    .A2(_10905_),
    .B1(_10956_),
    .B2(_10960_),
    .ZN(_10961_));
 INV_X1 _33481_ (.A(_10961_),
    .ZN(_10962_));
 OAI22_X1 _33482_ (.A1(\block_reg[1][30] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_10960_),
    .ZN(_10963_));
 MUX2_X1 _33483_ (.A(_10962_),
    .B(_10963_),
    .S(_03540_),
    .Z(_10964_));
 NOR3_X1 _33484_ (.A1(_10222_),
    .A2(_10685_),
    .A3(_10964_),
    .ZN(_10965_));
 AOI21_X1 _33485_ (.A(_10965_),
    .B1(_10686_),
    .B2(_10864_),
    .ZN(_00757_));
 INV_X1 _33486_ (.A(_08236_),
    .ZN(_10966_));
 XOR2_X1 _33487_ (.A(_10762_),
    .B(_10876_),
    .Z(_10967_));
 XNOR2_X1 _33488_ (.A(_10966_),
    .B(_10967_),
    .ZN(_10968_));
 MUX2_X1 _33489_ (.A(_09253_),
    .B(_10968_),
    .S(_07651_),
    .Z(_10969_));
 OAI22_X1 _33490_ (.A1(\block_reg[1][31] ),
    .A2(_09134_),
    .B1(_09222_),
    .B2(_10969_),
    .ZN(_10970_));
 NOR2_X1 _33491_ (.A1(_17168_),
    .A2(_10970_),
    .ZN(_10971_));
 AOI22_X1 _33492_ (.A1(\block_reg[1][31] ),
    .A2(_08116_),
    .B1(_08901_),
    .B2(_10969_),
    .ZN(_10972_));
 AOI21_X1 _33493_ (.A(_10971_),
    .B1(_10972_),
    .B2(_17168_),
    .ZN(_10973_));
 NOR3_X1 _33494_ (.A1(_10261_),
    .A2(_10685_),
    .A3(_10973_),
    .ZN(_10974_));
 INV_X1 _33495_ (.A(_09253_),
    .ZN(_10975_));
 AOI21_X1 _33496_ (.A(_10974_),
    .B1(_10686_),
    .B2(_10975_),
    .ZN(_00758_));
 XNOR2_X1 _33497_ (.A(_09240_),
    .B(_00403_),
    .ZN(_10976_));
 XNOR2_X1 _33498_ (.A(_10975_),
    .B(_10976_),
    .ZN(_10977_));
 XNOR2_X1 _33499_ (.A(_10720_),
    .B(_10977_),
    .ZN(_10978_));
 NAND2_X1 _33500_ (.A1(_07801_),
    .A2(_10978_),
    .ZN(_10979_));
 OAI21_X2 _33501_ (.A(_10979_),
    .B1(_10172_),
    .B2(_00369_),
    .ZN(_10980_));
 OAI221_X2 _33502_ (.A(_05282_),
    .B1(_10700_),
    .B2(_10980_),
    .C1(_10707_),
    .C2(\block_reg[1][3] ),
    .ZN(_10981_));
 AOI22_X1 _33503_ (.A1(\block_reg[1][3] ),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_10980_),
    .ZN(_10982_));
 OAI21_X1 _33504_ (.A(_10982_),
    .B1(_05281_),
    .B2(_05269_),
    .ZN(_10983_));
 AOI21_X2 _33505_ (.A(_10684_),
    .B1(_10981_),
    .B2(_10983_),
    .ZN(_10984_));
 AOI22_X1 _33506_ (.A1(_06722_),
    .A2(_10715_),
    .B1(_10984_),
    .B2(_10353_),
    .ZN(_00759_));
 XNOR2_X1 _33507_ (.A(_09233_),
    .B(_07321_),
    .ZN(_10985_));
 XNOR2_X1 _33508_ (.A(_10975_),
    .B(_10985_),
    .ZN(_10986_));
 XNOR2_X1 _33509_ (.A(_10738_),
    .B(_10986_),
    .ZN(_10987_));
 NAND2_X1 _33510_ (.A1(_10354_),
    .A2(_10987_),
    .ZN(_10988_));
 OAI21_X2 _33511_ (.A(_10988_),
    .B1(_10948_),
    .B2(_00349_),
    .ZN(_10989_));
 OAI22_X1 _33512_ (.A1(\block_reg[1][4] ),
    .A2(_10794_),
    .B1(_10795_),
    .B2(_10989_),
    .ZN(_10990_));
 NAND2_X1 _33513_ (.A1(_10891_),
    .A2(_10989_),
    .ZN(_10991_));
 CLKBUF_X3 _33514_ (.A(_07247_),
    .Z(_10992_));
 INV_X1 _33515_ (.A(\block_reg[1][4] ),
    .ZN(_10993_));
 OAI21_X1 _33516_ (.A(_10991_),
    .B1(_10992_),
    .B2(_10993_),
    .ZN(_10994_));
 MUX2_X1 _33517_ (.A(_10990_),
    .B(_10994_),
    .S(_05488_),
    .Z(_10995_));
 NOR2_X1 _33518_ (.A1(_10749_),
    .A2(_10995_),
    .ZN(_10996_));
 AOI22_X1 _33519_ (.A1(_06771_),
    .A2(_10715_),
    .B1(_10996_),
    .B2(_10414_),
    .ZN(_00760_));
 XNOR2_X1 _33520_ (.A(_09285_),
    .B(_10854_),
    .ZN(_10997_));
 XNOR2_X1 _33521_ (.A(_10752_),
    .B(_10997_),
    .ZN(_10998_));
 NAND2_X1 _33522_ (.A1(_10717_),
    .A2(_10998_),
    .ZN(_10999_));
 OAI21_X2 _33523_ (.A(_10999_),
    .B1(_07789_),
    .B2(_00352_),
    .ZN(_11000_));
 NAND2_X1 _33524_ (.A1(_10716_),
    .A2(_11000_),
    .ZN(_11001_));
 INV_X1 _33525_ (.A(\block_reg[1][5] ),
    .ZN(_11002_));
 OAI21_X1 _33526_ (.A(_11001_),
    .B1(_10729_),
    .B2(_11002_),
    .ZN(_11003_));
 OAI22_X1 _33527_ (.A1(\block_reg[1][5] ),
    .A2(_10476_),
    .B1(_07788_),
    .B2(_11000_),
    .ZN(_11004_));
 MUX2_X1 _33528_ (.A(_11003_),
    .B(_11004_),
    .S(_17197_),
    .Z(_11005_));
 NOR2_X1 _33529_ (.A1(_10749_),
    .A2(_11005_),
    .ZN(_11006_));
 AOI22_X1 _33530_ (.A1(_06764_),
    .A2(_10715_),
    .B1(_11006_),
    .B2(_10470_),
    .ZN(_00761_));
 XNOR2_X1 _33531_ (.A(_09277_),
    .B(_10865_),
    .ZN(_11007_));
 XNOR2_X1 _33532_ (.A(_10763_),
    .B(_11007_),
    .ZN(_11008_));
 NAND2_X1 _33533_ (.A1(_10717_),
    .A2(_11008_),
    .ZN(_11009_));
 OAI21_X2 _33534_ (.A(_11009_),
    .B1(_07789_),
    .B2(_00355_),
    .ZN(_11010_));
 NAND2_X1 _33535_ (.A1(_10716_),
    .A2(_11010_),
    .ZN(_11011_));
 INV_X1 _33536_ (.A(\block_reg[1][6] ),
    .ZN(_11012_));
 OAI21_X1 _33537_ (.A(_11011_),
    .B1(_10729_),
    .B2(_11012_),
    .ZN(_11013_));
 OAI22_X1 _33538_ (.A1(\block_reg[1][6] ),
    .A2(_10476_),
    .B1(_07788_),
    .B2(_11010_),
    .ZN(_11014_));
 MUX2_X1 _33539_ (.A(_11013_),
    .B(_11014_),
    .S(_16874_),
    .Z(_11015_));
 NOR2_X1 _33540_ (.A1(_10783_),
    .A2(_11015_),
    .ZN(_11016_));
 AOI22_X1 _33541_ (.A1(_06752_),
    .A2(_10715_),
    .B1(_11016_),
    .B2(_10527_),
    .ZN(_00762_));
 CLKBUF_X3 _33542_ (.A(_07253_),
    .Z(_11017_));
 XNOR2_X1 _33543_ (.A(_09260_),
    .B(_10722_),
    .ZN(_11018_));
 XNOR2_X1 _33544_ (.A(_10774_),
    .B(_11018_),
    .ZN(_11019_));
 NAND2_X1 _33545_ (.A1(_10354_),
    .A2(_11019_),
    .ZN(_11020_));
 OAI21_X2 _33546_ (.A(_11020_),
    .B1(_10948_),
    .B2(_00358_),
    .ZN(_11021_));
 OAI22_X1 _33547_ (.A1(\block_reg[1][7] ),
    .A2(_10794_),
    .B1(_11017_),
    .B2(_11021_),
    .ZN(_11022_));
 NAND2_X1 _33548_ (.A1(_10891_),
    .A2(_11021_),
    .ZN(_11023_));
 OAI21_X1 _33549_ (.A(_11023_),
    .B1(_10992_),
    .B2(_05675_),
    .ZN(_11024_));
 MUX2_X2 _33550_ (.A(_11022_),
    .B(_11024_),
    .S(_17184_),
    .Z(_11025_));
 NOR2_X1 _33551_ (.A1(_10783_),
    .A2(_11025_),
    .ZN(_11026_));
 AOI22_X1 _33552_ (.A1(_06741_),
    .A2(_10715_),
    .B1(_11026_),
    .B2(_10566_),
    .ZN(_00763_));
 XNOR2_X1 _33553_ (.A(_00392_),
    .B(_08178_),
    .ZN(_11027_));
 XNOR2_X1 _33554_ (.A(_10830_),
    .B(_11027_),
    .ZN(_11028_));
 XNOR2_X1 _33555_ (.A(_09323_),
    .B(_11028_),
    .ZN(_11029_));
 NAND2_X1 _33556_ (.A1(_10354_),
    .A2(_11029_),
    .ZN(_11030_));
 OAI21_X2 _33557_ (.A(_11030_),
    .B1(_07801_),
    .B2(_00394_),
    .ZN(_11031_));
 AOI22_X1 _33558_ (.A1(\block_reg[1][8] ),
    .A2(_09005_),
    .B1(_07908_),
    .B2(_11031_),
    .ZN(_11032_));
 NAND2_X1 _33559_ (.A1(_17011_),
    .A2(_11032_),
    .ZN(_11033_));
 OAI22_X1 _33560_ (.A1(\block_reg[1][8] ),
    .A2(_09221_),
    .B1(_09223_),
    .B2(_11031_),
    .ZN(_11034_));
 OAI21_X1 _33561_ (.A(_11033_),
    .B1(_11034_),
    .B2(_17011_),
    .ZN(_11035_));
 NAND2_X1 _33562_ (.A1(_10614_),
    .A2(_11035_),
    .ZN(_11036_));
 MUX2_X1 _33563_ (.A(_11036_),
    .B(_07267_),
    .S(_10783_),
    .Z(_00764_));
 XNOR2_X1 _33564_ (.A(\core.enc_block.block_w0_reg[1] ),
    .B(_10784_),
    .ZN(_11037_));
 XNOR2_X1 _33565_ (.A(_10832_),
    .B(_11037_),
    .ZN(_11038_));
 NAND2_X1 _33566_ (.A1(_08039_),
    .A2(_11038_),
    .ZN(_11039_));
 OAI21_X2 _33567_ (.A(_11039_),
    .B1(_07243_),
    .B2(_07296_),
    .ZN(_11040_));
 OAI22_X1 _33568_ (.A1(\block_reg[1][9] ),
    .A2(_09134_),
    .B1(_09222_),
    .B2(_11040_),
    .ZN(_11041_));
 NOR2_X1 _33569_ (.A1(_03574_),
    .A2(_11041_),
    .ZN(_11042_));
 AOI22_X1 _33570_ (.A1(\block_reg[1][9] ),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_11040_),
    .ZN(_11043_));
 AOI21_X1 _33571_ (.A(_11042_),
    .B1(_11043_),
    .B2(_03574_),
    .ZN(_11044_));
 NOR3_X1 _33572_ (.A1(_10670_),
    .A2(_10685_),
    .A3(_11044_),
    .ZN(_11045_));
 AOI21_X1 _33573_ (.A(_11045_),
    .B1(_10686_),
    .B2(_07295_),
    .ZN(_00765_));
 INV_X1 _33574_ (.A(_06861_),
    .ZN(_11046_));
 AOI21_X4 _33575_ (.A(_06692_),
    .B1(_07260_),
    .B2(_07264_),
    .ZN(_11047_));
 BUF_X4 _33576_ (.A(_11047_),
    .Z(_11048_));
 BUF_X4 _33577_ (.A(_11048_),
    .Z(_11049_));
 NOR2_X1 _33578_ (.A1(_06863_),
    .A2(_07789_),
    .ZN(_11050_));
 XNOR2_X2 _33579_ (.A(_09255_),
    .B(_09321_),
    .ZN(_11051_));
 BUF_X2 _33580_ (.A(\core.enc_block.block_w3_reg[16] ),
    .Z(_11052_));
 XNOR2_X2 _33581_ (.A(_11052_),
    .B(_10624_),
    .ZN(_11053_));
 XNOR2_X1 _33582_ (.A(_11051_),
    .B(_11053_),
    .ZN(_11054_));
 XNOR2_X2 _33583_ (.A(_00308_),
    .B(_11054_),
    .ZN(_11055_));
 AOI21_X4 _33584_ (.A(_11050_),
    .B1(_11055_),
    .B2(_10172_),
    .ZN(_11056_));
 OAI221_X2 _33585_ (.A(_17778_),
    .B1(_10700_),
    .B2(_11056_),
    .C1(_10707_),
    .C2(\block_reg[2][0] ),
    .ZN(_11057_));
 AOI22_X2 _33586_ (.A1(\block_reg[2][0] ),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_11056_),
    .ZN(_11058_));
 OAI21_X2 _33587_ (.A(_11058_),
    .B1(_17777_),
    .B2(_17776_),
    .ZN(_11059_));
 AOI21_X2 _33588_ (.A(_11048_),
    .B1(_11057_),
    .B2(_11059_),
    .ZN(_11060_));
 AOI22_X1 _33589_ (.A1(_11046_),
    .A2(_11049_),
    .B1(_11060_),
    .B2(_07223_),
    .ZN(_00766_));
 INV_X1 _33590_ (.A(_07274_),
    .ZN(_11061_));
 CLKBUF_X3 _33591_ (.A(_11047_),
    .Z(_11062_));
 XOR2_X2 _33592_ (.A(_09243_),
    .B(_06790_),
    .Z(_11063_));
 BUF_X2 _33593_ (.A(\core.enc_block.block_w3_reg[18] ),
    .Z(_11064_));
 XNOR2_X1 _33594_ (.A(_07298_),
    .B(_11064_),
    .ZN(_11065_));
 XNOR2_X1 _33595_ (.A(_11063_),
    .B(_11065_),
    .ZN(_11066_));
 XNOR2_X1 _33596_ (.A(_06802_),
    .B(_11066_),
    .ZN(_11067_));
 NAND2_X1 _33597_ (.A1(_10354_),
    .A2(_11067_),
    .ZN(_11068_));
 OAI21_X4 _33598_ (.A(_11068_),
    .B1(_10948_),
    .B2(_00399_),
    .ZN(_11069_));
 OAI22_X1 _33599_ (.A1(\block_reg[2][10] ),
    .A2(_10794_),
    .B1(_11017_),
    .B2(_11069_),
    .ZN(_11070_));
 NAND2_X1 _33600_ (.A1(_10891_),
    .A2(_11069_),
    .ZN(_11071_));
 OAI21_X1 _33601_ (.A(_11071_),
    .B1(_10992_),
    .B2(_17711_),
    .ZN(_11072_));
 MUX2_X1 _33602_ (.A(_11070_),
    .B(_11072_),
    .S(_17727_),
    .Z(_11073_));
 NOR2_X1 _33603_ (.A1(_11062_),
    .A2(_11073_),
    .ZN(_11074_));
 AOI22_X1 _33604_ (.A1(_11061_),
    .A2(_11049_),
    .B1(_11074_),
    .B2(_07642_),
    .ZN(_00767_));
 INV_X1 _33605_ (.A(_07283_),
    .ZN(_11075_));
 CLKBUF_X3 _33606_ (.A(_11048_),
    .Z(_11076_));
 XNOR2_X1 _33607_ (.A(_06721_),
    .B(_07258_),
    .ZN(_11077_));
 XNOR2_X1 _33608_ (.A(_09231_),
    .B(_11077_),
    .ZN(_11078_));
 XNOR2_X2 _33609_ (.A(_06740_),
    .B(_08121_),
    .ZN(_11079_));
 CLKBUF_X3 _33610_ (.A(\core.enc_block.block_w3_reg[19] ),
    .Z(_11080_));
 XNOR2_X1 _33611_ (.A(_06790_),
    .B(_11080_),
    .ZN(_11081_));
 XNOR2_X1 _33612_ (.A(_11079_),
    .B(_11081_),
    .ZN(_11082_));
 XNOR2_X1 _33613_ (.A(_11078_),
    .B(_11082_),
    .ZN(_11083_));
 NAND2_X1 _33614_ (.A1(_10717_),
    .A2(_11083_),
    .ZN(_11084_));
 OAI21_X2 _33615_ (.A(_11084_),
    .B1(_10948_),
    .B2(_00402_),
    .ZN(_11085_));
 OAI22_X1 _33616_ (.A1(\block_reg[2][11] ),
    .A2(_10794_),
    .B1(_11017_),
    .B2(_11085_),
    .ZN(_11086_));
 NAND2_X1 _33617_ (.A1(_10891_),
    .A2(_11085_),
    .ZN(_11087_));
 OAI21_X1 _33618_ (.A(_11087_),
    .B1(_10992_),
    .B2(_18065_),
    .ZN(_11088_));
 MUX2_X1 _33619_ (.A(_11086_),
    .B(_11088_),
    .S(_18076_),
    .Z(_11089_));
 NOR2_X1 _33620_ (.A1(_11062_),
    .A2(_11089_),
    .ZN(_11090_));
 AOI22_X1 _33621_ (.A1(_11075_),
    .A2(_11076_),
    .B1(_11090_),
    .B2(_07786_),
    .ZN(_00768_));
 INV_X1 _33622_ (.A(_07317_),
    .ZN(_11091_));
 OR2_X1 _33623_ (.A1(_07323_),
    .A2(_07242_),
    .ZN(_11092_));
 XNOR2_X2 _33624_ (.A(\core.enc_block.block_w2_reg[28] ),
    .B(\core.enc_block.block_w3_reg[20] ),
    .ZN(_11093_));
 XOR2_X2 _33625_ (.A(_06740_),
    .B(_06721_),
    .Z(_11094_));
 XNOR2_X2 _33626_ (.A(_11093_),
    .B(_11094_),
    .ZN(_11095_));
 XNOR2_X2 _33627_ (.A(_08121_),
    .B(_07659_),
    .ZN(_11096_));
 XNOR2_X1 _33628_ (.A(_06770_),
    .B(_11096_),
    .ZN(_11097_));
 XNOR2_X1 _33629_ (.A(_11095_),
    .B(_11097_),
    .ZN(_11098_));
 OAI21_X2 _33630_ (.A(_11092_),
    .B1(_11098_),
    .B2(_07902_),
    .ZN(_11099_));
 OAI22_X1 _33631_ (.A1(\block_reg[2][12] ),
    .A2(_10232_),
    .B1(_11017_),
    .B2(_11099_),
    .ZN(_11100_));
 NAND2_X1 _33632_ (.A1(_10891_),
    .A2(_11099_),
    .ZN(_11101_));
 INV_X1 _33633_ (.A(\block_reg[2][12] ),
    .ZN(_11102_));
 OAI21_X1 _33634_ (.A(_11101_),
    .B1(_10992_),
    .B2(_11102_),
    .ZN(_11103_));
 MUX2_X1 _33635_ (.A(_11100_),
    .B(_11103_),
    .S(_18240_),
    .Z(_11104_));
 NOR2_X1 _33636_ (.A1(_11062_),
    .A2(_11104_),
    .ZN(_11105_));
 AOI22_X1 _33637_ (.A1(_11091_),
    .A2(_11076_),
    .B1(_11105_),
    .B2(_07892_),
    .ZN(_00769_));
 INV_X1 _33638_ (.A(_07306_),
    .ZN(_11106_));
 CLKBUF_X3 _33639_ (.A(_11047_),
    .Z(_11107_));
 XOR2_X2 _33640_ (.A(_09275_),
    .B(_06763_),
    .Z(_11108_));
 CLKBUF_X3 _33641_ (.A(\core.enc_block.block_w3_reg[21] ),
    .Z(_11109_));
 XNOR2_X1 _33642_ (.A(_07323_),
    .B(_11109_),
    .ZN(_11110_));
 XNOR2_X1 _33643_ (.A(_11108_),
    .B(_11110_),
    .ZN(_11111_));
 XNOR2_X1 _33644_ (.A(_06770_),
    .B(_11111_),
    .ZN(_11112_));
 NAND2_X1 _33645_ (.A1(_10717_),
    .A2(_11112_),
    .ZN(_11113_));
 OAI21_X2 _33646_ (.A(_11113_),
    .B1(_07789_),
    .B2(_00385_),
    .ZN(_11114_));
 NAND2_X1 _33647_ (.A1(_10716_),
    .A2(_11114_),
    .ZN(_11115_));
 INV_X1 _33648_ (.A(\block_reg[2][13] ),
    .ZN(_11116_));
 OAI21_X1 _33649_ (.A(_11115_),
    .B1(_10729_),
    .B2(_11116_),
    .ZN(_11117_));
 OAI22_X1 _33650_ (.A1(\block_reg[2][13] ),
    .A2(_10476_),
    .B1(_07788_),
    .B2(_11114_),
    .ZN(_11118_));
 MUX2_X1 _33651_ (.A(_11117_),
    .B(_11118_),
    .S(_17823_),
    .Z(_11119_));
 NOR2_X1 _33652_ (.A1(_11107_),
    .A2(_11119_),
    .ZN(_11120_));
 AOI22_X1 _33653_ (.A1(_11106_),
    .A2(_11076_),
    .B1(_11120_),
    .B2(_08037_),
    .ZN(_00770_));
 INV_X1 _33654_ (.A(_07329_),
    .ZN(_11121_));
 XNOR2_X2 _33655_ (.A(_09262_),
    .B(_06751_),
    .ZN(_11122_));
 CLKBUF_X3 _33656_ (.A(\core.enc_block.block_w3_reg[22] ),
    .Z(_11123_));
 XOR2_X1 _33657_ (.A(_00385_),
    .B(_11123_),
    .Z(_11124_));
 XNOR2_X1 _33658_ (.A(_11122_),
    .B(_11124_),
    .ZN(_11125_));
 XNOR2_X1 _33659_ (.A(_06763_),
    .B(_11125_),
    .ZN(_11126_));
 NAND2_X1 _33660_ (.A1(_10354_),
    .A2(_11126_),
    .ZN(_11127_));
 OAI21_X2 _33661_ (.A(_11127_),
    .B1(_07801_),
    .B2(_00388_),
    .ZN(_11128_));
 OAI221_X1 _33662_ (.A(_17701_),
    .B1(_10700_),
    .B2(_11128_),
    .C1(_10707_),
    .C2(\block_reg[2][14] ),
    .ZN(_11129_));
 NAND2_X1 _33663_ (.A1(_09211_),
    .A2(_11128_),
    .ZN(_11130_));
 INV_X1 _33664_ (.A(\block_reg[2][14] ),
    .ZN(_11131_));
 OAI21_X1 _33665_ (.A(_11130_),
    .B1(_08888_),
    .B2(_11131_),
    .ZN(_11132_));
 OR2_X1 _33666_ (.A1(_17701_),
    .A2(_11132_),
    .ZN(_11133_));
 AOI21_X1 _33667_ (.A(_11048_),
    .B1(_11129_),
    .B2(_11133_),
    .ZN(_11134_));
 AOI22_X1 _33668_ (.A1(_11121_),
    .A2(_11076_),
    .B1(_11134_),
    .B2(_08102_),
    .ZN(_00771_));
 INV_X1 _33669_ (.A(_07338_),
    .ZN(_11135_));
 BUF_X4 _33670_ (.A(\core.enc_block.block_w3_reg[23] ),
    .Z(_11136_));
 XOR2_X2 _33671_ (.A(_09255_),
    .B(_11136_),
    .Z(_11137_));
 XNOR2_X1 _33672_ (.A(_06740_),
    .B(_00388_),
    .ZN(_11138_));
 XNOR2_X1 _33673_ (.A(_11137_),
    .B(_11138_),
    .ZN(_11139_));
 XNOR2_X1 _33674_ (.A(_06751_),
    .B(_11139_),
    .ZN(_11140_));
 NAND2_X1 _33675_ (.A1(_10265_),
    .A2(_11140_),
    .ZN(_11141_));
 OAI21_X2 _33676_ (.A(_11141_),
    .B1(_07789_),
    .B2(_00391_),
    .ZN(_11142_));
 NAND2_X1 _33677_ (.A1(_09126_),
    .A2(_11142_),
    .ZN(_11143_));
 INV_X1 _33678_ (.A(\block_reg[2][15] ),
    .ZN(_11144_));
 OAI21_X1 _33679_ (.A(_11143_),
    .B1(_10729_),
    .B2(_11144_),
    .ZN(_11145_));
 OAI22_X1 _33680_ (.A1(\block_reg[2][15] ),
    .A2(_10476_),
    .B1(_10795_),
    .B2(_11142_),
    .ZN(_11146_));
 MUX2_X1 _33681_ (.A(_11145_),
    .B(_11146_),
    .S(_17847_),
    .Z(_11147_));
 NOR2_X1 _33682_ (.A1(_11107_),
    .A2(_11147_),
    .ZN(_11148_));
 AOI22_X1 _33683_ (.A1(_11135_),
    .A2(_11076_),
    .B1(_11148_),
    .B2(_08164_),
    .ZN(_00772_));
 BUF_X4 _33684_ (.A(_11047_),
    .Z(_11149_));
 XNOR2_X2 _33685_ (.A(_11136_),
    .B(_08121_),
    .ZN(_11150_));
 XNOR2_X2 _33686_ (.A(_09321_),
    .B(_06863_),
    .ZN(_11151_));
 XNOR2_X1 _33687_ (.A(_11150_),
    .B(_11151_),
    .ZN(_11152_));
 XNOR2_X1 _33688_ (.A(_10624_),
    .B(_11152_),
    .ZN(_11153_));
 NAND2_X1 _33689_ (.A1(_08039_),
    .A2(_11153_),
    .ZN(_11154_));
 OAI21_X2 _33690_ (.A(_11154_),
    .B1(_07243_),
    .B2(_00424_),
    .ZN(_11155_));
 OAI22_X1 _33691_ (.A1(\block_reg[2][16] ),
    .A2(_09134_),
    .B1(_09222_),
    .B2(_11155_),
    .ZN(_11156_));
 NOR2_X1 _33692_ (.A1(_17905_),
    .A2(_11156_),
    .ZN(_11157_));
 AOI22_X2 _33693_ (.A1(\block_reg[2][16] ),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_11155_),
    .ZN(_11158_));
 AOI21_X2 _33694_ (.A(_11157_),
    .B1(_11158_),
    .B2(_17905_),
    .ZN(_11159_));
 NOR3_X1 _33695_ (.A1(_08598_),
    .A2(_11149_),
    .A3(_11159_),
    .ZN(_11160_));
 INV_X1 _33696_ (.A(_08178_),
    .ZN(_11161_));
 AOI21_X1 _33697_ (.A(_11160_),
    .B1(_11049_),
    .B2(_11161_),
    .ZN(_00773_));
 INV_X1 _33698_ (.A(_08185_),
    .ZN(_11162_));
 AND2_X1 _33699_ (.A1(_00427_),
    .A2(_10223_),
    .ZN(_11163_));
 XNOR2_X1 _33700_ (.A(_11136_),
    .B(_10682_),
    .ZN(_11164_));
 XNOR2_X1 _33701_ (.A(_06802_),
    .B(_11052_),
    .ZN(_11165_));
 XNOR2_X2 _33702_ (.A(_11164_),
    .B(_11165_),
    .ZN(_11166_));
 XNOR2_X2 _33703_ (.A(_10624_),
    .B(_08121_),
    .ZN(_11167_));
 XNOR2_X1 _33704_ (.A(_00309_),
    .B(_11167_),
    .ZN(_11168_));
 XNOR2_X2 _33705_ (.A(_11166_),
    .B(_11168_),
    .ZN(_11169_));
 AOI21_X4 _33706_ (.A(_11163_),
    .B1(_11169_),
    .B2(_07801_),
    .ZN(_11170_));
 OAI221_X2 _33707_ (.A(_18258_),
    .B1(_10700_),
    .B2(_11170_),
    .C1(_10707_),
    .C2(\block_reg[2][17] ),
    .ZN(_11171_));
 NAND2_X1 _33708_ (.A1(_09211_),
    .A2(_11170_),
    .ZN(_11172_));
 INV_X1 _33709_ (.A(\block_reg[2][17] ),
    .ZN(_11173_));
 OAI21_X1 _33710_ (.A(_11172_),
    .B1(_08888_),
    .B2(_11173_),
    .ZN(_11174_));
 OR2_X1 _33711_ (.A1(_18258_),
    .A2(_11174_),
    .ZN(_11175_));
 AOI21_X2 _33712_ (.A(_11048_),
    .B1(_11171_),
    .B2(_11175_),
    .ZN(_11176_));
 AOI22_X1 _33713_ (.A1(_11162_),
    .A2(_11076_),
    .B1(_11176_),
    .B2(_08716_),
    .ZN(_00774_));
 INV_X1 _33714_ (.A(_08199_),
    .ZN(_11177_));
 INV_X1 _33715_ (.A(\block_reg[2][18] ),
    .ZN(_11178_));
 CLKBUF_X3 _33716_ (.A(\core.enc_block.block_w3_reg[17] ),
    .Z(_11179_));
 XNOR2_X1 _33717_ (.A(_07258_),
    .B(_10682_),
    .ZN(_11180_));
 XNOR2_X2 _33718_ (.A(_11063_),
    .B(_11180_),
    .ZN(_11181_));
 XNOR2_X1 _33719_ (.A(_11179_),
    .B(_11181_),
    .ZN(_11182_));
 MUX2_X2 _33720_ (.A(_00430_),
    .B(_11182_),
    .S(_07232_),
    .Z(_11183_));
 OAI22_X1 _33721_ (.A1(_11178_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_11183_),
    .ZN(_11184_));
 NOR2_X1 _33722_ (.A1(_17562_),
    .A2(_11184_),
    .ZN(_11185_));
 AOI22_X2 _33723_ (.A1(_11178_),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_11183_),
    .ZN(_11186_));
 AOI21_X2 _33724_ (.A(_11185_),
    .B1(_11186_),
    .B2(_17562_),
    .ZN(_11187_));
 NOR2_X1 _33725_ (.A1(_11107_),
    .A2(_11187_),
    .ZN(_11188_));
 AOI22_X1 _33726_ (.A1(_11177_),
    .A2(_11076_),
    .B1(_11188_),
    .B2(_08804_),
    .ZN(_00775_));
 INV_X1 _33727_ (.A(_08207_),
    .ZN(_11189_));
 XNOR2_X1 _33728_ (.A(_11064_),
    .B(_07659_),
    .ZN(_11190_));
 XNOR2_X1 _33729_ (.A(_11150_),
    .B(_11190_),
    .ZN(_11191_));
 XNOR2_X1 _33730_ (.A(_11078_),
    .B(_11191_),
    .ZN(_11192_));
 NAND2_X1 _33731_ (.A1(_09217_),
    .A2(_11192_),
    .ZN(_11193_));
 OAI21_X2 _33732_ (.A(_11193_),
    .B1(_10172_),
    .B2(_00433_),
    .ZN(_11194_));
 OAI22_X1 _33733_ (.A1(\block_reg[2][19] ),
    .A2(_07905_),
    .B1(_08889_),
    .B2(_11194_),
    .ZN(_11195_));
 OR2_X1 _33734_ (.A1(_17810_),
    .A2(_11195_),
    .ZN(_11196_));
 AOI22_X1 _33735_ (.A1(\block_reg[2][19] ),
    .A2(_10695_),
    .B1(_10696_),
    .B2(_11194_),
    .ZN(_11197_));
 NAND2_X1 _33736_ (.A1(_17810_),
    .A2(_11197_),
    .ZN(_11198_));
 AOI21_X1 _33737_ (.A(_11048_),
    .B1(_11196_),
    .B2(_11198_),
    .ZN(_11199_));
 AOI22_X1 _33738_ (.A1(_11189_),
    .A2(_11076_),
    .B1(_11199_),
    .B2(_08887_),
    .ZN(_00776_));
 INV_X1 _33739_ (.A(_06800_),
    .ZN(_11200_));
 XNOR2_X1 _33740_ (.A(_06863_),
    .B(_11179_),
    .ZN(_11201_));
 XNOR2_X1 _33741_ (.A(_09310_),
    .B(_06740_),
    .ZN(_11202_));
 XNOR2_X1 _33742_ (.A(_11201_),
    .B(_11202_),
    .ZN(_11203_));
 XNOR2_X1 _33743_ (.A(_07298_),
    .B(_11051_),
    .ZN(_11204_));
 XOR2_X1 _33744_ (.A(_11203_),
    .B(_11204_),
    .Z(_11205_));
 MUX2_X2 _33745_ (.A(_06802_),
    .B(_11205_),
    .S(_07232_),
    .Z(_11206_));
 OAI22_X1 _33746_ (.A1(\block_reg[2][1] ),
    .A2(_10232_),
    .B1(_11017_),
    .B2(_11206_),
    .ZN(_11207_));
 NAND2_X1 _33747_ (.A1(_10891_),
    .A2(_11206_),
    .ZN(_11208_));
 OAI21_X1 _33748_ (.A(_11208_),
    .B1(_10992_),
    .B2(_05900_),
    .ZN(_11209_));
 MUX2_X1 _33749_ (.A(_11207_),
    .B(_11209_),
    .S(_17671_),
    .Z(_11210_));
 NOR2_X1 _33750_ (.A1(_11107_),
    .A2(_11210_),
    .ZN(_11211_));
 AOI22_X1 _33751_ (.A1(_11200_),
    .A2(_11076_),
    .B1(_11211_),
    .B2(_08997_),
    .ZN(_00777_));
 XOR2_X1 _33752_ (.A(_11136_),
    .B(_07813_),
    .Z(_11212_));
 XNOR2_X1 _33753_ (.A(_06770_),
    .B(_11080_),
    .ZN(_11213_));
 XNOR2_X1 _33754_ (.A(_11212_),
    .B(_11213_),
    .ZN(_11214_));
 XNOR2_X1 _33755_ (.A(_00310_),
    .B(_11096_),
    .ZN(_11215_));
 XNOR2_X1 _33756_ (.A(_11214_),
    .B(_11215_),
    .ZN(_11216_));
 NOR2_X1 _33757_ (.A1(_10223_),
    .A2(_11216_),
    .ZN(_11217_));
 AOI21_X2 _33758_ (.A(_11217_),
    .B1(_07902_),
    .B2(_00413_),
    .ZN(_11218_));
 AOI22_X1 _33759_ (.A1(\block_reg[2][20] ),
    .A2(_09005_),
    .B1(_07908_),
    .B2(_11218_),
    .ZN(_11219_));
 NAND2_X1 _33760_ (.A1(_18296_),
    .A2(_11219_),
    .ZN(_11220_));
 OAI22_X1 _33761_ (.A1(\block_reg[2][20] ),
    .A2(_09221_),
    .B1(_09223_),
    .B2(_11218_),
    .ZN(_11221_));
 OAI21_X1 _33762_ (.A(_11220_),
    .B1(_11221_),
    .B2(_18296_),
    .ZN(_11222_));
 NAND2_X1 _33763_ (.A1(_09059_),
    .A2(_11222_),
    .ZN(_11223_));
 MUX2_X1 _33764_ (.A(_11223_),
    .B(_08218_),
    .S(_11107_),
    .Z(_00778_));
 INV_X1 _33765_ (.A(_08225_),
    .ZN(_11224_));
 INV_X1 _33766_ (.A(\core.enc_block.block_w3_reg[20] ),
    .ZN(_11225_));
 XNOR2_X1 _33767_ (.A(_07913_),
    .B(_07813_),
    .ZN(_11226_));
 XNOR2_X1 _33768_ (.A(_11108_),
    .B(_11226_),
    .ZN(_11227_));
 XNOR2_X1 _33769_ (.A(_11225_),
    .B(_11227_),
    .ZN(_11228_));
 NOR2_X1 _33770_ (.A1(_07902_),
    .A2(_11228_),
    .ZN(_11229_));
 AOI21_X2 _33771_ (.A(_11229_),
    .B1(_07902_),
    .B2(_00416_),
    .ZN(_11230_));
 OAI221_X1 _33772_ (.A(_17890_),
    .B1(_10700_),
    .B2(_11230_),
    .C1(_10707_),
    .C2(\block_reg[2][21] ),
    .ZN(_11231_));
 MUX2_X2 _33773_ (.A(_00257_),
    .B(_17889_),
    .S(_16489_),
    .Z(_11232_));
 AOI22_X1 _33774_ (.A1(\block_reg[2][21] ),
    .A2(_10695_),
    .B1(_10696_),
    .B2(_11230_),
    .ZN(_11233_));
 NAND2_X1 _33775_ (.A1(_11232_),
    .A2(_11233_),
    .ZN(_11234_));
 AOI21_X1 _33776_ (.A(_11048_),
    .B1(_11231_),
    .B2(_11234_),
    .ZN(_11235_));
 AOI22_X1 _33777_ (.A1(_11224_),
    .A2(_11076_),
    .B1(_11235_),
    .B2(_09124_),
    .ZN(_00779_));
 XNOR2_X2 _33778_ (.A(_11109_),
    .B(_07913_),
    .ZN(_11236_));
 XNOR2_X1 _33779_ (.A(_11122_),
    .B(_11236_),
    .ZN(_11237_));
 XNOR2_X1 _33780_ (.A(_08056_),
    .B(_11237_),
    .ZN(_11238_));
 NAND2_X1 _33781_ (.A1(_08809_),
    .A2(_11238_),
    .ZN(_11239_));
 OAI21_X2 _33782_ (.A(_11239_),
    .B1(_10265_),
    .B2(_00419_),
    .ZN(_11240_));
 AOI22_X1 _33783_ (.A1(\block_reg[2][22] ),
    .A2(_10905_),
    .B1(_10956_),
    .B2(_11240_),
    .ZN(_11241_));
 INV_X1 _33784_ (.A(_11241_),
    .ZN(_11242_));
 OAI22_X1 _33785_ (.A1(\block_reg[2][22] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_11240_),
    .ZN(_11243_));
 MUX2_X1 _33786_ (.A(_11242_),
    .B(_11243_),
    .S(_17573_),
    .Z(_11244_));
 NOR3_X1 _33787_ (.A1(_09172_),
    .A2(_11149_),
    .A3(_11244_),
    .ZN(_11245_));
 AOI21_X1 _33788_ (.A(_11245_),
    .B1(_11049_),
    .B2(_10957_),
    .ZN(_00780_));
 XNOR2_X2 _33789_ (.A(_11123_),
    .B(_08056_),
    .ZN(_11246_));
 XNOR2_X1 _33790_ (.A(_11079_),
    .B(_11246_),
    .ZN(_11247_));
 XNOR2_X1 _33791_ (.A(_09255_),
    .B(_11247_),
    .ZN(_11248_));
 NAND2_X1 _33792_ (.A1(_10717_),
    .A2(_11248_),
    .ZN(_11249_));
 OAI21_X2 _33793_ (.A(_11249_),
    .B1(_10948_),
    .B2(_00422_),
    .ZN(_11250_));
 OAI22_X1 _33794_ (.A1(\block_reg[2][23] ),
    .A2(_10232_),
    .B1(_11017_),
    .B2(_11250_),
    .ZN(_11251_));
 NAND2_X1 _33795_ (.A1(_10891_),
    .A2(_11250_),
    .ZN(_11252_));
 OAI21_X1 _33796_ (.A(_11252_),
    .B1(_10992_),
    .B2(_06542_),
    .ZN(_11253_));
 MUX2_X1 _33797_ (.A(_11251_),
    .B(_11253_),
    .S(_17551_),
    .Z(_11254_));
 NOR2_X1 _33798_ (.A1(_11107_),
    .A2(_11254_),
    .ZN(_11255_));
 AOI22_X1 _33799_ (.A1(_10966_),
    .A2(_11062_),
    .B1(_11255_),
    .B2(_09210_),
    .ZN(_00781_));
 XOR2_X1 _33800_ (.A(_11053_),
    .B(_11137_),
    .Z(_11256_));
 XNOR2_X1 _33801_ (.A(_06863_),
    .B(_11256_),
    .ZN(_11257_));
 MUX2_X1 _33802_ (.A(_09321_),
    .B(_11257_),
    .S(_08038_),
    .Z(_11258_));
 AOI22_X1 _33803_ (.A1(\block_reg[2][24] ),
    .A2(_09125_),
    .B1(_07229_),
    .B2(_11258_),
    .ZN(_11259_));
 OAI22_X1 _33804_ (.A1(\block_reg[2][24] ),
    .A2(_07904_),
    .B1(_09007_),
    .B2(_11258_),
    .ZN(_11260_));
 INV_X1 _33805_ (.A(_11260_),
    .ZN(_11261_));
 MUX2_X1 _33806_ (.A(_11259_),
    .B(_11261_),
    .S(_17642_),
    .Z(_11262_));
 NAND2_X1 _33807_ (.A1(_09682_),
    .A2(_11262_),
    .ZN(_11263_));
 MUX2_X1 _33808_ (.A(_11263_),
    .B(_09321_),
    .S(_11149_),
    .Z(_00782_));
 INV_X1 _33809_ (.A(_09310_),
    .ZN(_11264_));
 AND2_X1 _33810_ (.A1(_00309_),
    .A2(_10223_),
    .ZN(_11265_));
 XNOR2_X1 _33811_ (.A(_00427_),
    .B(_11051_),
    .ZN(_11266_));
 XNOR2_X1 _33812_ (.A(_11166_),
    .B(_11266_),
    .ZN(_11267_));
 AOI21_X2 _33813_ (.A(_11265_),
    .B1(_11267_),
    .B2(_07801_),
    .ZN(_11268_));
 OAI221_X1 _33814_ (.A(_17795_),
    .B1(_10700_),
    .B2(_11268_),
    .C1(_10707_),
    .C2(\block_reg[2][25] ),
    .ZN(_11269_));
 NAND2_X1 _33815_ (.A1(_09211_),
    .A2(_11268_),
    .ZN(_11270_));
 INV_X1 _33816_ (.A(\block_reg[2][25] ),
    .ZN(_11271_));
 OAI21_X1 _33817_ (.A(_11270_),
    .B1(_08888_),
    .B2(_11271_),
    .ZN(_11272_));
 OR2_X1 _33818_ (.A1(_17795_),
    .A2(_11272_),
    .ZN(_11273_));
 AOI21_X1 _33819_ (.A(_11048_),
    .B1(_11269_),
    .B2(_11273_),
    .ZN(_11274_));
 AOI22_X1 _33820_ (.A1(_11264_),
    .A2(_11062_),
    .B1(_11274_),
    .B2(_09778_),
    .ZN(_00783_));
 XNOR2_X1 _33821_ (.A(_11064_),
    .B(_07258_),
    .ZN(_11275_));
 XNOR2_X1 _33822_ (.A(_09310_),
    .B(_11275_),
    .ZN(_11276_));
 XNOR2_X1 _33823_ (.A(_06790_),
    .B(_11179_),
    .ZN(_11277_));
 XNOR2_X1 _33824_ (.A(_11276_),
    .B(_11277_),
    .ZN(_11278_));
 MUX2_X1 _33825_ (.A(_09243_),
    .B(_11278_),
    .S(_09131_),
    .Z(_11279_));
 AOI22_X1 _33826_ (.A1(\block_reg[2][26] ),
    .A2(_10905_),
    .B1(_10956_),
    .B2(_11279_),
    .ZN(_11280_));
 INV_X1 _33827_ (.A(_11280_),
    .ZN(_11281_));
 OAI22_X1 _33828_ (.A1(\block_reg[2][26] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_11279_),
    .ZN(_11282_));
 MUX2_X1 _33829_ (.A(_11281_),
    .B(_11282_),
    .S(_17591_),
    .Z(_11283_));
 NOR3_X1 _33830_ (.A1(_09860_),
    .A2(_11149_),
    .A3(_11283_),
    .ZN(_11284_));
 AOI21_X1 _33831_ (.A(_11284_),
    .B1(_11049_),
    .B2(_09244_),
    .ZN(_00784_));
 XOR2_X1 _33832_ (.A(_11137_),
    .B(_11190_),
    .Z(_11285_));
 XNOR2_X1 _33833_ (.A(_06721_),
    .B(_00433_),
    .ZN(_11286_));
 XNOR2_X1 _33834_ (.A(_09244_),
    .B(_11286_),
    .ZN(_11287_));
 XNOR2_X1 _33835_ (.A(_11285_),
    .B(_11287_),
    .ZN(_11288_));
 MUX2_X1 _33836_ (.A(_09231_),
    .B(_11288_),
    .S(_07651_),
    .Z(_11289_));
 OAI22_X1 _33837_ (.A1(\block_reg[2][27] ),
    .A2(_09134_),
    .B1(_09222_),
    .B2(_11289_),
    .ZN(_11290_));
 NOR2_X1 _33838_ (.A1(_17921_),
    .A2(_11290_),
    .ZN(_11291_));
 AOI22_X1 _33839_ (.A1(\block_reg[2][27] ),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_11289_),
    .ZN(_11292_));
 AOI21_X2 _33840_ (.A(_11291_),
    .B1(_11292_),
    .B2(_17921_),
    .ZN(_11293_));
 NOR3_X1 _33841_ (.A1(_09950_),
    .A2(_11149_),
    .A3(_11293_),
    .ZN(_11294_));
 INV_X1 _33842_ (.A(_09231_),
    .ZN(_11295_));
 AOI21_X1 _33843_ (.A(_11294_),
    .B1(_11049_),
    .B2(_11295_),
    .ZN(_00785_));
 XNOR2_X2 _33844_ (.A(_09255_),
    .B(_09231_),
    .ZN(_11296_));
 XNOR2_X1 _33845_ (.A(_00413_),
    .B(_11296_),
    .ZN(_11297_));
 XNOR2_X1 _33846_ (.A(_11214_),
    .B(_11297_),
    .ZN(_11298_));
 NOR2_X1 _33847_ (.A1(_10223_),
    .A2(_11298_),
    .ZN(_11299_));
 AOI21_X2 _33848_ (.A(_11299_),
    .B1(_10223_),
    .B2(_00310_),
    .ZN(_11300_));
 AOI22_X1 _33849_ (.A1(\block_reg[2][28] ),
    .A2(_10905_),
    .B1(_10956_),
    .B2(_11300_),
    .ZN(_11301_));
 INV_X1 _33850_ (.A(_11301_),
    .ZN(_11302_));
 OAI22_X1 _33851_ (.A1(\block_reg[2][28] ),
    .A2(_10678_),
    .B1(_10269_),
    .B2(_11300_),
    .ZN(_11303_));
 MUX2_X1 _33852_ (.A(_11302_),
    .B(_11303_),
    .S(_18309_),
    .Z(_11304_));
 NOR3_X1 _33853_ (.A1(_10010_),
    .A2(_11149_),
    .A3(_11304_),
    .ZN(_11305_));
 INV_X1 _33854_ (.A(\core.enc_block.block_w2_reg[28] ),
    .ZN(_11306_));
 AOI21_X1 _33855_ (.A(_11305_),
    .B1(_11049_),
    .B2(_11306_),
    .ZN(_00786_));
 XNOR2_X1 _33856_ (.A(_11093_),
    .B(_11236_),
    .ZN(_11307_));
 XNOR2_X1 _33857_ (.A(_06763_),
    .B(_11307_),
    .ZN(_11308_));
 MUX2_X1 _33858_ (.A(_09275_),
    .B(_11308_),
    .S(_08038_),
    .Z(_11309_));
 AOI22_X1 _33859_ (.A1(\block_reg[2][29] ),
    .A2(_09125_),
    .B1(_07229_),
    .B2(_11309_),
    .ZN(_11310_));
 OAI22_X1 _33860_ (.A1(\block_reg[2][29] ),
    .A2(_07904_),
    .B1(_09007_),
    .B2(_11309_),
    .ZN(_11311_));
 INV_X1 _33861_ (.A(_11311_),
    .ZN(_11312_));
 MUX2_X1 _33862_ (.A(_11310_),
    .B(_11312_),
    .S(_17945_),
    .Z(_11313_));
 NAND2_X1 _33863_ (.A1(_10076_),
    .A2(_11313_),
    .ZN(_11314_));
 MUX2_X1 _33864_ (.A(_11314_),
    .B(_09275_),
    .S(_11149_),
    .Z(_00787_));
 INV_X1 _33865_ (.A(_06788_),
    .ZN(_11315_));
 XNOR2_X1 _33866_ (.A(_09243_),
    .B(_06802_),
    .ZN(_11316_));
 XNOR2_X1 _33867_ (.A(_11276_),
    .B(_11316_),
    .ZN(_11317_));
 MUX2_X2 _33868_ (.A(_06790_),
    .B(_11317_),
    .S(_08039_),
    .Z(_11318_));
 OAI22_X1 _33869_ (.A1(\block_reg[2][2] ),
    .A2(_07905_),
    .B1(_08889_),
    .B2(_11318_),
    .ZN(_11319_));
 OR2_X1 _33870_ (.A1(_17534_),
    .A2(_11319_),
    .ZN(_11320_));
 AOI22_X1 _33871_ (.A1(\block_reg[2][2] ),
    .A2(_10695_),
    .B1(_10696_),
    .B2(_11318_),
    .ZN(_11321_));
 NAND2_X1 _33872_ (.A1(_17534_),
    .A2(_11321_),
    .ZN(_11322_));
 AOI21_X1 _33873_ (.A(_11047_),
    .B1(_11320_),
    .B2(_11322_),
    .ZN(_11323_));
 AOI22_X1 _33874_ (.A1(_11315_),
    .A2(_11062_),
    .B1(_11323_),
    .B2(_10168_),
    .ZN(_00788_));
 XNOR2_X1 _33875_ (.A(_06751_),
    .B(_11109_),
    .ZN(_11324_));
 XNOR2_X1 _33876_ (.A(_11246_),
    .B(_11324_),
    .ZN(_11325_));
 XNOR2_X1 _33877_ (.A(_09275_),
    .B(_11325_),
    .ZN(_11326_));
 MUX2_X1 _33878_ (.A(_09262_),
    .B(_11326_),
    .S(_09131_),
    .Z(_11327_));
 AOI22_X1 _33879_ (.A1(\block_reg[2][30] ),
    .A2(_10905_),
    .B1(_10956_),
    .B2(_11327_),
    .ZN(_11328_));
 INV_X1 _33880_ (.A(_11328_),
    .ZN(_11329_));
 OAI22_X1 _33881_ (.A1(\block_reg[2][30] ),
    .A2(_10678_),
    .B1(_08105_),
    .B2(_11327_),
    .ZN(_11330_));
 MUX2_X1 _33882_ (.A(_11329_),
    .B(_11330_),
    .S(_17603_),
    .Z(_11331_));
 NOR3_X1 _33883_ (.A1(_10222_),
    .A2(_11149_),
    .A3(_11331_),
    .ZN(_11332_));
 AOI21_X1 _33884_ (.A(_11332_),
    .B1(_11049_),
    .B2(_09263_),
    .ZN(_00789_));
 XOR2_X1 _33885_ (.A(_00308_),
    .B(_11123_),
    .Z(_11333_));
 XNOR2_X1 _33886_ (.A(_11150_),
    .B(_11333_),
    .ZN(_11334_));
 XNOR2_X1 _33887_ (.A(_09262_),
    .B(_11334_),
    .ZN(_11335_));
 MUX2_X1 _33888_ (.A(_09255_),
    .B(_11335_),
    .S(_07651_),
    .Z(_11336_));
 OAI22_X1 _33889_ (.A1(\block_reg[2][31] ),
    .A2(_09134_),
    .B1(_09222_),
    .B2(_11336_),
    .ZN(_11337_));
 NOR2_X1 _33890_ (.A1(_17934_),
    .A2(_11337_),
    .ZN(_11338_));
 AOI22_X1 _33891_ (.A1(\block_reg[2][31] ),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_11336_),
    .ZN(_11339_));
 AOI21_X1 _33892_ (.A(_11338_),
    .B1(_11339_),
    .B2(_17934_),
    .ZN(_11340_));
 NOR3_X2 _33893_ (.A1(_10261_),
    .A2(_11048_),
    .A3(_11340_),
    .ZN(_11341_));
 AOI21_X1 _33894_ (.A(_11341_),
    .B1(_11049_),
    .B2(_09256_),
    .ZN(_00790_));
 XNOR2_X1 _33895_ (.A(_11063_),
    .B(_11296_),
    .ZN(_11342_));
 XNOR2_X1 _33896_ (.A(_00402_),
    .B(_11080_),
    .ZN(_11343_));
 XNOR2_X1 _33897_ (.A(_06741_),
    .B(_11343_),
    .ZN(_11344_));
 XNOR2_X1 _33898_ (.A(_11342_),
    .B(_11344_),
    .ZN(_11345_));
 MUX2_X1 _33899_ (.A(_06722_),
    .B(_11345_),
    .S(_07242_),
    .Z(_11346_));
 AOI221_X1 _33900_ (.A(_17861_),
    .B1(_07808_),
    .B2(_11346_),
    .C1(_09005_),
    .C2(_06058_),
    .ZN(_11347_));
 NOR2_X1 _33901_ (.A1(_09007_),
    .A2(_11346_),
    .ZN(_11348_));
 AOI21_X1 _33902_ (.A(_11348_),
    .B1(_08900_),
    .B2(\block_reg[2][3] ),
    .ZN(_11349_));
 AND2_X1 _33903_ (.A1(_17861_),
    .A2(_11349_),
    .ZN(_11350_));
 OAI21_X1 _33904_ (.A(_10353_),
    .B1(_11347_),
    .B2(_11350_),
    .ZN(_11351_));
 MUX2_X1 _33905_ (.A(_11351_),
    .B(_06714_),
    .S(_11149_),
    .Z(_00791_));
 INV_X1 _33906_ (.A(_06768_),
    .ZN(_11352_));
 XNOR2_X1 _33907_ (.A(_07323_),
    .B(_11296_),
    .ZN(_11353_));
 XNOR2_X1 _33908_ (.A(_11095_),
    .B(_11353_),
    .ZN(_11354_));
 MUX2_X2 _33909_ (.A(_06770_),
    .B(_11354_),
    .S(_07232_),
    .Z(_11355_));
 OAI22_X1 _33910_ (.A1(\block_reg[2][4] ),
    .A2(_10232_),
    .B1(_11017_),
    .B2(_11355_),
    .ZN(_11356_));
 NAND2_X1 _33911_ (.A1(_10716_),
    .A2(_11355_),
    .ZN(_11357_));
 INV_X1 _33912_ (.A(\block_reg[2][4] ),
    .ZN(_11358_));
 OAI21_X1 _33913_ (.A(_11357_),
    .B1(_10992_),
    .B2(_11358_),
    .ZN(_11359_));
 MUX2_X1 _33914_ (.A(_11356_),
    .B(_11359_),
    .S(_18281_),
    .Z(_11360_));
 NOR2_X1 _33915_ (.A1(_11107_),
    .A2(_11360_),
    .ZN(_11361_));
 AOI22_X1 _33916_ (.A1(_11352_),
    .A2(_11062_),
    .B1(_11361_),
    .B2(_10414_),
    .ZN(_00792_));
 INV_X1 _33917_ (.A(_06761_),
    .ZN(_11362_));
 XOR2_X1 _33918_ (.A(_09275_),
    .B(_06770_),
    .Z(_11363_));
 XNOR2_X1 _33919_ (.A(_11236_),
    .B(_11363_),
    .ZN(_11364_));
 XNOR2_X1 _33920_ (.A(_11306_),
    .B(_11364_),
    .ZN(_11365_));
 MUX2_X2 _33921_ (.A(_06763_),
    .B(_11365_),
    .S(_07232_),
    .Z(_11366_));
 NAND2_X1 _33922_ (.A1(_09126_),
    .A2(_11366_),
    .ZN(_11367_));
 INV_X1 _33923_ (.A(\block_reg[2][5] ),
    .ZN(_11368_));
 OAI21_X1 _33924_ (.A(_11367_),
    .B1(_07248_),
    .B2(_11368_),
    .ZN(_11369_));
 OAI22_X1 _33925_ (.A1(\block_reg[2][5] ),
    .A2(_10476_),
    .B1(_10795_),
    .B2(_11366_),
    .ZN(_11370_));
 MUX2_X1 _33926_ (.A(_11369_),
    .B(_11370_),
    .S(_17760_),
    .Z(_11371_));
 NOR2_X1 _33927_ (.A1(_11107_),
    .A2(_11371_),
    .ZN(_11372_));
 AOI22_X1 _33928_ (.A1(_11362_),
    .A2(_11062_),
    .B1(_11372_),
    .B2(_10470_),
    .ZN(_00793_));
 XOR2_X1 _33929_ (.A(_11108_),
    .B(_11246_),
    .Z(_11373_));
 XNOR2_X1 _33930_ (.A(_09262_),
    .B(_11373_),
    .ZN(_11374_));
 MUX2_X1 _33931_ (.A(_06751_),
    .B(_11374_),
    .S(_08038_),
    .Z(_11375_));
 AOI22_X1 _33932_ (.A1(\block_reg[2][6] ),
    .A2(_09125_),
    .B1(_07229_),
    .B2(_11375_),
    .ZN(_11376_));
 OAI22_X1 _33933_ (.A1(\block_reg[2][6] ),
    .A2(_07904_),
    .B1(_09007_),
    .B2(_11375_),
    .ZN(_11377_));
 INV_X1 _33934_ (.A(_11377_),
    .ZN(_11378_));
 MUX2_X1 _33935_ (.A(_11376_),
    .B(_11378_),
    .S(_17657_),
    .Z(_11379_));
 NAND2_X1 _33936_ (.A1(_10527_),
    .A2(_11379_),
    .ZN(_11380_));
 MUX2_X1 _33937_ (.A(_11380_),
    .B(_06748_),
    .S(_11149_),
    .Z(_00794_));
 INV_X1 _33938_ (.A(_06737_),
    .ZN(_11381_));
 XNOR2_X1 _33939_ (.A(_11122_),
    .B(_11150_),
    .ZN(_11382_));
 XNOR2_X1 _33940_ (.A(_09255_),
    .B(_11382_),
    .ZN(_11383_));
 NAND2_X1 _33941_ (.A1(_10717_),
    .A2(_11383_),
    .ZN(_11384_));
 OAI21_X2 _33942_ (.A(_11384_),
    .B1(_10948_),
    .B2(_00308_),
    .ZN(_11385_));
 OAI22_X1 _33943_ (.A1(\block_reg[2][7] ),
    .A2(_10232_),
    .B1(_11017_),
    .B2(_11385_),
    .ZN(_11386_));
 NAND2_X1 _33944_ (.A1(_10716_),
    .A2(_11385_),
    .ZN(_11387_));
 OAI21_X1 _33945_ (.A(_11387_),
    .B1(_10992_),
    .B2(_06105_),
    .ZN(_11388_));
 MUX2_X1 _33946_ (.A(_11386_),
    .B(_11388_),
    .S(_17517_),
    .Z(_11389_));
 NOR2_X1 _33947_ (.A1(_11107_),
    .A2(_11389_),
    .ZN(_11390_));
 AOI22_X1 _33948_ (.A1(_11381_),
    .A2(_11062_),
    .B1(_11390_),
    .B2(_10566_),
    .ZN(_00795_));
 INV_X1 _33949_ (.A(_07237_),
    .ZN(_11391_));
 XNOR2_X1 _33950_ (.A(_11079_),
    .B(_11151_),
    .ZN(_11392_));
 XNOR2_X1 _33951_ (.A(_11052_),
    .B(_11392_),
    .ZN(_11393_));
 NAND2_X1 _33952_ (.A1(_10717_),
    .A2(_11393_),
    .ZN(_11394_));
 OAI21_X2 _33953_ (.A(_11394_),
    .B1(_10948_),
    .B2(_00393_),
    .ZN(_11395_));
 OAI22_X1 _33954_ (.A1(\block_reg[2][8] ),
    .A2(_10232_),
    .B1(_11017_),
    .B2(_11395_),
    .ZN(_11396_));
 NAND2_X1 _33955_ (.A1(_10716_),
    .A2(_11395_),
    .ZN(_11397_));
 OAI21_X1 _33956_ (.A(_11397_),
    .B1(_10992_),
    .B2(_05716_),
    .ZN(_11398_));
 MUX2_X1 _33957_ (.A(_11396_),
    .B(_11398_),
    .S(_17617_),
    .Z(_11399_));
 NOR2_X1 _33958_ (.A1(_11107_),
    .A2(_11399_),
    .ZN(_11400_));
 AOI22_X1 _33959_ (.A1(_11391_),
    .A2(_11062_),
    .B1(_11400_),
    .B2(_10614_),
    .ZN(_00796_));
 XNOR2_X1 _33960_ (.A(_06802_),
    .B(_11167_),
    .ZN(_11401_));
 XNOR2_X1 _33961_ (.A(_11203_),
    .B(_11401_),
    .ZN(_11402_));
 NAND2_X1 _33962_ (.A1(_08809_),
    .A2(_11402_),
    .ZN(_11403_));
 OAI21_X2 _33963_ (.A(_11403_),
    .B1(_10265_),
    .B2(_07298_),
    .ZN(_11404_));
 AOI22_X1 _33964_ (.A1(\block_reg[2][9] ),
    .A2(_10905_),
    .B1(_10956_),
    .B2(_11404_),
    .ZN(_11405_));
 INV_X1 _33965_ (.A(_11405_),
    .ZN(_11406_));
 OAI22_X1 _33966_ (.A1(\block_reg[2][9] ),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_11404_),
    .ZN(_11407_));
 MUX2_X1 _33967_ (.A(_11406_),
    .B(_11407_),
    .S(_17688_),
    .Z(_11408_));
 NOR3_X1 _33968_ (.A1(_10670_),
    .A2(_11048_),
    .A3(_11408_),
    .ZN(_11409_));
 INV_X1 _33969_ (.A(_07292_),
    .ZN(_11410_));
 AOI21_X1 _33970_ (.A(_11409_),
    .B1(_11049_),
    .B2(_11410_),
    .ZN(_00797_));
 INV_X1 _33971_ (.A(\core.enc_block.block_w3_reg[0] ),
    .ZN(_11411_));
 AOI21_X4 _33972_ (.A(_06692_),
    .B1(_07260_),
    .B2(_16242_),
    .ZN(_11412_));
 BUF_X4 _33973_ (.A(_11412_),
    .Z(_11413_));
 BUF_X4 _33974_ (.A(_11413_),
    .Z(_11414_));
 CLKBUF_X3 _33975_ (.A(_11412_),
    .Z(_11415_));
 NOR2_X1 _33976_ (.A1(_06861_),
    .A2(_08896_),
    .ZN(_11416_));
 CLKBUF_X3 _33977_ (.A(\core.enc_block.block_w3_reg[31] ),
    .Z(_11417_));
 BUF_X2 _33978_ (.A(\core.enc_block.block_w3_reg[24] ),
    .Z(_11418_));
 XNOR2_X2 _33979_ (.A(_11417_),
    .B(_11418_),
    .ZN(_11419_));
 XNOR2_X2 _33980_ (.A(_07267_),
    .B(_08612_),
    .ZN(_11420_));
 XNOR2_X1 _33981_ (.A(_11419_),
    .B(_11420_),
    .ZN(_11421_));
 XNOR2_X1 _33982_ (.A(_00302_),
    .B(_11421_),
    .ZN(_11422_));
 AOI21_X2 _33983_ (.A(_11416_),
    .B1(_11422_),
    .B2(_08048_),
    .ZN(_11423_));
 NAND2_X1 _33984_ (.A1(_09126_),
    .A2(_11423_),
    .ZN(_11424_));
 INV_X1 _33985_ (.A(\block_reg[3][0] ),
    .ZN(_11425_));
 OAI21_X1 _33986_ (.A(_11424_),
    .B1(_07248_),
    .B2(_11425_),
    .ZN(_11426_));
 OAI22_X1 _33987_ (.A1(\block_reg[3][0] ),
    .A2(_10476_),
    .B1(_10795_),
    .B2(_11423_),
    .ZN(_11427_));
 MUX2_X1 _33988_ (.A(_11426_),
    .B(_11427_),
    .S(_19026_),
    .Z(_11428_));
 NOR2_X1 _33989_ (.A1(_11415_),
    .A2(_11428_),
    .ZN(_11429_));
 AOI22_X1 _33990_ (.A1(_11411_),
    .A2(_11414_),
    .B1(_11429_),
    .B2(_07223_),
    .ZN(_00798_));
 XOR2_X2 _33991_ (.A(\core.enc_block.block_w3_reg[26] ),
    .B(_06788_),
    .Z(_11430_));
 XNOR2_X1 _33992_ (.A(_08729_),
    .B(_00305_),
    .ZN(_11431_));
 XNOR2_X1 _33993_ (.A(_11430_),
    .B(_11431_),
    .ZN(_11432_));
 XNOR2_X1 _33994_ (.A(_06800_),
    .B(_11432_),
    .ZN(_11433_));
 MUX2_X1 _33995_ (.A(_07276_),
    .B(_11433_),
    .S(_08896_),
    .Z(_11434_));
 AOI22_X1 _33996_ (.A1(\block_reg[3][10] ),
    .A2(_09005_),
    .B1(_07908_),
    .B2(_11434_),
    .ZN(_11435_));
 NAND2_X1 _33997_ (.A1(_19411_),
    .A2(_11435_),
    .ZN(_11436_));
 OAI22_X1 _33998_ (.A1(\block_reg[3][10] ),
    .A2(_09221_),
    .B1(_09223_),
    .B2(_11434_),
    .ZN(_11437_));
 OAI21_X2 _33999_ (.A(_11436_),
    .B1(_11437_),
    .B2(_19411_),
    .ZN(_11438_));
 NAND2_X1 _34000_ (.A1(_07642_),
    .A2(_11438_),
    .ZN(_11439_));
 BUF_X4 _34001_ (.A(_11412_),
    .Z(_11440_));
 MUX2_X1 _34002_ (.A(_11439_),
    .B(_10721_),
    .S(_11440_),
    .Z(_00799_));
 INV_X1 _34003_ (.A(_10739_),
    .ZN(_11441_));
 XNOR2_X2 _34004_ (.A(_06737_),
    .B(_07340_),
    .ZN(_11442_));
 BUF_X2 _34005_ (.A(\core.enc_block.block_w3_reg[27] ),
    .Z(_11443_));
 XNOR2_X2 _34006_ (.A(_11443_),
    .B(_08905_),
    .ZN(_11444_));
 XNOR2_X1 _34007_ (.A(_11442_),
    .B(_11444_),
    .ZN(_11445_));
 XNOR2_X1 _34008_ (.A(_06714_),
    .B(_07276_),
    .ZN(_11446_));
 XNOR2_X1 _34009_ (.A(_06788_),
    .B(_11446_),
    .ZN(_11447_));
 XNOR2_X1 _34010_ (.A(_11445_),
    .B(_11447_),
    .ZN(_11448_));
 NAND2_X1 _34011_ (.A1(_10354_),
    .A2(_11448_),
    .ZN(_11449_));
 OAI21_X2 _34012_ (.A(_11449_),
    .B1(_07801_),
    .B2(_00303_),
    .ZN(_11450_));
 OAI221_X2 _34013_ (.A(_03343_),
    .B1(_10700_),
    .B2(_11450_),
    .C1(_10707_),
    .C2(\block_reg[3][11] ),
    .ZN(_11451_));
 NAND2_X1 _34014_ (.A1(_09211_),
    .A2(_11450_),
    .ZN(_11452_));
 INV_X1 _34015_ (.A(\block_reg[3][11] ),
    .ZN(_11453_));
 OAI21_X1 _34016_ (.A(_11452_),
    .B1(_08888_),
    .B2(_11453_),
    .ZN(_11454_));
 OR2_X1 _34017_ (.A1(_03343_),
    .A2(_11454_),
    .ZN(_11455_));
 AOI21_X2 _34018_ (.A(_11413_),
    .B1(_11451_),
    .B2(_11455_),
    .ZN(_11456_));
 AOI22_X1 _34019_ (.A1(_11441_),
    .A2(_11414_),
    .B1(_11456_),
    .B2(_07786_),
    .ZN(_00800_));
 BUF_X1 _34020_ (.A(\core.enc_block.block_w3_reg[28] ),
    .Z(_11457_));
 XNOR2_X1 _34021_ (.A(_11457_),
    .B(_09012_),
    .ZN(_11458_));
 XNOR2_X1 _34022_ (.A(_06737_),
    .B(_06714_),
    .ZN(_11459_));
 XNOR2_X1 _34023_ (.A(_11458_),
    .B(_11459_),
    .ZN(_11460_));
 XNOR2_X2 _34024_ (.A(_07340_),
    .B(_07285_),
    .ZN(_11461_));
 XNOR2_X1 _34025_ (.A(_06768_),
    .B(_11461_),
    .ZN(_11462_));
 XNOR2_X1 _34026_ (.A(_11460_),
    .B(_11462_),
    .ZN(_11463_));
 NAND2_X1 _34027_ (.A1(_10354_),
    .A2(_11463_),
    .ZN(_11464_));
 OAI21_X2 _34028_ (.A(_11464_),
    .B1(_07801_),
    .B2(_00304_),
    .ZN(_11465_));
 AOI22_X1 _34029_ (.A1(\block_reg[3][12] ),
    .A2(_09005_),
    .B1(_07908_),
    .B2(_11465_),
    .ZN(_11466_));
 NAND2_X1 _34030_ (.A1(_03774_),
    .A2(_11466_),
    .ZN(_11467_));
 OAI22_X1 _34031_ (.A1(\block_reg[3][12] ),
    .A2(_09221_),
    .B1(_09223_),
    .B2(_11465_),
    .ZN(_11468_));
 OAI21_X2 _34032_ (.A(_11467_),
    .B1(_11468_),
    .B2(_03774_),
    .ZN(_11469_));
 NAND2_X1 _34033_ (.A1(_07892_),
    .A2(_11469_),
    .ZN(_11470_));
 MUX2_X1 _34034_ (.A(_11470_),
    .B(_10841_),
    .S(_11440_),
    .Z(_00801_));
 INV_X1 _34035_ (.A(_10854_),
    .ZN(_11471_));
 BUF_X4 _34036_ (.A(_11413_),
    .Z(_11472_));
 BUF_X2 _34037_ (.A(\core.enc_block.block_w3_reg[29] ),
    .Z(_11473_));
 XOR2_X2 _34038_ (.A(_06761_),
    .B(_11473_),
    .Z(_11474_));
 XNOR2_X1 _34039_ (.A(_00304_),
    .B(_09139_),
    .ZN(_11475_));
 XNOR2_X1 _34040_ (.A(_11474_),
    .B(_11475_),
    .ZN(_11476_));
 XNOR2_X1 _34041_ (.A(_06768_),
    .B(_11476_),
    .ZN(_11477_));
 NAND2_X1 _34042_ (.A1(_09217_),
    .A2(_11477_),
    .ZN(_11478_));
 OAI21_X1 _34043_ (.A(_11478_),
    .B1(_10172_),
    .B2(_00306_),
    .ZN(_11479_));
 OAI22_X1 _34044_ (.A1(\block_reg[3][13] ),
    .A2(_07905_),
    .B1(_08889_),
    .B2(_11479_),
    .ZN(_11480_));
 OR2_X1 _34045_ (.A1(_18969_),
    .A2(_11480_),
    .ZN(_11481_));
 AOI22_X1 _34046_ (.A1(\block_reg[3][13] ),
    .A2(_10695_),
    .B1(_10696_),
    .B2(_11479_),
    .ZN(_11482_));
 NAND2_X1 _34047_ (.A1(_18969_),
    .A2(_11482_),
    .ZN(_11483_));
 AOI21_X1 _34048_ (.A(_11413_),
    .B1(_11481_),
    .B2(_11483_),
    .ZN(_11484_));
 AOI22_X1 _34049_ (.A1(_11471_),
    .A2(_11472_),
    .B1(_11484_),
    .B2(_08037_),
    .ZN(_00802_));
 INV_X1 _34050_ (.A(_10865_),
    .ZN(_11485_));
 BUF_X4 _34051_ (.A(_11412_),
    .Z(_11486_));
 BUF_X2 _34052_ (.A(\core.enc_block.block_w3_reg[30] ),
    .Z(_11487_));
 XNOR2_X2 _34053_ (.A(_06748_),
    .B(_11487_),
    .ZN(_11488_));
 XOR2_X1 _34054_ (.A(_09183_),
    .B(_00306_),
    .Z(_11489_));
 XNOR2_X1 _34055_ (.A(_11488_),
    .B(_11489_),
    .ZN(_11490_));
 XNOR2_X1 _34056_ (.A(_06761_),
    .B(_11490_),
    .ZN(_11491_));
 NAND2_X1 _34057_ (.A1(_09217_),
    .A2(_11491_),
    .ZN(_11492_));
 OAI21_X1 _34058_ (.A(_11492_),
    .B1(_10172_),
    .B2(_00307_),
    .ZN(_11493_));
 OAI22_X1 _34059_ (.A1(\block_reg[3][14] ),
    .A2(_07905_),
    .B1(_08889_),
    .B2(_11493_),
    .ZN(_11494_));
 OR2_X1 _34060_ (.A1(_19223_),
    .A2(_11494_),
    .ZN(_11495_));
 AOI22_X1 _34061_ (.A1(\block_reg[3][14] ),
    .A2(_10695_),
    .B1(_10696_),
    .B2(_11493_),
    .ZN(_11496_));
 NAND2_X1 _34062_ (.A1(_19223_),
    .A2(_11496_),
    .ZN(_11497_));
 AOI21_X1 _34063_ (.A(_11486_),
    .B1(_11495_),
    .B2(_11497_),
    .ZN(_11498_));
 AOI22_X1 _34064_ (.A1(_11485_),
    .A2(_11472_),
    .B1(_11498_),
    .B2(_08102_),
    .ZN(_00803_));
 XNOR2_X2 _34065_ (.A(_11417_),
    .B(_09227_),
    .ZN(_11499_));
 XOR2_X1 _34066_ (.A(_06737_),
    .B(_00307_),
    .Z(_11500_));
 XNOR2_X1 _34067_ (.A(_11499_),
    .B(_11500_),
    .ZN(_11501_));
 XNOR2_X1 _34068_ (.A(_06748_),
    .B(_11501_),
    .ZN(_11502_));
 MUX2_X1 _34069_ (.A(_07340_),
    .B(_11502_),
    .S(_08896_),
    .Z(_11503_));
 AOI22_X1 _34070_ (.A1(\block_reg[3][15] ),
    .A2(_09005_),
    .B1(_07908_),
    .B2(_11503_),
    .ZN(_11504_));
 NAND2_X1 _34071_ (.A1(_18941_),
    .A2(_11504_),
    .ZN(_11505_));
 OAI22_X1 _34072_ (.A1(\block_reg[3][15] ),
    .A2(_09221_),
    .B1(_09223_),
    .B2(_11503_),
    .ZN(_11506_));
 OAI21_X1 _34073_ (.A(_11505_),
    .B1(_11506_),
    .B2(_18941_),
    .ZN(_11507_));
 NAND2_X1 _34074_ (.A1(_08164_),
    .A2(_11507_),
    .ZN(_11508_));
 MUX2_X1 _34075_ (.A(_11508_),
    .B(_10722_),
    .S(_11440_),
    .Z(_00804_));
 XNOR2_X2 _34076_ (.A(_07340_),
    .B(_07267_),
    .ZN(_11509_));
 XNOR2_X2 _34077_ (.A(_06861_),
    .B(_11418_),
    .ZN(_11510_));
 XNOR2_X1 _34078_ (.A(_11509_),
    .B(_11510_),
    .ZN(_11511_));
 XNOR2_X1 _34079_ (.A(_09227_),
    .B(_11511_),
    .ZN(_11512_));
 NAND2_X1 _34080_ (.A1(_08809_),
    .A2(_11512_),
    .ZN(_11513_));
 OAI21_X2 _34081_ (.A(_11513_),
    .B1(_10265_),
    .B2(_00423_),
    .ZN(_11514_));
 AOI22_X1 _34082_ (.A1(\block_reg[3][16] ),
    .A2(_10905_),
    .B1(_10956_),
    .B2(_11514_),
    .ZN(_11515_));
 INV_X1 _34083_ (.A(_11515_),
    .ZN(_11516_));
 OAI22_X1 _34084_ (.A1(\block_reg[3][16] ),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_11514_),
    .ZN(_11517_));
 MUX2_X1 _34085_ (.A(_11516_),
    .B(_11517_),
    .S(_18859_),
    .Z(_11518_));
 NOR3_X1 _34086_ (.A1(_08598_),
    .A2(_11440_),
    .A3(_11518_),
    .ZN(_11519_));
 INV_X1 _34087_ (.A(_11052_),
    .ZN(_11520_));
 AOI21_X1 _34088_ (.A(_11519_),
    .B1(_11414_),
    .B2(_11520_),
    .ZN(_00805_));
 INV_X1 _34089_ (.A(_11179_),
    .ZN(_11521_));
 AND2_X1 _34090_ (.A1(_00426_),
    .A2(_10223_),
    .ZN(_11522_));
 XNOR2_X1 _34091_ (.A(_08612_),
    .B(_09227_),
    .ZN(_11523_));
 XNOR2_X1 _34092_ (.A(_06800_),
    .B(_07294_),
    .ZN(_11524_));
 XNOR2_X2 _34093_ (.A(_11523_),
    .B(_11524_),
    .ZN(_11525_));
 XNOR2_X1 _34094_ (.A(_00344_),
    .B(_11509_),
    .ZN(_11526_));
 XNOR2_X1 _34095_ (.A(_11525_),
    .B(_11526_),
    .ZN(_11527_));
 AOI21_X2 _34096_ (.A(_11522_),
    .B1(_11527_),
    .B2(_10172_),
    .ZN(_11528_));
 OAI221_X2 _34097_ (.A(_19210_),
    .B1(_07893_),
    .B2(_11528_),
    .C1(_07906_),
    .C2(\block_reg[3][17] ),
    .ZN(_11529_));
 MUX2_X1 _34098_ (.A(_00267_),
    .B(_19209_),
    .S(_16489_),
    .Z(_11530_));
 AOI22_X1 _34099_ (.A1(\block_reg[3][17] ),
    .A2(_10695_),
    .B1(_07809_),
    .B2(_11528_),
    .ZN(_11531_));
 NAND2_X1 _34100_ (.A1(_11530_),
    .A2(_11531_),
    .ZN(_11532_));
 AOI21_X2 _34101_ (.A(_11486_),
    .B1(_11529_),
    .B2(_11532_),
    .ZN(_11533_));
 AOI22_X1 _34102_ (.A1(_11521_),
    .A2(_11472_),
    .B1(_11533_),
    .B2(_08716_),
    .ZN(_00806_));
 INV_X1 _34103_ (.A(_11064_),
    .ZN(_11534_));
 NOR2_X1 _34104_ (.A1(\block_reg[3][18] ),
    .A2(_10729_),
    .ZN(_11535_));
 XNOR2_X1 _34105_ (.A(_07276_),
    .B(_08614_),
    .ZN(_11536_));
 XNOR2_X1 _34106_ (.A(_11430_),
    .B(_11536_),
    .ZN(_11537_));
 XNOR2_X1 _34107_ (.A(_07294_),
    .B(_11537_),
    .ZN(_11538_));
 MUX2_X1 _34108_ (.A(_00429_),
    .B(_11538_),
    .S(_07243_),
    .Z(_11539_));
 AOI21_X1 _34109_ (.A(_11535_),
    .B1(_11539_),
    .B2(_10696_),
    .ZN(_11540_));
 NAND2_X1 _34110_ (.A1(_19396_),
    .A2(_11540_),
    .ZN(_11541_));
 NAND2_X1 _34111_ (.A1(\block_reg[3][18] ),
    .A2(_09005_),
    .ZN(_11542_));
 OAI21_X1 _34112_ (.A(_11542_),
    .B1(_11539_),
    .B2(_08889_),
    .ZN(_11543_));
 OR2_X1 _34113_ (.A1(_19396_),
    .A2(_11543_),
    .ZN(_11544_));
 AOI21_X2 _34114_ (.A(_11486_),
    .B1(_11541_),
    .B2(_11544_),
    .ZN(_11545_));
 AOI22_X1 _34115_ (.A1(_11534_),
    .A2(_11472_),
    .B1(_11545_),
    .B2(_08804_),
    .ZN(_00807_));
 INV_X1 _34116_ (.A(_11080_),
    .ZN(_11546_));
 XNOR2_X1 _34117_ (.A(_09227_),
    .B(_11461_),
    .ZN(_11547_));
 XOR2_X2 _34118_ (.A(_07276_),
    .B(_08729_),
    .Z(_11548_));
 XNOR2_X1 _34119_ (.A(_00348_),
    .B(_06714_),
    .ZN(_11549_));
 XNOR2_X1 _34120_ (.A(_11548_),
    .B(_11549_),
    .ZN(_11550_));
 XNOR2_X1 _34121_ (.A(_11547_),
    .B(_11550_),
    .ZN(_11551_));
 NAND2_X1 _34122_ (.A1(_10265_),
    .A2(_11551_),
    .ZN(_11552_));
 OAI21_X2 _34123_ (.A(_11552_),
    .B1(_07789_),
    .B2(_00432_),
    .ZN(_11553_));
 NAND2_X1 _34124_ (.A1(_09126_),
    .A2(_11553_),
    .ZN(_11554_));
 INV_X1 _34125_ (.A(\block_reg[3][19] ),
    .ZN(_11555_));
 OAI21_X1 _34126_ (.A(_11554_),
    .B1(_07248_),
    .B2(_11555_),
    .ZN(_11556_));
 OAI22_X1 _34127_ (.A1(\block_reg[3][19] ),
    .A2(_10794_),
    .B1(_10795_),
    .B2(_11553_),
    .ZN(_11557_));
 MUX2_X1 _34128_ (.A(_11556_),
    .B(_11557_),
    .S(_03298_),
    .Z(_11558_));
 NOR2_X1 _34129_ (.A1(_11415_),
    .A2(_11558_),
    .ZN(_11559_));
 AOI22_X1 _34130_ (.A1(_11546_),
    .A2(_11472_),
    .B1(_11559_),
    .B2(_08887_),
    .ZN(_00808_));
 BUF_X2 _34131_ (.A(\core.enc_block.block_w3_reg[25] ),
    .Z(_11560_));
 XNOR2_X2 _34132_ (.A(_11560_),
    .B(_08614_),
    .ZN(_11561_));
 XNOR2_X1 _34133_ (.A(_06737_),
    .B(_06861_),
    .ZN(_11562_));
 XNOR2_X2 _34134_ (.A(_11561_),
    .B(_11562_),
    .ZN(_11563_));
 XNOR2_X1 _34135_ (.A(_07294_),
    .B(_11419_),
    .ZN(_11564_));
 XNOR2_X1 _34136_ (.A(_11563_),
    .B(_11564_),
    .ZN(_11565_));
 MUX2_X1 _34137_ (.A(_06800_),
    .B(_11565_),
    .S(_07232_),
    .Z(_11566_));
 NAND2_X1 _34138_ (.A1(_09126_),
    .A2(_11566_),
    .ZN(_11567_));
 INV_X1 _34139_ (.A(\block_reg[3][1] ),
    .ZN(_11568_));
 OAI21_X1 _34140_ (.A(_11567_),
    .B1(_07248_),
    .B2(_11568_),
    .ZN(_11569_));
 OAI22_X1 _34141_ (.A1(\block_reg[3][1] ),
    .A2(_10794_),
    .B1(_10795_),
    .B2(_11566_),
    .ZN(_11570_));
 MUX2_X1 _34142_ (.A(_11569_),
    .B(_11570_),
    .S(_19284_),
    .Z(_11571_));
 NOR2_X1 _34143_ (.A1(_11415_),
    .A2(_11571_),
    .ZN(_11572_));
 AOI22_X1 _34144_ (.A1(_10671_),
    .A2(_11472_),
    .B1(_11572_),
    .B2(_08997_),
    .ZN(_00809_));
 XNOR2_X1 _34145_ (.A(_06768_),
    .B(_07319_),
    .ZN(_11573_));
 XOR2_X1 _34146_ (.A(_00331_),
    .B(_08905_),
    .Z(_11574_));
 XNOR2_X1 _34147_ (.A(_11573_),
    .B(_11574_),
    .ZN(_11575_));
 XNOR2_X1 _34148_ (.A(_11547_),
    .B(_11575_),
    .ZN(_11576_));
 NAND2_X1 _34149_ (.A1(_10717_),
    .A2(_11576_),
    .ZN(_11577_));
 OAI21_X2 _34150_ (.A(_11577_),
    .B1(_10948_),
    .B2(_00412_),
    .ZN(_11578_));
 OAI22_X1 _34151_ (.A1(\block_reg[3][20] ),
    .A2(_10232_),
    .B1(_11017_),
    .B2(_11578_),
    .ZN(_11579_));
 NAND2_X1 _34152_ (.A1(_10716_),
    .A2(_11578_),
    .ZN(_11580_));
 OAI21_X1 _34153_ (.A(_11580_),
    .B1(_10729_),
    .B2(_03699_),
    .ZN(_11581_));
 MUX2_X1 _34154_ (.A(_11579_),
    .B(_11581_),
    .S(_03710_),
    .Z(_11582_));
 NOR2_X1 _34155_ (.A1(_11440_),
    .A2(_11582_),
    .ZN(_11583_));
 AOI22_X1 _34156_ (.A1(_11225_),
    .A2(_11472_),
    .B1(_11583_),
    .B2(_09059_),
    .ZN(_00810_));
 INV_X1 _34157_ (.A(_11109_),
    .ZN(_11584_));
 NOR2_X1 _34158_ (.A1(\block_reg[3][21] ),
    .A2(_10729_),
    .ZN(_11585_));
 XNOR2_X1 _34159_ (.A(_07308_),
    .B(_09012_),
    .ZN(_11586_));
 XNOR2_X1 _34160_ (.A(_11474_),
    .B(_11586_),
    .ZN(_11587_));
 XNOR2_X1 _34161_ (.A(_07319_),
    .B(_11587_),
    .ZN(_11588_));
 MUX2_X1 _34162_ (.A(_00415_),
    .B(_11588_),
    .S(_07243_),
    .Z(_11589_));
 AOI21_X1 _34163_ (.A(_11585_),
    .B1(_11589_),
    .B2(_10696_),
    .ZN(_11590_));
 NAND2_X1 _34164_ (.A1(_18908_),
    .A2(_11590_),
    .ZN(_11591_));
 NAND2_X1 _34165_ (.A1(\block_reg[3][21] ),
    .A2(_09125_),
    .ZN(_11592_));
 OAI21_X1 _34166_ (.A(_11592_),
    .B1(_11589_),
    .B2(_08889_),
    .ZN(_11593_));
 OR2_X1 _34167_ (.A1(_18908_),
    .A2(_11593_),
    .ZN(_11594_));
 AOI21_X1 _34168_ (.A(_11486_),
    .B1(_11591_),
    .B2(_11594_),
    .ZN(_11595_));
 AOI22_X1 _34169_ (.A1(_11584_),
    .A2(_11472_),
    .B1(_11595_),
    .B2(_09124_),
    .ZN(_00811_));
 XNOR2_X2 _34170_ (.A(_07308_),
    .B(_09139_),
    .ZN(_11596_));
 XNOR2_X1 _34171_ (.A(_11488_),
    .B(_11596_),
    .ZN(_11597_));
 XNOR2_X1 _34172_ (.A(_07331_),
    .B(_11597_),
    .ZN(_11598_));
 NAND2_X1 _34173_ (.A1(_08722_),
    .A2(_11598_),
    .ZN(_11599_));
 OAI21_X1 _34174_ (.A(_11599_),
    .B1(_07243_),
    .B2(_00418_),
    .ZN(_11600_));
 OAI22_X1 _34175_ (.A1(\block_reg[3][22] ),
    .A2(_09134_),
    .B1(_09222_),
    .B2(_11600_),
    .ZN(_11601_));
 NOR2_X1 _34176_ (.A1(_18920_),
    .A2(_11601_),
    .ZN(_11602_));
 AOI22_X1 _34177_ (.A1(\block_reg[3][22] ),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_11600_),
    .ZN(_11603_));
 AOI21_X2 _34178_ (.A(_11602_),
    .B1(_11603_),
    .B2(_18920_),
    .ZN(_11604_));
 NOR3_X1 _34179_ (.A1(_09172_),
    .A2(_11440_),
    .A3(_11604_),
    .ZN(_11605_));
 INV_X1 _34180_ (.A(_11123_),
    .ZN(_11606_));
 AOI21_X1 _34181_ (.A(_11605_),
    .B1(_11414_),
    .B2(_11606_),
    .ZN(_00812_));
 INV_X1 _34182_ (.A(_11136_),
    .ZN(_11607_));
 XNOR2_X2 _34183_ (.A(_07331_),
    .B(_09183_),
    .ZN(_11608_));
 XNOR2_X1 _34184_ (.A(_11442_),
    .B(_11608_),
    .ZN(_11609_));
 XNOR2_X1 _34185_ (.A(_11417_),
    .B(_11609_),
    .ZN(_11610_));
 NAND2_X1 _34186_ (.A1(_10354_),
    .A2(_11610_),
    .ZN(_11611_));
 OAI21_X2 _34187_ (.A(_11611_),
    .B1(_07801_),
    .B2(_00421_),
    .ZN(_11612_));
 OAI221_X2 _34188_ (.A(_18955_),
    .B1(_07893_),
    .B2(_11612_),
    .C1(_07906_),
    .C2(\block_reg[3][23] ),
    .ZN(_11613_));
 NAND2_X1 _34189_ (.A1(_09211_),
    .A2(_11612_),
    .ZN(_11614_));
 OAI21_X1 _34190_ (.A(_11614_),
    .B1(_08888_),
    .B2(_03956_),
    .ZN(_11615_));
 OR2_X1 _34191_ (.A1(_18955_),
    .A2(_11615_),
    .ZN(_11616_));
 AOI21_X2 _34192_ (.A(_11486_),
    .B1(_11613_),
    .B2(_11616_),
    .ZN(_11617_));
 AOI22_X1 _34193_ (.A1(_11607_),
    .A2(_11472_),
    .B1(_11617_),
    .B2(_09210_),
    .ZN(_00813_));
 INV_X1 _34194_ (.A(_11418_),
    .ZN(_11618_));
 XNOR2_X1 _34195_ (.A(_11420_),
    .B(_11499_),
    .ZN(_11619_));
 XNOR2_X1 _34196_ (.A(_06861_),
    .B(_11619_),
    .ZN(_11620_));
 NAND2_X1 _34197_ (.A1(_10717_),
    .A2(_11620_),
    .ZN(_11621_));
 OAI21_X2 _34198_ (.A(_11621_),
    .B1(_10948_),
    .B2(_00341_),
    .ZN(_11622_));
 OAI22_X1 _34199_ (.A1(\block_reg[3][24] ),
    .A2(_10232_),
    .B1(_07254_),
    .B2(_11622_),
    .ZN(_11623_));
 NAND2_X1 _34200_ (.A1(_10716_),
    .A2(_11622_),
    .ZN(_11624_));
 OAI21_X1 _34201_ (.A(_11624_),
    .B1(_10729_),
    .B2(_06546_),
    .ZN(_11625_));
 MUX2_X1 _34202_ (.A(_11623_),
    .B(_11625_),
    .S(_18981_),
    .Z(_11626_));
 NOR2_X1 _34203_ (.A1(_11440_),
    .A2(_11626_),
    .ZN(_11627_));
 AOI22_X1 _34204_ (.A1(_11618_),
    .A2(_11472_),
    .B1(_11627_),
    .B2(_09682_),
    .ZN(_00814_));
 INV_X1 _34205_ (.A(_11560_),
    .ZN(_11628_));
 AND2_X1 _34206_ (.A1(_00344_),
    .A2(_10223_),
    .ZN(_11629_));
 XNOR2_X1 _34207_ (.A(_00426_),
    .B(_11419_),
    .ZN(_11630_));
 XNOR2_X1 _34208_ (.A(_11525_),
    .B(_11630_),
    .ZN(_11631_));
 AOI21_X2 _34209_ (.A(_11629_),
    .B1(_11631_),
    .B2(_09217_),
    .ZN(_11632_));
 OAI221_X1 _34210_ (.A(_19298_),
    .B1(_07893_),
    .B2(_11632_),
    .C1(_07906_),
    .C2(\block_reg[3][25] ),
    .ZN(_11633_));
 NAND2_X1 _34211_ (.A1(_09211_),
    .A2(_11632_),
    .ZN(_11634_));
 INV_X1 _34212_ (.A(\block_reg[3][25] ),
    .ZN(_11635_));
 OAI21_X1 _34213_ (.A(_11634_),
    .B1(_08888_),
    .B2(_11635_),
    .ZN(_11636_));
 OR2_X1 _34214_ (.A1(_19298_),
    .A2(_11636_),
    .ZN(_11637_));
 AOI21_X1 _34215_ (.A(_11486_),
    .B1(_11633_),
    .B2(_11637_),
    .ZN(_11638_));
 AOI22_X1 _34216_ (.A1(_11628_),
    .A2(_11415_),
    .B1(_11638_),
    .B2(_09778_),
    .ZN(_00815_));
 XOR2_X1 _34217_ (.A(_11548_),
    .B(_11561_),
    .Z(_11639_));
 XNOR2_X1 _34218_ (.A(_06788_),
    .B(_11639_),
    .ZN(_11640_));
 MUX2_X1 _34219_ (.A(\core.enc_block.block_w3_reg[26] ),
    .B(_11640_),
    .S(_09131_),
    .Z(_11641_));
 AOI22_X1 _34220_ (.A1(\block_reg[3][26] ),
    .A2(_07805_),
    .B1(_10956_),
    .B2(_11641_),
    .ZN(_11642_));
 INV_X1 _34221_ (.A(_11642_),
    .ZN(_11643_));
 OAI22_X1 _34222_ (.A1(\block_reg[3][26] ),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_11641_),
    .ZN(_11644_));
 MUX2_X1 _34223_ (.A(_11643_),
    .B(_11644_),
    .S(_19428_),
    .Z(_11645_));
 NOR3_X1 _34224_ (.A1(_09860_),
    .A2(_11413_),
    .A3(_11645_),
    .ZN(_11646_));
 AOI21_X1 _34225_ (.A(_11646_),
    .B1(_11414_),
    .B2(_09245_),
    .ZN(_00816_));
 XNOR2_X1 _34226_ (.A(_00432_),
    .B(_08729_),
    .ZN(_11647_));
 XNOR2_X1 _34227_ (.A(_11499_),
    .B(_11647_),
    .ZN(_11648_));
 XNOR2_X1 _34228_ (.A(_06714_),
    .B(_07285_),
    .ZN(_11649_));
 XNOR2_X1 _34229_ (.A(_09245_),
    .B(_11649_),
    .ZN(_11650_));
 XNOR2_X1 _34230_ (.A(_11648_),
    .B(_11650_),
    .ZN(_11651_));
 MUX2_X1 _34231_ (.A(_11443_),
    .B(_11651_),
    .S(_09131_),
    .Z(_11652_));
 AOI22_X1 _34232_ (.A1(\block_reg[3][27] ),
    .A2(_07805_),
    .B1(_10956_),
    .B2(_11652_),
    .ZN(_11653_));
 INV_X1 _34233_ (.A(_11653_),
    .ZN(_11654_));
 OAI22_X1 _34234_ (.A1(\block_reg[3][27] ),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_11652_),
    .ZN(_11655_));
 MUX2_X1 _34235_ (.A(_11654_),
    .B(_11655_),
    .S(_03325_),
    .Z(_11656_));
 NOR3_X1 _34236_ (.A1(_09950_),
    .A2(_11413_),
    .A3(_11656_),
    .ZN(_11657_));
 INV_X1 _34237_ (.A(_11443_),
    .ZN(_11658_));
 AOI21_X1 _34238_ (.A(_11657_),
    .B1(_11414_),
    .B2(_11658_),
    .ZN(_00817_));
 XOR2_X1 _34239_ (.A(_11499_),
    .B(_11573_),
    .Z(_11659_));
 XNOR2_X1 _34240_ (.A(_00412_),
    .B(_11444_),
    .ZN(_11660_));
 XNOR2_X1 _34241_ (.A(_11659_),
    .B(_11660_),
    .ZN(_11661_));
 NAND2_X1 _34242_ (.A1(_08809_),
    .A2(_11661_),
    .ZN(_11662_));
 OAI21_X1 _34243_ (.A(_11662_),
    .B1(_10265_),
    .B2(_00331_),
    .ZN(_11663_));
 AOI22_X1 _34244_ (.A1(\block_reg[3][28] ),
    .A2(_07805_),
    .B1(_10956_),
    .B2(_11663_),
    .ZN(_11664_));
 INV_X1 _34245_ (.A(_11664_),
    .ZN(_11665_));
 OAI22_X1 _34246_ (.A1(\block_reg[3][28] ),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_11663_),
    .ZN(_11666_));
 MUX2_X1 _34247_ (.A(_11665_),
    .B(_11666_),
    .S(_03738_),
    .Z(_11667_));
 NOR3_X1 _34248_ (.A1(_10010_),
    .A2(_11413_),
    .A3(_11667_),
    .ZN(_11668_));
 INV_X1 _34249_ (.A(_11457_),
    .ZN(_11669_));
 AOI21_X1 _34250_ (.A(_11668_),
    .B1(_11414_),
    .B2(_11669_),
    .ZN(_00818_));
 INV_X1 _34251_ (.A(_11473_),
    .ZN(_11670_));
 XNOR2_X1 _34252_ (.A(_11458_),
    .B(_11596_),
    .ZN(_11671_));
 XNOR2_X1 _34253_ (.A(_06761_),
    .B(_11671_),
    .ZN(_11672_));
 NAND2_X1 _34254_ (.A1(_09217_),
    .A2(_11672_),
    .ZN(_11673_));
 OAI21_X1 _34255_ (.A(_11673_),
    .B1(_10172_),
    .B2(_00334_),
    .ZN(_11674_));
 OAI22_X1 _34256_ (.A1(\block_reg[3][29] ),
    .A2(_07905_),
    .B1(_08889_),
    .B2(_11674_),
    .ZN(_11675_));
 OR2_X1 _34257_ (.A1(_19001_),
    .A2(_11675_),
    .ZN(_11676_));
 AOI22_X1 _34258_ (.A1(\block_reg[3][29] ),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_11674_),
    .ZN(_11677_));
 NAND2_X1 _34259_ (.A1(_19001_),
    .A2(_11677_),
    .ZN(_11678_));
 AOI21_X1 _34260_ (.A(_11486_),
    .B1(_11676_),
    .B2(_11678_),
    .ZN(_11679_));
 AOI22_X1 _34261_ (.A1(_11670_),
    .A2(_11415_),
    .B1(_11679_),
    .B2(_10076_),
    .ZN(_00819_));
 INV_X1 _34262_ (.A(_07648_),
    .ZN(_11680_));
 XNOR2_X1 _34263_ (.A(_06800_),
    .B(_11560_),
    .ZN(_11681_));
 XNOR2_X1 _34264_ (.A(_11548_),
    .B(_11681_),
    .ZN(_11682_));
 XNOR2_X1 _34265_ (.A(_09245_),
    .B(_11682_),
    .ZN(_11683_));
 MUX2_X1 _34266_ (.A(_06788_),
    .B(_11683_),
    .S(_08722_),
    .Z(_11684_));
 OAI221_X1 _34267_ (.A(_19457_),
    .B1(_07893_),
    .B2(_11684_),
    .C1(_07906_),
    .C2(\block_reg[3][2] ),
    .ZN(_11685_));
 NAND2_X1 _34268_ (.A1(_09211_),
    .A2(_11684_),
    .ZN(_11686_));
 INV_X1 _34269_ (.A(\block_reg[3][2] ),
    .ZN(_11687_));
 OAI21_X1 _34270_ (.A(_11686_),
    .B1(_07905_),
    .B2(_11687_),
    .ZN(_11688_));
 OR2_X1 _34271_ (.A1(_19457_),
    .A2(_11688_),
    .ZN(_11689_));
 AOI21_X1 _34272_ (.A(_11486_),
    .B1(_11685_),
    .B2(_11689_),
    .ZN(_11690_));
 AOI22_X1 _34273_ (.A1(_11680_),
    .A2(_11415_),
    .B1(_11690_),
    .B2(_10168_),
    .ZN(_00820_));
 INV_X1 _34274_ (.A(\block_reg[3][30] ),
    .ZN(_11691_));
 XOR2_X1 _34275_ (.A(_11473_),
    .B(_09139_),
    .Z(_11692_));
 XNOR2_X1 _34276_ (.A(_11608_),
    .B(_11692_),
    .ZN(_11693_));
 XNOR2_X1 _34277_ (.A(_06748_),
    .B(_11693_),
    .ZN(_11694_));
 MUX2_X1 _34278_ (.A(_00337_),
    .B(_11694_),
    .S(_07651_),
    .Z(_11695_));
 OAI22_X1 _34279_ (.A1(_11691_),
    .A2(_09134_),
    .B1(_09222_),
    .B2(_11695_),
    .ZN(_11696_));
 NOR2_X1 _34280_ (.A1(_19245_),
    .A2(_11696_),
    .ZN(_11697_));
 AOI22_X1 _34281_ (.A1(_11691_),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_11695_),
    .ZN(_11698_));
 AOI21_X1 _34282_ (.A(_11697_),
    .B1(_11698_),
    .B2(_19245_),
    .ZN(_11699_));
 NOR3_X1 _34283_ (.A1(_10222_),
    .A2(_11413_),
    .A3(_11699_),
    .ZN(_11700_));
 INV_X1 _34284_ (.A(_11487_),
    .ZN(_11701_));
 AOI21_X1 _34285_ (.A(_11700_),
    .B1(_11414_),
    .B2(_11701_),
    .ZN(_00821_));
 XOR2_X1 _34286_ (.A(_09183_),
    .B(_09227_),
    .Z(_11702_));
 XNOR2_X1 _34287_ (.A(_11442_),
    .B(_11702_),
    .ZN(_11703_));
 XNOR2_X1 _34288_ (.A(_11701_),
    .B(_11703_),
    .ZN(_11704_));
 NOR2_X1 _34289_ (.A1(_10223_),
    .A2(_11704_),
    .ZN(_11705_));
 AOI21_X2 _34290_ (.A(_11705_),
    .B1(_10223_),
    .B2(_00340_),
    .ZN(_11706_));
 NAND2_X1 _34291_ (.A1(_07808_),
    .A2(_11706_),
    .ZN(_11707_));
 INV_X1 _34292_ (.A(\block_reg[3][31] ),
    .ZN(_11708_));
 OAI21_X1 _34293_ (.A(_11707_),
    .B1(_07251_),
    .B2(_11708_),
    .ZN(_11709_));
 OAI22_X1 _34294_ (.A1(\block_reg[3][31] ),
    .A2(_08104_),
    .B1(_08105_),
    .B2(_11706_),
    .ZN(_11710_));
 MUX2_X1 _34295_ (.A(_11709_),
    .B(_11710_),
    .S(_19440_),
    .Z(_11711_));
 NOR3_X1 _34296_ (.A1(_10261_),
    .A2(_11413_),
    .A3(_11711_),
    .ZN(_11712_));
 INV_X1 _34297_ (.A(_11417_),
    .ZN(_11713_));
 AOI21_X1 _34298_ (.A(_11712_),
    .B1(_11414_),
    .B2(_11713_),
    .ZN(_00822_));
 INV_X1 _34299_ (.A(_07790_),
    .ZN(_11714_));
 XNOR2_X1 _34300_ (.A(_11430_),
    .B(_11444_),
    .ZN(_11715_));
 XNOR2_X1 _34301_ (.A(_11417_),
    .B(_00303_),
    .ZN(_11716_));
 XNOR2_X1 _34302_ (.A(_06737_),
    .B(_11716_),
    .ZN(_11717_));
 XNOR2_X1 _34303_ (.A(_11715_),
    .B(_11717_),
    .ZN(_11718_));
 MUX2_X2 _34304_ (.A(_06714_),
    .B(_11718_),
    .S(_07243_),
    .Z(_11719_));
 OAI221_X1 _34305_ (.A(_03357_),
    .B1(_07893_),
    .B2(_11719_),
    .C1(_07906_),
    .C2(\block_reg[3][3] ),
    .ZN(_11720_));
 AOI22_X1 _34306_ (.A1(\block_reg[3][3] ),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_11719_),
    .ZN(_11721_));
 OAI21_X1 _34307_ (.A(_11721_),
    .B1(_03356_),
    .B2(_03355_),
    .ZN(_11722_));
 AOI21_X1 _34308_ (.A(_11486_),
    .B1(_11720_),
    .B2(_11722_),
    .ZN(_11723_));
 AOI22_X1 _34309_ (.A1(_11714_),
    .A2(_11415_),
    .B1(_11723_),
    .B2(_10353_),
    .ZN(_00823_));
 INV_X1 _34310_ (.A(_07897_),
    .ZN(_11724_));
 XNOR2_X1 _34311_ (.A(_11443_),
    .B(_00304_),
    .ZN(_11725_));
 XNOR2_X1 _34312_ (.A(_11713_),
    .B(_11725_),
    .ZN(_11726_));
 XNOR2_X1 _34313_ (.A(_11460_),
    .B(_11726_),
    .ZN(_11727_));
 MUX2_X2 _34314_ (.A(_06768_),
    .B(_11727_),
    .S(_07243_),
    .Z(_11728_));
 OAI221_X1 _34315_ (.A(_03759_),
    .B1(_07893_),
    .B2(_11728_),
    .C1(_07906_),
    .C2(\block_reg[3][4] ),
    .ZN(_11729_));
 AOI22_X1 _34316_ (.A1(\block_reg[3][4] ),
    .A2(_08116_),
    .B1(_08117_),
    .B2(_11728_),
    .ZN(_11730_));
 OAI21_X1 _34317_ (.A(_11730_),
    .B1(_03758_),
    .B2(_03757_),
    .ZN(_11731_));
 AOI21_X1 _34318_ (.A(_11486_),
    .B1(_11729_),
    .B2(_11731_),
    .ZN(_11732_));
 AOI22_X1 _34319_ (.A1(_11724_),
    .A2(_11415_),
    .B1(_11732_),
    .B2(_10414_),
    .ZN(_00824_));
 INV_X1 _34320_ (.A(_08043_),
    .ZN(_11733_));
 NOR2_X1 _34321_ (.A1(_06761_),
    .A2(_08896_),
    .ZN(_11734_));
 XOR2_X1 _34322_ (.A(_11457_),
    .B(_11473_),
    .Z(_11735_));
 XNOR2_X1 _34323_ (.A(_11596_),
    .B(_11735_),
    .ZN(_11736_));
 XNOR2_X1 _34324_ (.A(_06768_),
    .B(_11736_),
    .ZN(_11737_));
 AOI21_X2 _34325_ (.A(_11734_),
    .B1(_11737_),
    .B2(_08048_),
    .ZN(_11738_));
 OAI22_X1 _34326_ (.A1(\block_reg[3][5] ),
    .A2(_10232_),
    .B1(_07254_),
    .B2(_11738_),
    .ZN(_11739_));
 NAND2_X1 _34327_ (.A1(_10716_),
    .A2(_11738_),
    .ZN(_11740_));
 OAI21_X1 _34328_ (.A(_11740_),
    .B1(_10729_),
    .B2(_06362_),
    .ZN(_11741_));
 MUX2_X1 _34329_ (.A(_11739_),
    .B(_11741_),
    .S(_18895_),
    .Z(_11742_));
 NOR2_X1 _34330_ (.A1(_11440_),
    .A2(_11742_),
    .ZN(_11743_));
 AOI22_X1 _34331_ (.A1(_11733_),
    .A2(_11415_),
    .B1(_11743_),
    .B2(_10470_),
    .ZN(_00825_));
 XOR2_X1 _34332_ (.A(_11474_),
    .B(_11608_),
    .Z(_11744_));
 XNOR2_X1 _34333_ (.A(_11487_),
    .B(_11744_),
    .ZN(_11745_));
 MUX2_X1 _34334_ (.A(_06748_),
    .B(_11745_),
    .S(_08038_),
    .Z(_11746_));
 AOI22_X1 _34335_ (.A1(\block_reg[3][6] ),
    .A2(_09125_),
    .B1(_07229_),
    .B2(_11746_),
    .ZN(_11747_));
 OAI22_X1 _34336_ (.A1(\block_reg[3][6] ),
    .A2(_07904_),
    .B1(_09007_),
    .B2(_11746_),
    .ZN(_11748_));
 INV_X1 _34337_ (.A(_11748_),
    .ZN(_11749_));
 MUX2_X1 _34338_ (.A(_11747_),
    .B(_11749_),
    .S(_18883_),
    .Z(_11750_));
 NAND2_X1 _34339_ (.A1(_10527_),
    .A2(_11750_),
    .ZN(_11751_));
 MUX2_X1 _34340_ (.A(_11751_),
    .B(_08110_),
    .S(_11440_),
    .Z(_00826_));
 INV_X1 _34341_ (.A(_07791_),
    .ZN(_11752_));
 XNOR2_X1 _34342_ (.A(_11488_),
    .B(_11499_),
    .ZN(_11753_));
 XNOR2_X1 _34343_ (.A(_07340_),
    .B(_11753_),
    .ZN(_11754_));
 NAND2_X1 _34344_ (.A1(_09217_),
    .A2(_11754_),
    .ZN(_11755_));
 OAI21_X1 _34345_ (.A(_11755_),
    .B1(_10172_),
    .B2(_00302_),
    .ZN(_11756_));
 OAI22_X1 _34346_ (.A1(\block_reg[3][7] ),
    .A2(_07905_),
    .B1(_07788_),
    .B2(_11756_),
    .ZN(_11757_));
 OR2_X1 _34347_ (.A1(_19259_),
    .A2(_11757_),
    .ZN(_11758_));
 AOI22_X1 _34348_ (.A1(\block_reg[3][7] ),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_11756_),
    .ZN(_11759_));
 NAND2_X1 _34349_ (.A1(_19259_),
    .A2(_11759_),
    .ZN(_11760_));
 AOI21_X1 _34350_ (.A(_11412_),
    .B1(_11758_),
    .B2(_11760_),
    .ZN(_11761_));
 AOI22_X1 _34351_ (.A1(_11752_),
    .A2(_11415_),
    .B1(_11761_),
    .B2(_10566_),
    .ZN(_00827_));
 XNOR2_X1 _34352_ (.A(_11442_),
    .B(_11510_),
    .ZN(_11762_));
 XNOR2_X1 _34353_ (.A(_08612_),
    .B(_11762_),
    .ZN(_11763_));
 MUX2_X1 _34354_ (.A(_07267_),
    .B(_11763_),
    .S(_08038_),
    .Z(_11764_));
 AOI22_X1 _34355_ (.A1(\block_reg[3][8] ),
    .A2(_07806_),
    .B1(_07229_),
    .B2(_11764_),
    .ZN(_11765_));
 OAI22_X1 _34356_ (.A1(\block_reg[3][8] ),
    .A2(_07904_),
    .B1(_07253_),
    .B2(_11764_),
    .ZN(_11766_));
 INV_X1 _34357_ (.A(_11766_),
    .ZN(_11767_));
 MUX2_X1 _34358_ (.A(_11765_),
    .B(_11767_),
    .S(_19015_),
    .Z(_11768_));
 NAND2_X1 _34359_ (.A1(_10614_),
    .A2(_11768_),
    .ZN(_11769_));
 MUX2_X1 _34360_ (.A(_11769_),
    .B(\core.enc_block.block_w3_reg[8] ),
    .S(_11440_),
    .Z(_00828_));
 XNOR2_X1 _34361_ (.A(_06800_),
    .B(_11509_),
    .ZN(_11770_));
 XNOR2_X1 _34362_ (.A(_11563_),
    .B(_11770_),
    .ZN(_11771_));
 NAND2_X1 _34363_ (.A1(_08722_),
    .A2(_11771_),
    .ZN(_11772_));
 OAI21_X1 _34364_ (.A(_11772_),
    .B1(_07243_),
    .B2(_00305_),
    .ZN(_11773_));
 OAI22_X1 _34365_ (.A1(\block_reg[3][9] ),
    .A2(_09134_),
    .B1(_09222_),
    .B2(_11773_),
    .ZN(_11774_));
 NOR2_X1 _34366_ (.A1(_19273_),
    .A2(_11774_),
    .ZN(_11775_));
 AOI22_X1 _34367_ (.A1(\block_reg[3][9] ),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_11773_),
    .ZN(_11776_));
 AOI21_X1 _34368_ (.A(_11775_),
    .B1(_11776_),
    .B2(_19273_),
    .ZN(_11777_));
 NOR3_X2 _34369_ (.A1(_10670_),
    .A2(_11413_),
    .A3(_11777_),
    .ZN(_11778_));
 INV_X1 _34370_ (.A(_10796_),
    .ZN(_11779_));
 AOI21_X1 _34371_ (.A(_11778_),
    .B1(_11414_),
    .B2(_11779_),
    .ZN(_00829_));
 INV_X1 _34372_ (.A(\core.enc_block.ready ),
    .ZN(_11780_));
 OAI21_X1 _34373_ (.A(_16246_),
    .B1(_16241_),
    .B2(_11780_),
    .ZN(_00830_));
 XNOR2_X1 _34374_ (.A(_16409_),
    .B(_16249_),
    .ZN(_11781_));
 NOR2_X1 _34375_ (.A1(_16241_),
    .A2(_11781_),
    .ZN(_00831_));
 NAND2_X1 _34376_ (.A1(_16236_),
    .A2(_16249_),
    .ZN(_11782_));
 OAI21_X1 _34377_ (.A(_22115_),
    .B1(_16232_),
    .B2(_16234_),
    .ZN(_11783_));
 AOI21_X1 _34378_ (.A(_16241_),
    .B1(_11782_),
    .B2(_11783_),
    .ZN(_00832_));
 OAI21_X1 _34379_ (.A(_22114_),
    .B1(_16232_),
    .B2(_16234_),
    .ZN(_11784_));
 XNOR2_X1 _34380_ (.A(_16426_),
    .B(_11784_),
    .ZN(_11785_));
 NOR2_X1 _34381_ (.A1(_16241_),
    .A2(_11785_),
    .ZN(_00833_));
 NAND3_X1 _34382_ (.A1(_16236_),
    .A2(_16373_),
    .A3(_16380_),
    .ZN(_11786_));
 XNOR2_X1 _34383_ (.A(_00323_),
    .B(_11786_),
    .ZN(_11787_));
 MUX2_X1 _34384_ (.A(_11787_),
    .B(_16477_),
    .S(_16249_),
    .Z(_11788_));
 NOR2_X1 _34385_ (.A1(_16241_),
    .A2(_11788_),
    .ZN(_00834_));
 NOR3_X1 _34386_ (.A1(_06693_),
    .A2(_16239_),
    .A3(\core.enc_block.sword_ctr_reg[0] ),
    .ZN(_11789_));
 AOI21_X1 _34387_ (.A(_11789_),
    .B1(\core.enc_block.sword_ctr_reg[0] ),
    .B2(_16239_),
    .ZN(_11790_));
 NOR3_X1 _34388_ (.A1(_16234_),
    .A2(_16232_),
    .A3(_11790_),
    .ZN(_00835_));
 MUX2_X1 _34389_ (.A(_22119_),
    .B(\core.enc_block.sword_ctr_reg[1] ),
    .S(_16239_),
    .Z(_11791_));
 AND2_X1 _34390_ (.A1(_16249_),
    .A2(_11791_),
    .ZN(_00836_));
 INV_X4 _34391_ (.A(_00318_),
    .ZN(_11792_));
 BUF_X4 _34392_ (.A(_22106_),
    .Z(_11793_));
 BUF_X4 _34393_ (.A(\core.keymem.round_ctr_reg[3] ),
    .Z(_11794_));
 NOR2_X4 _34394_ (.A1(_11794_),
    .A2(_16218_),
    .ZN(_11795_));
 AND2_X1 _34395_ (.A1(_11793_),
    .A2(_11795_),
    .ZN(_11796_));
 BUF_X4 _34396_ (.A(_11796_),
    .Z(_11797_));
 BUF_X4 _34397_ (.A(_11797_),
    .Z(_11798_));
 BUF_X4 _34398_ (.A(_11798_),
    .Z(_11799_));
 BUF_X8 _34399_ (.A(_11799_),
    .Z(_11800_));
 NAND2_X4 _34400_ (.A1(_11792_),
    .A2(_11800_),
    .ZN(_11801_));
 BUF_X8 _34401_ (.A(_11801_),
    .Z(_11802_));
 INV_X2 _34402_ (.A(_16222_),
    .ZN(_11803_));
 BUF_X8 _34403_ (.A(_11803_),
    .Z(_11804_));
 BUF_X4 _34404_ (.A(_11804_),
    .Z(_11805_));
 NOR2_X4 _34405_ (.A1(_11805_),
    .A2(_11801_),
    .ZN(_11806_));
 XOR2_X2 _34406_ (.A(\core.keymem.prev_key1_reg[32] ),
    .B(\core.keymem.prev_key1_reg[64] ),
    .Z(_11807_));
 XNOR2_X1 _34407_ (.A(_06858_),
    .B(_00328_),
    .ZN(_11808_));
 XNOR2_X1 _34408_ (.A(_11807_),
    .B(_11808_),
    .ZN(_11809_));
 XNOR2_X1 _34409_ (.A(_09681_),
    .B(_11809_),
    .ZN(_11810_));
 INV_X8 _34410_ (.A(_16219_),
    .ZN(_11811_));
 BUF_X8 _34411_ (.A(_11795_),
    .Z(_11812_));
 NAND2_X4 _34412_ (.A1(_11793_),
    .A2(_11812_),
    .ZN(_11813_));
 NAND2_X4 _34413_ (.A1(_11811_),
    .A2(_11813_),
    .ZN(_11814_));
 NOR2_X1 _34414_ (.A1(_11810_),
    .A2(_11814_),
    .ZN(_11815_));
 BUF_X4 _34415_ (.A(_22110_),
    .Z(_11816_));
 AND2_X1 _34416_ (.A1(_11816_),
    .A2(_11795_),
    .ZN(_11817_));
 BUF_X4 _34417_ (.A(_11817_),
    .Z(_11818_));
 BUF_X4 _34418_ (.A(_11818_),
    .Z(_11819_));
 BUF_X4 _34419_ (.A(_11819_),
    .Z(_11820_));
 NAND2_X1 _34420_ (.A1(\core.key[0] ),
    .A2(_11820_),
    .ZN(_11821_));
 NOR2_X4 _34421_ (.A1(_11811_),
    .A2(_11797_),
    .ZN(_11822_));
 BUF_X4 _34422_ (.A(_11822_),
    .Z(_11823_));
 AND2_X1 _34423_ (.A1(_11821_),
    .A2(_11823_),
    .ZN(_11824_));
 NAND2_X4 _34424_ (.A1(_11816_),
    .A2(_11795_),
    .ZN(_11825_));
 BUF_X4 _34425_ (.A(_11825_),
    .Z(_11826_));
 BUF_X4 _34426_ (.A(_11826_),
    .Z(_11827_));
 BUF_X4 _34427_ (.A(_11827_),
    .Z(_11828_));
 BUF_X4 _34428_ (.A(\core.keymem.round_ctr_reg[0] ),
    .Z(_11829_));
 CLKBUF_X3 _34429_ (.A(_11829_),
    .Z(_11830_));
 BUF_X4 _34430_ (.A(_11830_),
    .Z(_11831_));
 BUF_X4 _34431_ (.A(_11831_),
    .Z(_11832_));
 NAND4_X1 _34432_ (.A1(_11831_),
    .A2(_07116_),
    .A3(_07171_),
    .A4(_07220_),
    .ZN(_11833_));
 OAI33_X1 _34433_ (.A1(_11832_),
    .A2(_09569_),
    .A3(_09680_),
    .B1(_11833_),
    .B2(_07073_),
    .B3(_07044_),
    .ZN(_11834_));
 XNOR2_X2 _34434_ (.A(\core.keymem.prev_key0_reg[96] ),
    .B(net12),
    .ZN(_11835_));
 XNOR2_X2 _34435_ (.A(\core.keymem.prev_key0_reg[32] ),
    .B(\core.keymem.prev_key0_reg[64] ),
    .ZN(_11836_));
 XOR2_X1 _34436_ (.A(\core.keymem.prev_key0_reg[0] ),
    .B(_11836_),
    .Z(_11837_));
 XNOR2_X1 _34437_ (.A(_11835_),
    .B(_11837_),
    .ZN(_11838_));
 NAND2_X1 _34438_ (.A1(_11828_),
    .A2(_11838_),
    .ZN(_11839_));
 BUF_X4 _34439_ (.A(_11797_),
    .Z(_11840_));
 BUF_X4 _34440_ (.A(_11840_),
    .Z(_11841_));
 BUF_X8 _34441_ (.A(_11841_),
    .Z(_11842_));
 AOI221_X2 _34442_ (.A(_11815_),
    .B1(_11824_),
    .B2(_11839_),
    .C1(_00327_),
    .C2(_11842_),
    .ZN(_11843_));
 BUF_X2 _34443_ (.A(_11843_),
    .Z(_11844_));
 AOI22_X1 _34444_ (.A1(\core.keymem.key_mem[0][0] ),
    .A2(_11802_),
    .B1(_11806_),
    .B2(_11844_),
    .ZN(_11845_));
 INV_X1 _34445_ (.A(_11845_),
    .ZN(_00837_));
 BUF_X4 _34446_ (.A(_11811_),
    .Z(_11846_));
 BUF_X8 _34447_ (.A(_11846_),
    .Z(_11847_));
 BUF_X4 _34448_ (.A(_11826_),
    .Z(_11848_));
 NOR2_X1 _34449_ (.A1(\core.key[100] ),
    .A2(_11848_),
    .ZN(_11849_));
 INV_X4 _34450_ (.A(_11829_),
    .ZN(_11850_));
 BUF_X4 _34451_ (.A(_11850_),
    .Z(_11851_));
 OR2_X1 _34452_ (.A1(_09570_),
    .A2(_09964_),
    .ZN(_11852_));
 OAI21_X1 _34453_ (.A(_11852_),
    .B1(_09973_),
    .B2(_09660_),
    .ZN(_11853_));
 AND4_X1 _34454_ (.A1(_09670_),
    .A2(_09988_),
    .A3(_10000_),
    .A4(_10007_),
    .ZN(_11854_));
 NAND3_X2 _34455_ (.A1(_11851_),
    .A2(_11853_),
    .A3(_11854_),
    .ZN(_11855_));
 BUF_X4 _34456_ (.A(_11850_),
    .Z(_11856_));
 BUF_X4 _34457_ (.A(_11856_),
    .Z(_11857_));
 OAI21_X4 _34458_ (.A(_11855_),
    .B1(_10413_),
    .B2(_11857_),
    .ZN(_11858_));
 XOR2_X2 _34459_ (.A(\core.keymem.prev_key0_reg[100] ),
    .B(_11858_),
    .Z(_11859_));
 BUF_X4 _34460_ (.A(_11826_),
    .Z(_11860_));
 AOI221_X2 _34461_ (.A(_11849_),
    .B1(_11859_),
    .B2(_11860_),
    .C1(_11793_),
    .C2(_11812_),
    .ZN(_11861_));
 BUF_X4 _34462_ (.A(_11813_),
    .Z(_11862_));
 BUF_X4 _34463_ (.A(_11862_),
    .Z(_11863_));
 NOR2_X1 _34464_ (.A1(_00127_),
    .A2(_11863_),
    .ZN(_11864_));
 NOR3_X2 _34465_ (.A1(_11847_),
    .A2(_11861_),
    .A3(_11864_),
    .ZN(_11865_));
 BUF_X8 _34466_ (.A(_11846_),
    .Z(_11866_));
 XNOR2_X1 _34467_ (.A(_00128_),
    .B(_10009_),
    .ZN(_11867_));
 BUF_X4 _34468_ (.A(_11813_),
    .Z(_11868_));
 MUX2_X1 _34469_ (.A(_00127_),
    .B(_11867_),
    .S(_11868_),
    .Z(_11869_));
 NAND2_X1 _34470_ (.A1(_11866_),
    .A2(_11869_),
    .ZN(_11870_));
 NAND2_X1 _34471_ (.A1(_16228_),
    .A2(_11870_),
    .ZN(_11871_));
 NOR2_X4 _34472_ (.A1(_11865_),
    .A2(_11871_),
    .ZN(_11872_));
 BUF_X2 _34473_ (.A(_11872_),
    .Z(_11873_));
 BUF_X8 _34474_ (.A(_11813_),
    .Z(_11874_));
 BUF_X4 _34475_ (.A(_11874_),
    .Z(_11875_));
 NOR2_X2 _34476_ (.A1(_16224_),
    .A2(_11875_),
    .ZN(_11876_));
 BUF_X4 _34477_ (.A(_11876_),
    .Z(_11877_));
 BUF_X4 _34478_ (.A(_11877_),
    .Z(_11878_));
 MUX2_X1 _34479_ (.A(\core.keymem.key_mem[0][100] ),
    .B(_11873_),
    .S(_11878_),
    .Z(_00838_));
 INV_X2 _34480_ (.A(_00129_),
    .ZN(_11879_));
 CLKBUF_X3 _34481_ (.A(_11877_),
    .Z(_11880_));
 NAND3_X1 _34482_ (.A1(_16286_),
    .A2(_11879_),
    .A3(_11880_),
    .ZN(_11881_));
 BUF_X4 _34483_ (.A(_11877_),
    .Z(_11882_));
 CLKBUF_X3 _34484_ (.A(_11882_),
    .Z(_11883_));
 INV_X1 _34485_ (.A(\core.keymem.key_mem[0][101] ),
    .ZN(_11884_));
 OAI21_X1 _34486_ (.A(_11881_),
    .B1(_11883_),
    .B2(_11884_),
    .ZN(_00839_));
 BUF_X4 _34487_ (.A(_11874_),
    .Z(_11885_));
 NOR2_X1 _34488_ (.A1(_00130_),
    .A2(_11885_),
    .ZN(_11886_));
 XNOR2_X2 _34489_ (.A(\core.keymem.prev_key1_reg[102] ),
    .B(_10221_),
    .ZN(_11887_));
 NOR2_X4 _34490_ (.A1(_16219_),
    .A2(_11840_),
    .ZN(_11888_));
 BUF_X8 _34491_ (.A(_11888_),
    .Z(_11889_));
 AOI21_X2 _34492_ (.A(_11886_),
    .B1(_11887_),
    .B2(_11889_),
    .ZN(_11890_));
 BUF_X4 _34493_ (.A(_11818_),
    .Z(_11891_));
 BUF_X4 _34494_ (.A(_11891_),
    .Z(_11892_));
 AND2_X1 _34495_ (.A1(\core.key[102] ),
    .A2(_11892_),
    .ZN(_11893_));
 BUF_X2 _34496_ (.A(\core.keymem.prev_key0_reg[102] ),
    .Z(_11894_));
 OR4_X4 _34497_ (.A1(_11856_),
    .A2(_07044_),
    .A3(_08916_),
    .A4(_10525_),
    .ZN(_11895_));
 AND4_X1 _34498_ (.A1(_10194_),
    .A2(_10198_),
    .A3(_10204_),
    .A4(_10219_),
    .ZN(_11896_));
 NAND3_X2 _34499_ (.A1(_11851_),
    .A2(_09708_),
    .A3(_11896_),
    .ZN(_11897_));
 NAND2_X1 _34500_ (.A1(_11895_),
    .A2(_11897_),
    .ZN(_11898_));
 XNOR2_X2 _34501_ (.A(_11894_),
    .B(_11898_),
    .ZN(_11899_));
 BUF_X8 _34502_ (.A(_11827_),
    .Z(_11900_));
 BUF_X8 _34503_ (.A(_11900_),
    .Z(_11901_));
 AOI21_X2 _34504_ (.A(_11893_),
    .B1(_11899_),
    .B2(_11901_),
    .ZN(_11902_));
 NAND2_X4 _34505_ (.A1(_16219_),
    .A2(_11813_),
    .ZN(_11903_));
 BUF_X4 _34506_ (.A(_11903_),
    .Z(_11904_));
 OAI21_X4 _34507_ (.A(_11890_),
    .B1(_11902_),
    .B2(_11904_),
    .ZN(_11905_));
 BUF_X2 _34508_ (.A(_11905_),
    .Z(_11906_));
 AOI22_X1 _34509_ (.A1(\core.keymem.key_mem[0][102] ),
    .A2(_11802_),
    .B1(_11806_),
    .B2(_11906_),
    .ZN(_11907_));
 INV_X1 _34510_ (.A(_11907_),
    .ZN(_00840_));
 BUF_X4 _34511_ (.A(_16219_),
    .Z(_11908_));
 BUF_X4 _34512_ (.A(_11908_),
    .Z(_11909_));
 OR2_X2 _34513_ (.A1(_10253_),
    .A2(_10259_),
    .ZN(_11910_));
 XNOR2_X1 _34514_ (.A(_00132_),
    .B(_11910_),
    .ZN(_11911_));
 NOR2_X1 _34515_ (.A1(_11798_),
    .A2(_11911_),
    .ZN(_11912_));
 AOI21_X2 _34516_ (.A(_11912_),
    .B1(_11841_),
    .B2(_00131_),
    .ZN(_11913_));
 OAI21_X2 _34517_ (.A(_16228_),
    .B1(_11909_),
    .B2(_11913_),
    .ZN(_11914_));
 OR2_X1 _34518_ (.A1(_00131_),
    .A2(_11885_),
    .ZN(_11915_));
 BUF_X8 _34519_ (.A(_11811_),
    .Z(_11916_));
 BUF_X8 _34520_ (.A(_11874_),
    .Z(_11917_));
 CLKBUF_X2 _34521_ (.A(\core.keymem.prev_key0_reg[103] ),
    .Z(_11918_));
 INV_X1 _34522_ (.A(_11918_),
    .ZN(_11919_));
 BUF_X8 _34523_ (.A(_11851_),
    .Z(_11920_));
 NOR2_X2 _34524_ (.A1(_11920_),
    .A2(_10565_),
    .ZN(_11921_));
 NOR3_X2 _34525_ (.A1(_11832_),
    .A2(_10253_),
    .A3(_10259_),
    .ZN(_11922_));
 NOR2_X1 _34526_ (.A1(_11921_),
    .A2(_11922_),
    .ZN(_11923_));
 XNOR2_X2 _34527_ (.A(_11919_),
    .B(_11923_),
    .ZN(_11924_));
 BUF_X4 _34528_ (.A(_11826_),
    .Z(_11925_));
 MUX2_X1 _34529_ (.A(\core.key[103] ),
    .B(_11924_),
    .S(_11925_),
    .Z(_11926_));
 AOI21_X2 _34530_ (.A(_11916_),
    .B1(_11917_),
    .B2(_11926_),
    .ZN(_11927_));
 AOI21_X4 _34531_ (.A(_11914_),
    .B1(_11915_),
    .B2(_11927_),
    .ZN(_11928_));
 BUF_X2 _34532_ (.A(_11928_),
    .Z(_11929_));
 MUX2_X1 _34533_ (.A(\core.keymem.key_mem[0][103] ),
    .B(_11929_),
    .S(_11878_),
    .Z(_00841_));
 BUF_X4 _34534_ (.A(_11805_),
    .Z(_11930_));
 NOR2_X1 _34535_ (.A1(_11930_),
    .A2(_00133_),
    .ZN(_11931_));
 MUX2_X1 _34536_ (.A(\core.keymem.key_mem[0][104] ),
    .B(_11931_),
    .S(_11878_),
    .Z(_00842_));
 NOR2_X1 _34537_ (.A1(_11930_),
    .A2(_00134_),
    .ZN(_11932_));
 MUX2_X1 _34538_ (.A(\core.keymem.key_mem[0][105] ),
    .B(_11932_),
    .S(_11878_),
    .Z(_00843_));
 BUF_X4 _34539_ (.A(_11801_),
    .Z(_11933_));
 NAND2_X1 _34540_ (.A1(\core.keymem.key_mem[0][106] ),
    .A2(_11933_),
    .ZN(_11934_));
 OR2_X4 _34541_ (.A1(_00135_),
    .A2(_11868_),
    .ZN(_11935_));
 BUF_X8 _34542_ (.A(_11823_),
    .Z(_11936_));
 BUF_X2 _34543_ (.A(\core.keymem.prev_key0_reg[106] ),
    .Z(_11937_));
 OR3_X2 _34544_ (.A1(_11857_),
    .A2(_07613_),
    .A3(_07641_),
    .ZN(_11938_));
 NOR4_X4 _34545_ (.A1(_10116_),
    .A2(_10133_),
    .A3(_10140_),
    .A4(_10156_),
    .ZN(_11939_));
 NAND2_X1 _34546_ (.A1(_07062_),
    .A2(_10322_),
    .ZN(_11940_));
 OAI21_X4 _34547_ (.A(_11940_),
    .B1(_10166_),
    .B2(_07062_),
    .ZN(_11941_));
 NAND3_X2 _34548_ (.A1(_11920_),
    .A2(_11939_),
    .A3(_11941_),
    .ZN(_11942_));
 NAND2_X1 _34549_ (.A1(_11938_),
    .A2(_11942_),
    .ZN(_11943_));
 XNOR2_X2 _34550_ (.A(_11937_),
    .B(_11943_),
    .ZN(_11944_));
 BUF_X4 _34551_ (.A(_11848_),
    .Z(_11945_));
 MUX2_X1 _34552_ (.A(\core.key[106] ),
    .B(_11944_),
    .S(_11945_),
    .Z(_11946_));
 NOR2_X4 _34553_ (.A1(_10157_),
    .A2(_10167_),
    .ZN(_11947_));
 XNOR2_X1 _34554_ (.A(_00136_),
    .B(_11947_),
    .ZN(_11948_));
 OAI21_X2 _34555_ (.A(_11935_),
    .B1(_11948_),
    .B2(_11841_),
    .ZN(_11949_));
 AOI22_X4 _34556_ (.A1(_11936_),
    .A2(_11946_),
    .B1(_11949_),
    .B2(_11866_),
    .ZN(_11950_));
 AND2_X1 _34557_ (.A1(_11935_),
    .A2(_11950_),
    .ZN(_11951_));
 BUF_X4 _34558_ (.A(_16229_),
    .Z(_11952_));
 NAND2_X2 _34559_ (.A1(_11952_),
    .A2(_11876_),
    .ZN(_11953_));
 BUF_X4 _34560_ (.A(_11953_),
    .Z(_11954_));
 OAI21_X1 _34561_ (.A(_11934_),
    .B1(_11951_),
    .B2(_11954_),
    .ZN(_00844_));
 NAND2_X1 _34562_ (.A1(_00137_),
    .A2(_11798_),
    .ZN(_11955_));
 XNOR2_X1 _34563_ (.A(_00138_),
    .B(_10352_),
    .ZN(_11956_));
 NAND2_X1 _34564_ (.A1(_11862_),
    .A2(_11956_),
    .ZN(_11957_));
 AOI21_X2 _34565_ (.A(_11908_),
    .B1(_11955_),
    .B2(_11957_),
    .ZN(_11958_));
 OR2_X1 _34566_ (.A1(_00137_),
    .A2(_11874_),
    .ZN(_11959_));
 BUF_X8 _34567_ (.A(_11868_),
    .Z(_11960_));
 NOR2_X4 _34568_ (.A1(_07753_),
    .A2(_07785_),
    .ZN(_11961_));
 MUX2_X2 _34569_ (.A(_11961_),
    .B(_10352_),
    .S(_11857_),
    .Z(_11962_));
 XNOR2_X1 _34570_ (.A(\core.keymem.prev_key0_reg[107] ),
    .B(_11962_),
    .ZN(_11963_));
 MUX2_X1 _34571_ (.A(\core.key[107] ),
    .B(_11963_),
    .S(_11860_),
    .Z(_11964_));
 AOI21_X2 _34572_ (.A(_11846_),
    .B1(_11960_),
    .B2(_11964_),
    .ZN(_11965_));
 AOI211_X2 _34573_ (.A(_11804_),
    .B(_11958_),
    .C1(_11959_),
    .C2(_11965_),
    .ZN(_11966_));
 BUF_X2 _34574_ (.A(_11966_),
    .Z(_11967_));
 MUX2_X1 _34575_ (.A(\core.keymem.key_mem[0][107] ),
    .B(_11967_),
    .S(_11878_),
    .Z(_00845_));
 NAND2_X1 _34576_ (.A1(\core.key[108] ),
    .A2(_11819_),
    .ZN(_11968_));
 BUF_X2 _34577_ (.A(\core.keymem.prev_key0_reg[108] ),
    .Z(_11969_));
 INV_X1 _34578_ (.A(_11969_),
    .ZN(_11970_));
 NOR3_X2 _34579_ (.A1(_11856_),
    .A2(_07828_),
    .A3(_07891_),
    .ZN(_11971_));
 NOR2_X1 _34580_ (.A1(_11831_),
    .A2(_10413_),
    .ZN(_11972_));
 OR2_X2 _34581_ (.A1(_11971_),
    .A2(_11972_),
    .ZN(_11973_));
 XNOR2_X2 _34582_ (.A(_11970_),
    .B(_11973_),
    .ZN(_11974_));
 OAI21_X1 _34583_ (.A(_11968_),
    .B1(_11974_),
    .B2(_11891_),
    .ZN(_11975_));
 AOI21_X2 _34584_ (.A(_11846_),
    .B1(_11874_),
    .B2(_11975_),
    .ZN(_11976_));
 OR2_X1 _34585_ (.A1(_00139_),
    .A2(_11868_),
    .ZN(_11977_));
 XOR2_X1 _34586_ (.A(_00140_),
    .B(_10413_),
    .Z(_11978_));
 MUX2_X1 _34587_ (.A(_00139_),
    .B(_11978_),
    .S(_11862_),
    .Z(_11979_));
 AOI221_X2 _34588_ (.A(_11804_),
    .B1(_11976_),
    .B2(_11977_),
    .C1(_11979_),
    .C2(_11866_),
    .ZN(_11980_));
 CLKBUF_X2 _34589_ (.A(_11980_),
    .Z(_11981_));
 MUX2_X1 _34590_ (.A(\core.keymem.key_mem[0][108] ),
    .B(_11981_),
    .S(_11878_),
    .Z(_00846_));
 NOR2_X1 _34591_ (.A1(_11930_),
    .A2(_00141_),
    .ZN(_11982_));
 MUX2_X1 _34592_ (.A(\core.keymem.key_mem[0][109] ),
    .B(_11982_),
    .S(_11878_),
    .Z(_00847_));
 CLKBUF_X3 _34593_ (.A(_00405_),
    .Z(_11983_));
 NOR2_X1 _34594_ (.A1(_11930_),
    .A2(_11983_),
    .ZN(_11984_));
 MUX2_X1 _34595_ (.A(\core.keymem.key_mem[0][10] ),
    .B(_11984_),
    .S(_11878_),
    .Z(_00848_));
 NAND2_X1 _34596_ (.A1(\core.keymem.key_mem[0][110] ),
    .A2(_11933_),
    .ZN(_11985_));
 BUF_X4 _34597_ (.A(_11952_),
    .Z(_11986_));
 BUF_X4 _34598_ (.A(_11903_),
    .Z(_11987_));
 BUF_X4 _34599_ (.A(_11819_),
    .Z(_11988_));
 BUF_X8 _34600_ (.A(_11988_),
    .Z(_11989_));
 INV_X1 _34601_ (.A(\core.key[110] ),
    .ZN(_11990_));
 AOI21_X1 _34602_ (.A(_11987_),
    .B1(_11989_),
    .B2(_11990_),
    .ZN(_11991_));
 BUF_X2 _34603_ (.A(\core.keymem.prev_key0_reg[110] ),
    .Z(_11992_));
 AOI21_X1 _34604_ (.A(_11829_),
    .B1(_10466_),
    .B2(_10463_),
    .ZN(_11993_));
 NAND4_X2 _34605_ (.A1(_10494_),
    .A2(_10505_),
    .A3(_10524_),
    .A4(_11993_),
    .ZN(_11994_));
 OAI33_X1 _34606_ (.A1(_11850_),
    .A2(_07974_),
    .A3(_08100_),
    .B1(_08916_),
    .B2(_11994_),
    .B3(_07044_),
    .ZN(_11995_));
 XNOR2_X2 _34607_ (.A(_11992_),
    .B(net11),
    .ZN(_11996_));
 BUF_X8 _34608_ (.A(_11892_),
    .Z(_11997_));
 OAI21_X2 _34609_ (.A(_11991_),
    .B1(_11996_),
    .B2(_11997_),
    .ZN(_11998_));
 CLKBUF_X2 _34610_ (.A(\core.keymem.prev_key1_reg[110] ),
    .Z(_11999_));
 XOR2_X2 _34611_ (.A(_11999_),
    .B(_10526_),
    .Z(_12000_));
 BUF_X4 _34612_ (.A(_11814_),
    .Z(_12001_));
 BUF_X4 _34613_ (.A(_11885_),
    .Z(_12002_));
 OAI221_X2 _34614_ (.A(_11998_),
    .B1(_12000_),
    .B2(_12001_),
    .C1(_12002_),
    .C2(_00142_),
    .ZN(_12003_));
 NAND2_X1 _34615_ (.A1(_11986_),
    .A2(_12003_),
    .ZN(_12004_));
 BUF_X8 _34616_ (.A(_11801_),
    .Z(_12005_));
 OAI21_X1 _34617_ (.A(_11985_),
    .B1(_12004_),
    .B2(_12005_),
    .ZN(_00849_));
 NAND2_X1 _34618_ (.A1(_00143_),
    .A2(_11798_),
    .ZN(_12006_));
 XOR2_X1 _34619_ (.A(_00144_),
    .B(_10565_),
    .Z(_12007_));
 NAND2_X1 _34620_ (.A1(_11868_),
    .A2(_12007_),
    .ZN(_12008_));
 AOI21_X1 _34621_ (.A(_06676_),
    .B1(_12006_),
    .B2(_12008_),
    .ZN(_12009_));
 OR2_X1 _34622_ (.A1(_11804_),
    .A2(_12009_),
    .ZN(_12010_));
 OR2_X1 _34623_ (.A1(_00143_),
    .A2(_11885_),
    .ZN(_12011_));
 MUX2_X1 _34624_ (.A(_08163_),
    .B(_10565_),
    .S(_11850_),
    .Z(_12012_));
 XOR2_X2 _34625_ (.A(\core.keymem.prev_key0_reg[111] ),
    .B(_12012_),
    .Z(_12013_));
 MUX2_X1 _34626_ (.A(\core.key[111] ),
    .B(_12013_),
    .S(_11925_),
    .Z(_12014_));
 AOI21_X2 _34627_ (.A(_11916_),
    .B1(_11917_),
    .B2(_12014_),
    .ZN(_12015_));
 AOI21_X4 _34628_ (.A(_12010_),
    .B1(_12011_),
    .B2(_12015_),
    .ZN(_12016_));
 BUF_X2 _34629_ (.A(_12016_),
    .Z(_12017_));
 BUF_X4 _34630_ (.A(_11877_),
    .Z(_12018_));
 MUX2_X1 _34631_ (.A(\core.keymem.key_mem[0][111] ),
    .B(_12017_),
    .S(_12018_),
    .Z(_00850_));
 NAND4_X2 _34632_ (.A1(_11856_),
    .A2(_10592_),
    .A3(_10605_),
    .A4(_10611_),
    .ZN(_12019_));
 OAI33_X1 _34633_ (.A1(_11857_),
    .A2(_08483_),
    .A3(_08596_),
    .B1(_12019_),
    .B2(_07982_),
    .B3(_07974_),
    .ZN(_12020_));
 XNOR2_X2 _34634_ (.A(\core.keymem.prev_key0_reg[112] ),
    .B(net13),
    .ZN(_12021_));
 MUX2_X1 _34635_ (.A(\core.key[112] ),
    .B(_12021_),
    .S(_11828_),
    .Z(_12022_));
 NAND2_X1 _34636_ (.A1(_11936_),
    .A2(_12022_),
    .ZN(_12023_));
 NOR2_X1 _34637_ (.A1(_00145_),
    .A2(_11863_),
    .ZN(_12024_));
 BUF_X2 _34638_ (.A(\core.keymem.prev_key1_reg[112] ),
    .Z(_12025_));
 XNOR2_X2 _34639_ (.A(_12025_),
    .B(_10613_),
    .ZN(_12026_));
 BUF_X8 _34640_ (.A(_11888_),
    .Z(_12027_));
 BUF_X8 _34641_ (.A(_12027_),
    .Z(_12028_));
 AOI21_X2 _34642_ (.A(_12024_),
    .B1(_12026_),
    .B2(_12028_),
    .ZN(_12029_));
 NAND2_X4 _34643_ (.A1(_12023_),
    .A2(_12029_),
    .ZN(_12030_));
 BUF_X2 _34644_ (.A(_12030_),
    .Z(_12031_));
 AOI22_X1 _34645_ (.A1(\core.keymem.key_mem[0][112] ),
    .A2(_11802_),
    .B1(_11806_),
    .B2(_12031_),
    .ZN(_12032_));
 INV_X1 _34646_ (.A(_12032_),
    .ZN(_00851_));
 NOR2_X1 _34647_ (.A1(_11930_),
    .A2(_00146_),
    .ZN(_12033_));
 MUX2_X1 _34648_ (.A(\core.keymem.key_mem[0][113] ),
    .B(_12033_),
    .S(_12018_),
    .Z(_00852_));
 NAND2_X1 _34649_ (.A1(\core.keymem.key_mem[0][114] ),
    .A2(_11933_),
    .ZN(_12034_));
 BUF_X8 _34650_ (.A(_11960_),
    .Z(_12035_));
 INV_X1 _34651_ (.A(\core.key[114] ),
    .ZN(_12036_));
 CLKBUF_X3 _34652_ (.A(\core.keymem.prev_key0_reg[114] ),
    .Z(_12037_));
 INV_X2 _34653_ (.A(_12037_),
    .ZN(_12038_));
 AND2_X1 _34654_ (.A1(_11831_),
    .A2(_08803_),
    .ZN(_12039_));
 BUF_X4 _34655_ (.A(_11830_),
    .Z(_12040_));
 NOR3_X4 _34656_ (.A1(_12040_),
    .A2(_07613_),
    .A3(_07641_),
    .ZN(_12041_));
 OR2_X2 _34657_ (.A1(_12039_),
    .A2(_12041_),
    .ZN(_12042_));
 XNOR2_X2 _34658_ (.A(_12038_),
    .B(_12042_),
    .ZN(_12043_));
 BUF_X4 _34659_ (.A(_11848_),
    .Z(_12044_));
 MUX2_X1 _34660_ (.A(_12036_),
    .B(_12043_),
    .S(_12044_),
    .Z(_12045_));
 NOR2_X4 _34661_ (.A1(_07613_),
    .A2(_07641_),
    .ZN(_12046_));
 XNOR2_X1 _34662_ (.A(_00148_),
    .B(_12046_),
    .ZN(_12047_));
 OAI222_X2 _34663_ (.A1(_00147_),
    .A2(_12035_),
    .B1(_11904_),
    .B2(_12045_),
    .C1(_12047_),
    .C2(_12001_),
    .ZN(_12048_));
 NAND2_X1 _34664_ (.A1(_16285_),
    .A2(_12048_),
    .ZN(_12049_));
 OAI21_X1 _34665_ (.A(_12034_),
    .B1(_12049_),
    .B2(_12005_),
    .ZN(_00853_));
 NAND2_X1 _34666_ (.A1(\core.key[115] ),
    .A2(_11819_),
    .ZN(_12050_));
 MUX2_X1 _34667_ (.A(_11961_),
    .B(_08886_),
    .S(_11831_),
    .Z(_12051_));
 XOR2_X2 _34668_ (.A(\core.keymem.prev_key0_reg[115] ),
    .B(_12051_),
    .Z(_12052_));
 OAI21_X1 _34669_ (.A(_12050_),
    .B1(_12052_),
    .B2(_11891_),
    .ZN(_12053_));
 AOI21_X2 _34670_ (.A(_11811_),
    .B1(_11874_),
    .B2(_12053_),
    .ZN(_12054_));
 OR2_X1 _34671_ (.A1(_00149_),
    .A2(_11868_),
    .ZN(_12055_));
 XNOR2_X1 _34672_ (.A(_00150_),
    .B(_11961_),
    .ZN(_12056_));
 MUX2_X1 _34673_ (.A(_00149_),
    .B(_12056_),
    .S(_11862_),
    .Z(_12057_));
 AOI221_X2 _34674_ (.A(_11804_),
    .B1(_12054_),
    .B2(_12055_),
    .C1(_12057_),
    .C2(_11866_),
    .ZN(_12058_));
 CLKBUF_X2 _34675_ (.A(_12058_),
    .Z(_12059_));
 MUX2_X1 _34676_ (.A(\core.keymem.key_mem[0][115] ),
    .B(_12059_),
    .S(_12018_),
    .Z(_00854_));
 NAND2_X1 _34677_ (.A1(\core.key[116] ),
    .A2(_11819_),
    .ZN(_12060_));
 CLKBUF_X2 _34678_ (.A(\core.keymem.prev_key0_reg[116] ),
    .Z(_12061_));
 INV_X1 _34679_ (.A(_12061_),
    .ZN(_12062_));
 BUF_X4 _34680_ (.A(_11829_),
    .Z(_12063_));
 NOR3_X4 _34681_ (.A1(_08836_),
    .A2(_09019_),
    .A3(_09026_),
    .ZN(_12064_));
 NOR4_X4 _34682_ (.A1(_09030_),
    .A2(_09038_),
    .A3(_09048_),
    .A4(_09057_),
    .ZN(_12065_));
 NAND3_X2 _34683_ (.A1(_12063_),
    .A2(_12064_),
    .A3(_12065_),
    .ZN(_12066_));
 OR3_X2 _34684_ (.A1(_11829_),
    .A2(_07828_),
    .A3(_07891_),
    .ZN(_12067_));
 NAND2_X1 _34685_ (.A1(_12066_),
    .A2(_12067_),
    .ZN(_12068_));
 XNOR2_X2 _34686_ (.A(_12062_),
    .B(_12068_),
    .ZN(_12069_));
 OAI21_X1 _34687_ (.A(_12060_),
    .B1(_12069_),
    .B2(_11891_),
    .ZN(_12070_));
 AOI21_X2 _34688_ (.A(_11811_),
    .B1(_11874_),
    .B2(_12070_),
    .ZN(_12071_));
 OR2_X1 _34689_ (.A1(_00151_),
    .A2(_11868_),
    .ZN(_12072_));
 NOR2_X2 _34690_ (.A1(_07828_),
    .A2(_07891_),
    .ZN(_12073_));
 XNOR2_X1 _34691_ (.A(_00152_),
    .B(_12073_),
    .ZN(_12074_));
 MUX2_X1 _34692_ (.A(_00151_),
    .B(_12074_),
    .S(_11862_),
    .Z(_12075_));
 AOI221_X2 _34693_ (.A(_11804_),
    .B1(_12071_),
    .B2(_12072_),
    .C1(_12075_),
    .C2(_11866_),
    .ZN(_12076_));
 CLKBUF_X2 _34694_ (.A(_12076_),
    .Z(_12077_));
 MUX2_X1 _34695_ (.A(\core.keymem.key_mem[0][116] ),
    .B(_12077_),
    .S(_12018_),
    .Z(_00855_));
 NOR2_X1 _34696_ (.A1(_11930_),
    .A2(_00153_),
    .ZN(_12078_));
 MUX2_X1 _34697_ (.A(\core.keymem.key_mem[0][117] ),
    .B(_12078_),
    .S(_12018_),
    .Z(_00856_));
 INV_X1 _34698_ (.A(_00154_),
    .ZN(_12079_));
 NAND3_X1 _34699_ (.A1(_16286_),
    .A2(_12079_),
    .A3(_11880_),
    .ZN(_12080_));
 INV_X1 _34700_ (.A(\core.keymem.key_mem[0][118] ),
    .ZN(_12081_));
 OAI21_X1 _34701_ (.A(_12080_),
    .B1(_11883_),
    .B2(_12081_),
    .ZN(_00857_));
 NAND2_X1 _34702_ (.A1(_00155_),
    .A2(_11840_),
    .ZN(_12082_));
 XOR2_X1 _34703_ (.A(_00156_),
    .B(_08163_),
    .Z(_12083_));
 NAND2_X1 _34704_ (.A1(_11868_),
    .A2(_12083_),
    .ZN(_12084_));
 AOI21_X1 _34705_ (.A(_06676_),
    .B1(_12082_),
    .B2(_12084_),
    .ZN(_12085_));
 OR2_X1 _34706_ (.A1(_11804_),
    .A2(_12085_),
    .ZN(_12086_));
 OR2_X1 _34707_ (.A1(_00155_),
    .A2(_11885_),
    .ZN(_12087_));
 NAND2_X1 _34708_ (.A1(\core.key[119] ),
    .A2(_11988_),
    .ZN(_12088_));
 CLKBUF_X3 _34709_ (.A(\core.keymem.prev_key0_reg[119] ),
    .Z(_12089_));
 MUX2_X2 _34710_ (.A(_08163_),
    .B(_09209_),
    .S(_12063_),
    .Z(_12090_));
 XNOR2_X2 _34711_ (.A(_12089_),
    .B(_12090_),
    .ZN(_12091_));
 BUF_X4 _34712_ (.A(_11820_),
    .Z(_12092_));
 OAI21_X2 _34713_ (.A(_12088_),
    .B1(_12091_),
    .B2(_12092_),
    .ZN(_12093_));
 AOI21_X4 _34714_ (.A(_11916_),
    .B1(_11917_),
    .B2(_12093_),
    .ZN(_12094_));
 AOI21_X4 _34715_ (.A(_12086_),
    .B1(_12087_),
    .B2(_12094_),
    .ZN(_12095_));
 CLKBUF_X2 _34716_ (.A(_12095_),
    .Z(_12096_));
 MUX2_X1 _34717_ (.A(\core.keymem.key_mem[0][119] ),
    .B(_12096_),
    .S(_12018_),
    .Z(_00858_));
 NOR2_X1 _34718_ (.A1(_11930_),
    .A2(_00406_),
    .ZN(_12097_));
 MUX2_X1 _34719_ (.A(\core.keymem.key_mem[0][11] ),
    .B(_12097_),
    .S(_12018_),
    .Z(_00859_));
 BUF_X4 _34720_ (.A(_11823_),
    .Z(_12098_));
 BUF_X4 _34721_ (.A(_12044_),
    .Z(_12099_));
 NOR2_X1 _34722_ (.A1(_00158_),
    .A2(_12099_),
    .ZN(_12100_));
 BUF_X4 _34723_ (.A(_11820_),
    .Z(_12101_));
 INV_X1 _34724_ (.A(\core.keymem.prev_key0_reg[120] ),
    .ZN(_12102_));
 NOR2_X1 _34725_ (.A1(_11857_),
    .A2(_12102_),
    .ZN(_12103_));
 OAI21_X1 _34726_ (.A(_12103_),
    .B1(_09680_),
    .B2(_09569_),
    .ZN(_12104_));
 OR4_X1 _34727_ (.A1(_11851_),
    .A2(\core.keymem.prev_key0_reg[120] ),
    .A3(_09569_),
    .A4(_09680_),
    .ZN(_12105_));
 BUF_X2 _34728_ (.A(\core.keymem.rcon_reg[0] ),
    .Z(_12106_));
 AND3_X1 _34729_ (.A1(_11856_),
    .A2(_12106_),
    .A3(_12102_),
    .ZN(_12107_));
 NOR3_X1 _34730_ (.A1(_11831_),
    .A2(_12106_),
    .A3(_12102_),
    .ZN(_12108_));
 OAI22_X2 _34731_ (.A1(_08483_),
    .A2(_08596_),
    .B1(_12107_),
    .B2(_12108_),
    .ZN(_12109_));
 INV_X1 _34732_ (.A(_08314_),
    .ZN(_12110_));
 AND4_X2 _34733_ (.A1(_08353_),
    .A2(_08376_),
    .A3(_08404_),
    .A4(_08437_),
    .ZN(_12111_));
 AND4_X2 _34734_ (.A1(_08446_),
    .A2(_08458_),
    .A3(_08468_),
    .A4(_08481_),
    .ZN(_12112_));
 AOI21_X2 _34735_ (.A(_12110_),
    .B1(_12111_),
    .B2(_12112_),
    .ZN(_12113_));
 NOR4_X4 _34736_ (.A1(_08495_),
    .A2(_08527_),
    .A3(_08560_),
    .A4(_08595_),
    .ZN(_12114_));
 NOR3_X1 _34737_ (.A1(_11831_),
    .A2(_12106_),
    .A3(\core.keymem.prev_key0_reg[120] ),
    .ZN(_12115_));
 AND3_X1 _34738_ (.A1(_11856_),
    .A2(_12106_),
    .A3(\core.keymem.prev_key0_reg[120] ),
    .ZN(_12116_));
 OAI211_X2 _34739_ (.A(_12113_),
    .B(_12114_),
    .C1(_12115_),
    .C2(_12116_),
    .ZN(_12117_));
 NAND4_X4 _34740_ (.A1(_12104_),
    .A2(_12105_),
    .A3(_12109_),
    .A4(_12117_),
    .ZN(_12118_));
 NOR2_X1 _34741_ (.A1(_12101_),
    .A2(_12118_),
    .ZN(_12119_));
 OAI21_X1 _34742_ (.A(_12098_),
    .B1(_12100_),
    .B2(_12119_),
    .ZN(_12120_));
 XNOR2_X2 _34743_ (.A(_12106_),
    .B(_08597_),
    .ZN(_12121_));
 XNOR2_X2 _34744_ (.A(\core.keymem.prev_key1_reg[120] ),
    .B(_12121_),
    .ZN(_12122_));
 OAI221_X2 _34745_ (.A(_12120_),
    .B1(_12122_),
    .B2(_12001_),
    .C1(_12035_),
    .C2(_00157_),
    .ZN(_12123_));
 BUF_X2 _34746_ (.A(_12123_),
    .Z(_12124_));
 AOI22_X1 _34747_ (.A1(\core.keymem.key_mem[0][120] ),
    .A2(_11802_),
    .B1(_11806_),
    .B2(_12124_),
    .ZN(_12125_));
 INV_X1 _34748_ (.A(_12125_),
    .ZN(_00860_));
 BUF_X1 _34749_ (.A(\core.keymem.prev_key0_reg[121] ),
    .Z(_12126_));
 INV_X1 _34750_ (.A(_12126_),
    .ZN(_12127_));
 NOR2_X1 _34751_ (.A1(_11920_),
    .A2(_12127_),
    .ZN(_12128_));
 NAND3_X1 _34752_ (.A1(_09734_),
    .A2(_09753_),
    .A3(_09775_),
    .ZN(_12129_));
 OAI21_X2 _34753_ (.A(_12128_),
    .B1(_12129_),
    .B2(_10179_),
    .ZN(_12130_));
 NAND4_X2 _34754_ (.A1(_11832_),
    .A2(_12127_),
    .A3(_09708_),
    .A4(_09776_),
    .ZN(_12131_));
 BUF_X2 _34755_ (.A(\core.keymem.rcon_logic.tmp_rcon[2] ),
    .Z(_12132_));
 NAND2_X1 _34756_ (.A1(_11850_),
    .A2(_12132_),
    .ZN(_12133_));
 NOR2_X1 _34757_ (.A1(_12126_),
    .A2(_12133_),
    .ZN(_12134_));
 NOR2_X1 _34758_ (.A1(_12063_),
    .A2(_12132_),
    .ZN(_12135_));
 AND2_X1 _34759_ (.A1(_12126_),
    .A2(_12135_),
    .ZN(_12136_));
 OAI21_X2 _34760_ (.A(_08705_),
    .B1(_12134_),
    .B2(_12136_),
    .ZN(_12137_));
 NOR2_X2 _34761_ (.A1(_08653_),
    .A2(_08704_),
    .ZN(_12138_));
 NAND2_X1 _34762_ (.A1(_08708_),
    .A2(_08713_),
    .ZN(_12139_));
 AOI21_X4 _34763_ (.A(_12139_),
    .B1(_12111_),
    .B2(_12112_),
    .ZN(_12140_));
 NAND4_X2 _34764_ (.A1(_12127_),
    .A2(_12138_),
    .A3(_12140_),
    .A4(_12135_),
    .ZN(_12141_));
 NAND4_X4 _34765_ (.A1(_12130_),
    .A2(_12131_),
    .A3(_12137_),
    .A4(_12141_),
    .ZN(_12142_));
 OR4_X1 _34766_ (.A1(_12127_),
    .A2(_08705_),
    .A3(_08715_),
    .A4(_12133_),
    .ZN(_12143_));
 NAND2_X1 _34767_ (.A1(_08715_),
    .A2(_12134_),
    .ZN(_12144_));
 NAND2_X1 _34768_ (.A1(_08715_),
    .A2(_12136_),
    .ZN(_12145_));
 NAND3_X2 _34769_ (.A1(_12143_),
    .A2(_12144_),
    .A3(_12145_),
    .ZN(_12146_));
 NOR3_X2 _34770_ (.A1(_12092_),
    .A2(_12142_),
    .A3(_12146_),
    .ZN(_12147_));
 BUF_X4 _34771_ (.A(_06676_),
    .Z(_12148_));
 BUF_X4 _34772_ (.A(_12044_),
    .Z(_12149_));
 OAI21_X1 _34773_ (.A(_12148_),
    .B1(_00160_),
    .B2(_12149_),
    .ZN(_12150_));
 INV_X1 _34774_ (.A(_12132_),
    .ZN(_12151_));
 AOI21_X2 _34775_ (.A(_12151_),
    .B1(_12138_),
    .B2(_12140_),
    .ZN(_12152_));
 NOR3_X2 _34776_ (.A1(_12132_),
    .A2(_08705_),
    .A3(_08715_),
    .ZN(_12153_));
 NOR2_X2 _34777_ (.A1(_12152_),
    .A2(_12153_),
    .ZN(_12154_));
 XOR2_X2 _34778_ (.A(\core.keymem.prev_key1_reg[121] ),
    .B(_12154_),
    .Z(_12155_));
 BUF_X4 _34779_ (.A(_11908_),
    .Z(_12156_));
 OAI221_X2 _34780_ (.A(_12035_),
    .B1(_12147_),
    .B2(_12150_),
    .C1(_12155_),
    .C2(_12156_),
    .ZN(_12157_));
 BUF_X4 _34781_ (.A(_11917_),
    .Z(_12158_));
 OAI21_X4 _34782_ (.A(_12157_),
    .B1(_12158_),
    .B2(_00159_),
    .ZN(_12159_));
 BUF_X2 _34783_ (.A(_12159_),
    .Z(_12160_));
 AOI22_X1 _34784_ (.A1(\core.keymem.key_mem[0][121] ),
    .A2(_11802_),
    .B1(_11806_),
    .B2(_12160_),
    .ZN(_12161_));
 INV_X1 _34785_ (.A(_12161_),
    .ZN(_00861_));
 INV_X2 _34786_ (.A(_00161_),
    .ZN(_12162_));
 NAND3_X1 _34787_ (.A1(_16286_),
    .A2(_12162_),
    .A3(_11880_),
    .ZN(_12163_));
 INV_X1 _34788_ (.A(\core.keymem.key_mem[0][122] ),
    .ZN(_12164_));
 OAI21_X1 _34789_ (.A(_12163_),
    .B1(_11883_),
    .B2(_12164_),
    .ZN(_00862_));
 NAND2_X1 _34790_ (.A1(\core.keymem.key_mem[0][123] ),
    .A2(_11933_),
    .ZN(_12165_));
 CLKBUF_X3 _34791_ (.A(\core.keymem.rcon_reg[3] ),
    .Z(_12166_));
 XNOR2_X2 _34792_ (.A(_12166_),
    .B(_08886_),
    .ZN(_12167_));
 XNOR2_X2 _34793_ (.A(\core.keymem.prev_key1_reg[123] ),
    .B(_12167_),
    .ZN(_12168_));
 AOI22_X2 _34794_ (.A1(_00163_),
    .A2(_11800_),
    .B1(_11889_),
    .B2(_12168_),
    .ZN(_12169_));
 BUF_X8 _34795_ (.A(_12149_),
    .Z(_12170_));
 OAI21_X2 _34796_ (.A(_11936_),
    .B1(_12170_),
    .B2(_00164_),
    .ZN(_12171_));
 BUF_X4 _34797_ (.A(_12092_),
    .Z(_12172_));
 BUF_X2 _34798_ (.A(\core.keymem.prev_key0_reg[123] ),
    .Z(_12173_));
 INV_X2 _34799_ (.A(_12173_),
    .ZN(_12174_));
 BUF_X4 _34800_ (.A(_11857_),
    .Z(_12175_));
 BUF_X4 _34801_ (.A(_12175_),
    .Z(_12176_));
 NOR2_X1 _34802_ (.A1(_12176_),
    .A2(_09949_),
    .ZN(_12177_));
 AOI21_X1 _34803_ (.A(_12177_),
    .B1(_12167_),
    .B2(_12176_),
    .ZN(_12178_));
 XNOR2_X1 _34804_ (.A(_12174_),
    .B(_12178_),
    .ZN(_12179_));
 NOR2_X1 _34805_ (.A1(_12172_),
    .A2(_12179_),
    .ZN(_12180_));
 OAI21_X4 _34806_ (.A(_12169_),
    .B1(_12171_),
    .B2(_12180_),
    .ZN(_12181_));
 BUF_X2 _34807_ (.A(_12181_),
    .Z(_12182_));
 OAI21_X1 _34808_ (.A(_12165_),
    .B1(_12182_),
    .B2(_11954_),
    .ZN(_00863_));
 BUF_X8 _34809_ (.A(_11804_),
    .Z(_12183_));
 BUF_X8 _34810_ (.A(_11874_),
    .Z(_12184_));
 BUF_X4 _34811_ (.A(_12184_),
    .Z(_12185_));
 BUF_X4 _34812_ (.A(_12185_),
    .Z(_12186_));
 NOR4_X2 _34813_ (.A1(_12183_),
    .A2(_16224_),
    .A3(_00165_),
    .A4(_12186_),
    .ZN(_12187_));
 AOI21_X1 _34814_ (.A(_12187_),
    .B1(_12005_),
    .B2(\core.keymem.key_mem[0][124] ),
    .ZN(_12188_));
 INV_X1 _34815_ (.A(_12188_),
    .ZN(_00864_));
 CLKBUF_X3 _34816_ (.A(_00167_),
    .Z(_12189_));
 NOR4_X4 _34817_ (.A1(_12183_),
    .A2(_16224_),
    .A3(_12189_),
    .A4(_12186_),
    .ZN(_12190_));
 AOI21_X1 _34818_ (.A(_12190_),
    .B1(_11933_),
    .B2(\core.keymem.key_mem[0][125] ),
    .ZN(_12191_));
 INV_X1 _34819_ (.A(_12191_),
    .ZN(_00865_));
 NAND2_X1 _34820_ (.A1(\core.keymem.key_mem[0][126] ),
    .A2(_11933_),
    .ZN(_12192_));
 BUF_X4 _34821_ (.A(_11799_),
    .Z(_12193_));
 BUF_X2 _34822_ (.A(\core.keymem.rcon_logic.tmp_rcon[7] ),
    .Z(_12194_));
 XNOR2_X2 _34823_ (.A(_12194_),
    .B(_09171_),
    .ZN(_12195_));
 XNOR2_X2 _34824_ (.A(\core.keymem.prev_key1_reg[126] ),
    .B(_12195_),
    .ZN(_12196_));
 AOI22_X2 _34825_ (.A1(_00169_),
    .A2(_12193_),
    .B1(_11889_),
    .B2(_12196_),
    .ZN(_12197_));
 NOR2_X1 _34826_ (.A1(_00170_),
    .A2(_11828_),
    .ZN(_12198_));
 OR2_X1 _34827_ (.A1(_11904_),
    .A2(_12198_),
    .ZN(_12199_));
 CLKBUF_X3 _34828_ (.A(\core.keymem.prev_key0_reg[126] ),
    .Z(_12200_));
 INV_X2 _34829_ (.A(_12200_),
    .ZN(_12201_));
 NOR2_X1 _34830_ (.A1(_12176_),
    .A2(_10221_),
    .ZN(_12202_));
 AOI21_X1 _34831_ (.A(_12202_),
    .B1(_12195_),
    .B2(_12176_),
    .ZN(_12203_));
 XNOR2_X1 _34832_ (.A(_12201_),
    .B(_12203_),
    .ZN(_12204_));
 NOR2_X2 _34833_ (.A1(_12172_),
    .A2(_12204_),
    .ZN(_12205_));
 OAI21_X4 _34834_ (.A(_12197_),
    .B1(_12199_),
    .B2(_12205_),
    .ZN(_12206_));
 CLKBUF_X3 _34835_ (.A(_12206_),
    .Z(_12207_));
 OAI21_X1 _34836_ (.A(_12192_),
    .B1(_12207_),
    .B2(_11954_),
    .ZN(_00866_));
 INV_X2 _34837_ (.A(_00171_),
    .ZN(_12208_));
 NAND3_X1 _34838_ (.A1(_16286_),
    .A2(_12208_),
    .A3(_11880_),
    .ZN(_12209_));
 INV_X1 _34839_ (.A(\core.keymem.key_mem[0][127] ),
    .ZN(_12210_));
 OAI21_X1 _34840_ (.A(_12209_),
    .B1(_11883_),
    .B2(_12210_),
    .ZN(_00867_));
 BUF_X4 _34841_ (.A(_11805_),
    .Z(_12211_));
 NOR2_X1 _34842_ (.A1(_12211_),
    .A2(_00407_),
    .ZN(_12212_));
 MUX2_X1 _34843_ (.A(\core.keymem.key_mem[0][12] ),
    .B(_12212_),
    .S(_12018_),
    .Z(_00868_));
 INV_X1 _34844_ (.A(_00408_),
    .ZN(_12213_));
 NAND3_X1 _34845_ (.A1(_16286_),
    .A2(_12213_),
    .A3(_11880_),
    .ZN(_12214_));
 INV_X1 _34846_ (.A(\core.keymem.key_mem[0][13] ),
    .ZN(_12215_));
 OAI21_X1 _34847_ (.A(_12214_),
    .B1(_11883_),
    .B2(_12215_),
    .ZN(_00869_));
 NOR2_X1 _34848_ (.A1(_12211_),
    .A2(_00409_),
    .ZN(_12216_));
 MUX2_X1 _34849_ (.A(\core.keymem.key_mem[0][14] ),
    .B(_12216_),
    .S(_12018_),
    .Z(_00870_));
 INV_X1 _34850_ (.A(_00410_),
    .ZN(_12217_));
 NAND3_X1 _34851_ (.A1(_16286_),
    .A2(_12217_),
    .A3(_11880_),
    .ZN(_12218_));
 INV_X1 _34852_ (.A(\core.keymem.key_mem[0][15] ),
    .ZN(_12219_));
 OAI21_X1 _34853_ (.A(_12218_),
    .B1(_11883_),
    .B2(_12219_),
    .ZN(_00871_));
 NOR2_X1 _34854_ (.A1(_12211_),
    .A2(_00411_),
    .ZN(_12220_));
 MUX2_X1 _34855_ (.A(\core.keymem.key_mem[0][16] ),
    .B(_12220_),
    .S(_12018_),
    .Z(_00872_));
 NOR2_X1 _34856_ (.A1(_12211_),
    .A2(_00434_),
    .ZN(_12221_));
 BUF_X4 _34857_ (.A(_11877_),
    .Z(_12222_));
 MUX2_X1 _34858_ (.A(\core.keymem.key_mem[0][17] ),
    .B(_12221_),
    .S(_12222_),
    .Z(_00873_));
 NOR2_X1 _34859_ (.A1(_12211_),
    .A2(_00435_),
    .ZN(_12223_));
 MUX2_X1 _34860_ (.A(\core.keymem.key_mem[0][18] ),
    .B(_12223_),
    .S(_12222_),
    .Z(_00874_));
 INV_X1 _34861_ (.A(_00436_),
    .ZN(_12224_));
 NAND3_X1 _34862_ (.A1(_16286_),
    .A2(_12224_),
    .A3(_11880_),
    .ZN(_12225_));
 INV_X1 _34863_ (.A(\core.keymem.key_mem[0][19] ),
    .ZN(_12226_));
 OAI21_X1 _34864_ (.A(_12225_),
    .B1(_11883_),
    .B2(_12226_),
    .ZN(_00875_));
 INV_X1 _34865_ (.A(_00371_),
    .ZN(_12227_));
 NAND3_X1 _34866_ (.A1(_16286_),
    .A2(_12227_),
    .A3(_11880_),
    .ZN(_12228_));
 INV_X1 _34867_ (.A(\core.keymem.key_mem[0][1] ),
    .ZN(_12229_));
 OAI21_X1 _34868_ (.A(_12228_),
    .B1(_11883_),
    .B2(_12229_),
    .ZN(_00876_));
 CLKBUF_X3 _34869_ (.A(_16285_),
    .Z(_12230_));
 INV_X1 _34870_ (.A(_00437_),
    .ZN(_12231_));
 NAND3_X1 _34871_ (.A1(_12230_),
    .A2(_12231_),
    .A3(_11880_),
    .ZN(_12232_));
 INV_X1 _34872_ (.A(\core.keymem.key_mem[0][20] ),
    .ZN(_12233_));
 OAI21_X1 _34873_ (.A(_12232_),
    .B1(_11883_),
    .B2(_12233_),
    .ZN(_00877_));
 NOR2_X1 _34874_ (.A1(_12211_),
    .A2(_00438_),
    .ZN(_12234_));
 MUX2_X1 _34875_ (.A(\core.keymem.key_mem[0][21] ),
    .B(_12234_),
    .S(_12222_),
    .Z(_00878_));
 INV_X2 _34876_ (.A(_00015_),
    .ZN(_12235_));
 CLKBUF_X3 _34877_ (.A(_11877_),
    .Z(_12236_));
 NAND3_X1 _34878_ (.A1(_12230_),
    .A2(_12235_),
    .A3(_12236_),
    .ZN(_12237_));
 BUF_X4 _34879_ (.A(_11882_),
    .Z(_12238_));
 INV_X1 _34880_ (.A(\core.keymem.key_mem[0][22] ),
    .ZN(_12239_));
 OAI21_X1 _34881_ (.A(_12237_),
    .B1(_12238_),
    .B2(_12239_),
    .ZN(_00879_));
 NAND2_X1 _34882_ (.A1(\core.keymem.key_mem[0][23] ),
    .A2(_11933_),
    .ZN(_12240_));
 NAND2_X4 _34883_ (.A1(_12044_),
    .A2(_11822_),
    .ZN(_12241_));
 CLKBUF_X2 _34884_ (.A(\core.keymem.prev_key0_reg[55] ),
    .Z(_12242_));
 INV_X1 _34885_ (.A(_12242_),
    .ZN(_12243_));
 BUF_X2 _34886_ (.A(\core.keymem.prev_key0_reg[87] ),
    .Z(_12244_));
 NOR4_X1 _34887_ (.A1(_12243_),
    .A2(_12244_),
    .A3(_12089_),
    .A4(_12090_),
    .ZN(_12245_));
 INV_X1 _34888_ (.A(_12244_),
    .ZN(_12246_));
 NOR4_X1 _34889_ (.A1(_12242_),
    .A2(_12246_),
    .A3(_12089_),
    .A4(_12090_),
    .ZN(_12247_));
 NAND3_X1 _34890_ (.A1(_12243_),
    .A2(_12246_),
    .A3(_12089_),
    .ZN(_12248_));
 NAND3_X1 _34891_ (.A1(_12242_),
    .A2(_12244_),
    .A3(_12089_),
    .ZN(_12249_));
 AOI21_X1 _34892_ (.A(_12090_),
    .B1(_12248_),
    .B2(_12249_),
    .ZN(_12250_));
 NAND4_X1 _34893_ (.A1(_12040_),
    .A2(_09188_),
    .A3(_09193_),
    .A4(_09208_),
    .ZN(_12251_));
 NOR3_X1 _34894_ (.A1(_12242_),
    .A2(_12244_),
    .A3(_12089_),
    .ZN(_12252_));
 NOR3_X1 _34895_ (.A1(_12243_),
    .A2(_12246_),
    .A3(_12089_),
    .ZN(_12253_));
 OAI221_X1 _34896_ (.A(_12251_),
    .B1(_12252_),
    .B2(_12253_),
    .C1(_08163_),
    .C2(_11832_),
    .ZN(_12254_));
 AND3_X1 _34897_ (.A1(_12242_),
    .A2(_12246_),
    .A3(_12089_),
    .ZN(_12255_));
 AND3_X1 _34898_ (.A1(_12243_),
    .A2(_12244_),
    .A3(_12089_),
    .ZN(_12256_));
 OAI221_X1 _34899_ (.A(_12251_),
    .B1(_12255_),
    .B2(_12256_),
    .C1(_08163_),
    .C2(_11832_),
    .ZN(_12257_));
 NAND2_X1 _34900_ (.A1(_12254_),
    .A2(_12257_),
    .ZN(_12258_));
 OR4_X2 _34901_ (.A1(_12245_),
    .A2(_12247_),
    .A3(_12250_),
    .A4(_12258_),
    .ZN(_12259_));
 XNOR2_X1 _34902_ (.A(\core.keymem.prev_key0_reg[23] ),
    .B(_12259_),
    .ZN(_12260_));
 NOR2_X2 _34903_ (.A1(_12241_),
    .A2(_12260_),
    .ZN(_12261_));
 BUF_X8 _34904_ (.A(_12184_),
    .Z(_12262_));
 BUF_X8 _34905_ (.A(_11814_),
    .Z(_12263_));
 XNOR2_X1 _34906_ (.A(\core.keymem.prev_key1_reg[87] ),
    .B(\core.keymem.prev_key1_reg[119] ),
    .ZN(_12264_));
 XNOR2_X2 _34907_ (.A(_08163_),
    .B(_12264_),
    .ZN(_12265_));
 XNOR2_X2 _34908_ (.A(\core.keymem.prev_key1_reg[55] ),
    .B(_12265_),
    .ZN(_12266_));
 XNOR2_X1 _34909_ (.A(_08293_),
    .B(_12266_),
    .ZN(_12267_));
 OAI22_X2 _34910_ (.A1(_00016_),
    .A2(_12262_),
    .B1(_12263_),
    .B2(_12267_),
    .ZN(_12268_));
 NOR2_X4 _34911_ (.A1(_11860_),
    .A2(_11903_),
    .ZN(_12269_));
 NAND2_X1 _34912_ (.A1(\core.key[23] ),
    .A2(_12269_),
    .ZN(_12270_));
 INV_X1 _34913_ (.A(_12270_),
    .ZN(_12271_));
 NOR3_X4 _34914_ (.A1(_12261_),
    .A2(_12268_),
    .A3(_12271_),
    .ZN(_12272_));
 OAI21_X1 _34915_ (.A(_12240_),
    .B1(_12272_),
    .B2(_11954_),
    .ZN(_00880_));
 NOR2_X1 _34916_ (.A1(_12211_),
    .A2(_00017_),
    .ZN(_12273_));
 MUX2_X1 _34917_ (.A(\core.keymem.key_mem[0][24] ),
    .B(_12273_),
    .S(_12222_),
    .Z(_00881_));
 INV_X1 _34918_ (.A(_00020_),
    .ZN(_12274_));
 NAND3_X1 _34919_ (.A1(_12230_),
    .A2(_12274_),
    .A3(_12236_),
    .ZN(_12275_));
 INV_X1 _34920_ (.A(\core.keymem.key_mem[0][25] ),
    .ZN(_12276_));
 OAI21_X1 _34921_ (.A(_12275_),
    .B1(_12238_),
    .B2(_12276_),
    .ZN(_00882_));
 NOR2_X2 _34922_ (.A1(_00023_),
    .A2(_11863_),
    .ZN(_12277_));
 XNOR2_X2 _34923_ (.A(\core.keymem.rcon_reg[2] ),
    .B(_08803_),
    .ZN(_12278_));
 BUF_X2 _34924_ (.A(\core.keymem.prev_key1_reg[90] ),
    .Z(_12279_));
 XOR2_X2 _34925_ (.A(\core.keymem.prev_key1_reg[58] ),
    .B(_12279_),
    .Z(_12280_));
 XOR2_X1 _34926_ (.A(\core.keymem.prev_key1_reg[26] ),
    .B(_00024_),
    .Z(_12281_));
 XNOR2_X1 _34927_ (.A(_12280_),
    .B(_12281_),
    .ZN(_12282_));
 XNOR2_X1 _34928_ (.A(_12278_),
    .B(_12282_),
    .ZN(_12283_));
 NOR2_X2 _34929_ (.A1(_11799_),
    .A2(_12283_),
    .ZN(_12284_));
 AOI21_X4 _34930_ (.A(_12277_),
    .B1(_12284_),
    .B2(_11847_),
    .ZN(_12285_));
 NOR2_X1 _34931_ (.A1(_11953_),
    .A2(_12285_),
    .ZN(_12286_));
 AOI21_X1 _34932_ (.A(_12286_),
    .B1(_11933_),
    .B2(\core.keymem.key_mem[0][26] ),
    .ZN(_12287_));
 INV_X1 _34933_ (.A(_12287_),
    .ZN(_00883_));
 NOR2_X1 _34934_ (.A1(_12211_),
    .A2(_00026_),
    .ZN(_12288_));
 MUX2_X1 _34935_ (.A(\core.keymem.key_mem[0][27] ),
    .B(_12288_),
    .S(_12222_),
    .Z(_00884_));
 NOR2_X1 _34936_ (.A1(_12211_),
    .A2(_00029_),
    .ZN(_12289_));
 MUX2_X1 _34937_ (.A(\core.keymem.key_mem[0][28] ),
    .B(_12289_),
    .S(_12222_),
    .Z(_00885_));
 NAND2_X1 _34938_ (.A1(\core.keymem.key_mem[0][29] ),
    .A2(_11933_),
    .ZN(_12290_));
 NOR2_X2 _34939_ (.A1(_00032_),
    .A2(_11813_),
    .ZN(_12291_));
 BUF_X8 _34940_ (.A(_11866_),
    .Z(_12292_));
 XOR2_X2 _34941_ (.A(\core.keymem.rcon_logic.tmp_rcon[6] ),
    .B(_09123_),
    .Z(_12293_));
 CLKBUF_X2 _34942_ (.A(\core.keymem.prev_key1_reg[93] ),
    .Z(_12294_));
 XOR2_X2 _34943_ (.A(\core.keymem.prev_key1_reg[61] ),
    .B(_12294_),
    .Z(_12295_));
 XNOR2_X1 _34944_ (.A(\core.keymem.prev_key1_reg[29] ),
    .B(_00033_),
    .ZN(_12296_));
 XNOR2_X1 _34945_ (.A(_12295_),
    .B(_12296_),
    .ZN(_12297_));
 XNOR2_X1 _34946_ (.A(_12293_),
    .B(_12297_),
    .ZN(_12298_));
 AOI21_X1 _34947_ (.A(_12291_),
    .B1(_12298_),
    .B2(_11862_),
    .ZN(_12299_));
 NAND2_X1 _34948_ (.A1(_12292_),
    .A2(_12299_),
    .ZN(_12300_));
 BUF_X4 _34949_ (.A(_06677_),
    .Z(_12301_));
 NAND2_X2 _34950_ (.A1(_11813_),
    .A2(_11819_),
    .ZN(_12302_));
 OR2_X1 _34951_ (.A1(_00034_),
    .A2(_12302_),
    .ZN(_12303_));
 NAND2_X1 _34952_ (.A1(_12301_),
    .A2(_12303_),
    .ZN(_12304_));
 MUX2_X1 _34953_ (.A(_10075_),
    .B(_12293_),
    .S(_11920_),
    .Z(_12305_));
 XOR2_X2 _34954_ (.A(\core.keymem.prev_key0_reg[125] ),
    .B(_12305_),
    .Z(_12306_));
 BUF_X2 _34955_ (.A(\core.keymem.prev_key0_reg[93] ),
    .Z(_12307_));
 XNOR2_X2 _34956_ (.A(\core.keymem.prev_key0_reg[61] ),
    .B(_12307_),
    .ZN(_12308_));
 XNOR2_X2 _34957_ (.A(\core.keymem.prev_key0_reg[29] ),
    .B(_12308_),
    .ZN(_12309_));
 XOR2_X1 _34958_ (.A(_12306_),
    .B(_12309_),
    .Z(_12310_));
 NOR2_X4 _34959_ (.A1(_11820_),
    .A2(_11903_),
    .ZN(_12311_));
 AOI221_X2 _34960_ (.A(_12291_),
    .B1(_12300_),
    .B2(_12304_),
    .C1(_12310_),
    .C2(_12311_),
    .ZN(_12312_));
 OAI21_X1 _34961_ (.A(_12290_),
    .B1(_12312_),
    .B2(_11954_),
    .ZN(_00886_));
 BUF_X4 _34962_ (.A(_11801_),
    .Z(_12313_));
 NAND2_X1 _34963_ (.A1(\core.keymem.key_mem[0][2] ),
    .A2(_12313_),
    .ZN(_12314_));
 XNOR2_X1 _34964_ (.A(\core.keymem.prev_key1_reg[66] ),
    .B(\core.keymem.prev_key1_reg[98] ),
    .ZN(_12315_));
 XNOR2_X2 _34965_ (.A(_09859_),
    .B(_12315_),
    .ZN(_12316_));
 XNOR2_X2 _34966_ (.A(\core.keymem.prev_key1_reg[34] ),
    .B(_12316_),
    .ZN(_12317_));
 XNOR2_X1 _34967_ (.A(\core.keymem.prev_key1_reg[2] ),
    .B(_12317_),
    .ZN(_12318_));
 OAI22_X2 _34968_ (.A1(_00373_),
    .A2(_12262_),
    .B1(_12263_),
    .B2(_12318_),
    .ZN(_12319_));
 INV_X1 _34969_ (.A(\core.keymem.prev_key0_reg[98] ),
    .ZN(_12320_));
 NAND3_X4 _34970_ (.A1(_11832_),
    .A2(_11939_),
    .A3(_11941_),
    .ZN(_12321_));
 NAND3_X2 _34971_ (.A1(_11857_),
    .A2(_09808_),
    .A3(_09858_),
    .ZN(_12322_));
 NAND2_X2 _34972_ (.A1(_12321_),
    .A2(_12322_),
    .ZN(_12323_));
 XNOR2_X2 _34973_ (.A(_12320_),
    .B(_12323_),
    .ZN(_12324_));
 CLKBUF_X2 _34974_ (.A(\core.keymem.prev_key0_reg[66] ),
    .Z(_12325_));
 INV_X1 _34975_ (.A(_12325_),
    .ZN(_12326_));
 NAND2_X1 _34976_ (.A1(\core.keymem.prev_key0_reg[34] ),
    .A2(_12326_),
    .ZN(_12327_));
 INV_X1 _34977_ (.A(\core.keymem.prev_key0_reg[34] ),
    .ZN(_12328_));
 NAND2_X1 _34978_ (.A1(_12328_),
    .A2(_12325_),
    .ZN(_12329_));
 AND2_X1 _34979_ (.A1(_12327_),
    .A2(_12329_),
    .ZN(_12330_));
 XNOR2_X1 _34980_ (.A(\core.keymem.prev_key0_reg[2] ),
    .B(_12330_),
    .ZN(_12331_));
 XNOR2_X1 _34981_ (.A(_12324_),
    .B(_12331_),
    .ZN(_12332_));
 BUF_X4 _34982_ (.A(_11945_),
    .Z(_12333_));
 MUX2_X2 _34983_ (.A(\core.key[2] ),
    .B(_12332_),
    .S(_12333_),
    .Z(_12334_));
 BUF_X8 _34984_ (.A(_12098_),
    .Z(_12335_));
 BUF_X4 _34985_ (.A(_12335_),
    .Z(_12336_));
 AOI21_X4 _34986_ (.A(_12319_),
    .B1(_12334_),
    .B2(_12336_),
    .ZN(_12337_));
 OAI21_X1 _34987_ (.A(_12314_),
    .B1(_12337_),
    .B2(_11954_),
    .ZN(_00887_));
 NOR2_X1 _34988_ (.A1(_12211_),
    .A2(_00035_),
    .ZN(_12338_));
 MUX2_X1 _34989_ (.A(\core.keymem.key_mem[0][30] ),
    .B(_12338_),
    .S(_12222_),
    .Z(_00888_));
 CLKBUF_X3 _34990_ (.A(_11805_),
    .Z(_12339_));
 NOR2_X1 _34991_ (.A1(_12339_),
    .A2(_00038_),
    .ZN(_12340_));
 MUX2_X1 _34992_ (.A(\core.keymem.key_mem[0][31] ),
    .B(_12340_),
    .S(_12222_),
    .Z(_00889_));
 NAND2_X1 _34993_ (.A1(\core.keymem.key_mem[0][32] ),
    .A2(_12313_),
    .ZN(_12341_));
 INV_X1 _34994_ (.A(\core.key[32] ),
    .ZN(_12342_));
 AOI21_X1 _34995_ (.A(_11987_),
    .B1(_11989_),
    .B2(_12342_),
    .ZN(_12343_));
 XNOR2_X1 _34996_ (.A(_11835_),
    .B(_11836_),
    .ZN(_12344_));
 BUF_X4 _34997_ (.A(_12092_),
    .Z(_12345_));
 OAI21_X2 _34998_ (.A(_12343_),
    .B1(_12344_),
    .B2(_12345_),
    .ZN(_12346_));
 BUF_X8 _34999_ (.A(_11874_),
    .Z(_12347_));
 OR2_X1 _35000_ (.A1(_00041_),
    .A2(_12347_),
    .ZN(_12348_));
 BUF_X4 _35001_ (.A(_06676_),
    .Z(_12349_));
 INV_X1 _35002_ (.A(\core.keymem.prev_key1_reg[96] ),
    .ZN(_12350_));
 XNOR2_X2 _35003_ (.A(_12350_),
    .B(_09681_),
    .ZN(_12351_));
 XNOR2_X1 _35004_ (.A(_11807_),
    .B(_12351_),
    .ZN(_12352_));
 OR3_X2 _35005_ (.A1(_12349_),
    .A2(_11799_),
    .A3(_12352_),
    .ZN(_12353_));
 NAND3_X4 _35006_ (.A1(_12346_),
    .A2(_12348_),
    .A3(_12353_),
    .ZN(_12354_));
 NAND2_X1 _35007_ (.A1(_16285_),
    .A2(_12354_),
    .ZN(_12355_));
 OAI21_X1 _35008_ (.A(_12341_),
    .B1(_12355_),
    .B2(_12005_),
    .ZN(_00890_));
 NAND2_X1 _35009_ (.A1(\core.keymem.key_mem[0][33] ),
    .A2(_12313_),
    .ZN(_12356_));
 NOR2_X2 _35010_ (.A1(_00042_),
    .A2(_11960_),
    .ZN(_12357_));
 XOR2_X2 _35011_ (.A(\core.keymem.prev_key1_reg[97] ),
    .B(_09777_),
    .Z(_12358_));
 XNOR2_X2 _35012_ (.A(\core.keymem.prev_key1_reg[33] ),
    .B(\core.keymem.prev_key1_reg[65] ),
    .ZN(_12359_));
 XNOR2_X2 _35013_ (.A(_12358_),
    .B(_12359_),
    .ZN(_12360_));
 AOI21_X4 _35014_ (.A(_12357_),
    .B1(_12360_),
    .B2(_12027_),
    .ZN(_12361_));
 OAI21_X1 _35015_ (.A(_12356_),
    .B1(_12361_),
    .B2(_11954_),
    .ZN(_00891_));
 NAND2_X1 _35016_ (.A1(\core.keymem.key_mem[0][34] ),
    .A2(_12313_),
    .ZN(_12362_));
 NOR2_X1 _35017_ (.A1(_00043_),
    .A2(_11960_),
    .ZN(_12363_));
 AOI21_X2 _35018_ (.A(_12363_),
    .B1(_12317_),
    .B2(_11889_),
    .ZN(_12364_));
 BUF_X8 _35019_ (.A(_11828_),
    .Z(_12365_));
 OAI21_X2 _35020_ (.A(_12098_),
    .B1(_12365_),
    .B2(\core.key[34] ),
    .ZN(_12366_));
 AOI221_X1 _35021_ (.A(\core.keymem.prev_key0_reg[98] ),
    .B1(_12321_),
    .B2(_12322_),
    .C1(_12327_),
    .C2(_12329_),
    .ZN(_12367_));
 NAND2_X1 _35022_ (.A1(_12328_),
    .A2(_12326_),
    .ZN(_12368_));
 NAND2_X1 _35023_ (.A1(\core.keymem.prev_key0_reg[34] ),
    .A2(_12325_),
    .ZN(_12369_));
 AOI221_X1 _35024_ (.A(_12320_),
    .B1(_12321_),
    .B2(_12322_),
    .C1(_12368_),
    .C2(_12369_),
    .ZN(_12370_));
 OR2_X1 _35025_ (.A1(_12367_),
    .A2(_12370_),
    .ZN(_12371_));
 AOI211_X2 _35026_ (.A(\core.keymem.prev_key0_reg[98] ),
    .B(_12323_),
    .C1(_12368_),
    .C2(_12369_),
    .ZN(_12372_));
 AOI211_X2 _35027_ (.A(_12320_),
    .B(_12323_),
    .C1(_12327_),
    .C2(_12329_),
    .ZN(_12373_));
 NOR4_X4 _35028_ (.A1(_11989_),
    .A2(_12371_),
    .A3(_12372_),
    .A4(_12373_),
    .ZN(_12374_));
 OAI21_X4 _35029_ (.A(_12364_),
    .B1(_12366_),
    .B2(_12374_),
    .ZN(_12375_));
 NAND2_X1 _35030_ (.A1(_16285_),
    .A2(_12375_),
    .ZN(_12376_));
 OAI21_X1 _35031_ (.A(_12362_),
    .B1(_12376_),
    .B2(_12005_),
    .ZN(_00892_));
 NAND2_X1 _35032_ (.A1(\core.keymem.key_mem[0][35] ),
    .A2(_12313_),
    .ZN(_12377_));
 NAND3_X2 _35033_ (.A1(_12040_),
    .A2(_10329_),
    .A3(_10351_),
    .ZN(_12378_));
 AND4_X1 _35034_ (.A1(_09877_),
    .A2(_09890_),
    .A3(_09904_),
    .A4(_09933_),
    .ZN(_12379_));
 NOR3_X1 _35035_ (.A1(_09718_),
    .A2(_09941_),
    .A3(_09947_),
    .ZN(_12380_));
 NAND3_X1 _35036_ (.A1(_11851_),
    .A2(_12379_),
    .A3(_12380_),
    .ZN(_12381_));
 NAND2_X1 _35037_ (.A1(_12378_),
    .A2(_12381_),
    .ZN(_12382_));
 BUF_X2 _35038_ (.A(\core.keymem.prev_key0_reg[35] ),
    .Z(_12383_));
 BUF_X2 _35039_ (.A(\core.keymem.prev_key0_reg[67] ),
    .Z(_12384_));
 CLKBUF_X2 _35040_ (.A(\core.keymem.prev_key0_reg[99] ),
    .Z(_12385_));
 NOR4_X1 _35041_ (.A1(_12383_),
    .A2(_12384_),
    .A3(_12385_),
    .A4(_11820_),
    .ZN(_12386_));
 NAND2_X1 _35042_ (.A1(_12383_),
    .A2(_12384_),
    .ZN(_12387_));
 NOR3_X1 _35043_ (.A1(_12385_),
    .A2(_11892_),
    .A3(_12387_),
    .ZN(_12388_));
 OAI21_X1 _35044_ (.A(_12382_),
    .B1(_12386_),
    .B2(_12388_),
    .ZN(_12389_));
 AND3_X1 _35045_ (.A1(_12063_),
    .A2(_10329_),
    .A3(_10351_),
    .ZN(_12390_));
 NOR3_X2 _35046_ (.A1(_11831_),
    .A2(_09934_),
    .A3(_09948_),
    .ZN(_12391_));
 INV_X1 _35047_ (.A(_12383_),
    .ZN(_12392_));
 INV_X1 _35048_ (.A(_12385_),
    .ZN(_12393_));
 NOR3_X1 _35049_ (.A1(_12392_),
    .A2(_12384_),
    .A3(_12393_),
    .ZN(_12394_));
 INV_X1 _35050_ (.A(_12384_),
    .ZN(_12395_));
 NOR3_X1 _35051_ (.A1(_12383_),
    .A2(_12395_),
    .A3(_12393_),
    .ZN(_12396_));
 OAI221_X2 _35052_ (.A(_12333_),
    .B1(_12390_),
    .B2(_12391_),
    .C1(_12394_),
    .C2(_12396_),
    .ZN(_12397_));
 NAND3_X1 _35053_ (.A1(_12383_),
    .A2(_12395_),
    .A3(_12393_),
    .ZN(_12398_));
 NAND3_X1 _35054_ (.A1(_12392_),
    .A2(_12384_),
    .A3(_12393_),
    .ZN(_12399_));
 AOI221_X2 _35055_ (.A(_12382_),
    .B1(_12398_),
    .B2(_12399_),
    .C1(_11812_),
    .C2(_11816_),
    .ZN(_12400_));
 NAND4_X1 _35056_ (.A1(_12392_),
    .A2(_12395_),
    .A3(_12385_),
    .A4(_11925_),
    .ZN(_12401_));
 OR3_X1 _35057_ (.A1(_12393_),
    .A2(_11819_),
    .A3(_12387_),
    .ZN(_12402_));
 AOI21_X1 _35058_ (.A(_12382_),
    .B1(_12401_),
    .B2(_12402_),
    .ZN(_12403_));
 NOR2_X1 _35059_ (.A1(_12400_),
    .A2(_12403_),
    .ZN(_12404_));
 INV_X1 _35060_ (.A(\core.key[35] ),
    .ZN(_12405_));
 AOI21_X2 _35061_ (.A(_11987_),
    .B1(_11989_),
    .B2(_12405_),
    .ZN(_12406_));
 NAND4_X4 _35062_ (.A1(_12389_),
    .A2(_12397_),
    .A3(_12404_),
    .A4(_12406_),
    .ZN(_12407_));
 NOR2_X1 _35063_ (.A1(_00044_),
    .A2(_11863_),
    .ZN(_12408_));
 XNOR2_X1 _35064_ (.A(\core.keymem.prev_key1_reg[67] ),
    .B(\core.keymem.prev_key1_reg[99] ),
    .ZN(_12409_));
 XNOR2_X2 _35065_ (.A(_09949_),
    .B(_12409_),
    .ZN(_12410_));
 XNOR2_X2 _35066_ (.A(\core.keymem.prev_key1_reg[35] ),
    .B(_12410_),
    .ZN(_12411_));
 AOI21_X2 _35067_ (.A(_12408_),
    .B1(_12411_),
    .B2(_11889_),
    .ZN(_12412_));
 AND2_X2 _35068_ (.A1(_12407_),
    .A2(_12412_),
    .ZN(_12413_));
 OAI21_X1 _35069_ (.A(_12377_),
    .B1(_12413_),
    .B2(_11954_),
    .ZN(_00893_));
 NOR2_X1 _35070_ (.A1(_00045_),
    .A2(_11960_),
    .ZN(_12414_));
 XNOR2_X1 _35071_ (.A(\core.keymem.prev_key1_reg[68] ),
    .B(\core.keymem.prev_key1_reg[100] ),
    .ZN(_12415_));
 XNOR2_X2 _35072_ (.A(_10009_),
    .B(_12415_),
    .ZN(_12416_));
 XNOR2_X2 _35073_ (.A(\core.keymem.prev_key1_reg[36] ),
    .B(_12416_),
    .ZN(_12417_));
 XNOR2_X2 _35074_ (.A(\core.keymem.prev_key0_reg[68] ),
    .B(\core.keymem.prev_key0_reg[100] ),
    .ZN(_12418_));
 XNOR2_X2 _35075_ (.A(\core.keymem.prev_key0_reg[36] ),
    .B(_12418_),
    .ZN(_12419_));
 XNOR2_X1 _35076_ (.A(_11858_),
    .B(_12419_),
    .ZN(_12420_));
 MUX2_X1 _35077_ (.A(\core.key[36] ),
    .B(_12420_),
    .S(_11945_),
    .Z(_12421_));
 AOI221_X2 _35078_ (.A(_12414_),
    .B1(_12417_),
    .B2(_12027_),
    .C1(_12421_),
    .C2(_11936_),
    .ZN(_12422_));
 NOR2_X1 _35079_ (.A1(_12183_),
    .A2(_12422_),
    .ZN(_12423_));
 MUX2_X1 _35080_ (.A(\core.keymem.key_mem[0][36] ),
    .B(_12423_),
    .S(_12222_),
    .Z(_00894_));
 NAND2_X1 _35081_ (.A1(\core.keymem.key_mem[0][37] ),
    .A2(_12313_),
    .ZN(_12424_));
 OAI21_X1 _35082_ (.A(_11823_),
    .B1(_11900_),
    .B2(\core.key[37] ),
    .ZN(_12425_));
 NAND4_X1 _35083_ (.A1(_11830_),
    .A2(_10431_),
    .A3(_10449_),
    .A4(_10467_),
    .ZN(_12426_));
 OAI33_X1 _35084_ (.A1(_12040_),
    .A2(_09569_),
    .A3(_10074_),
    .B1(_12426_),
    .B2(_07073_),
    .B3(_07044_),
    .ZN(_12427_));
 XNOR2_X2 _35085_ (.A(\core.keymem.prev_key0_reg[101] ),
    .B(net10),
    .ZN(_12428_));
 XOR2_X2 _35086_ (.A(\core.keymem.prev_key0_reg[69] ),
    .B(_12428_),
    .Z(_12429_));
 XNOR2_X1 _35087_ (.A(\core.keymem.prev_key0_reg[37] ),
    .B(_12429_),
    .ZN(_12430_));
 AOI21_X2 _35088_ (.A(_12425_),
    .B1(_12430_),
    .B2(_12333_),
    .ZN(_12431_));
 NOR2_X2 _35089_ (.A1(_00046_),
    .A2(_11863_),
    .ZN(_12432_));
 XOR2_X2 _35090_ (.A(\core.keymem.prev_key1_reg[101] ),
    .B(_10075_),
    .Z(_12433_));
 BUF_X2 _35091_ (.A(\core.keymem.prev_key1_reg[69] ),
    .Z(_12434_));
 XNOR2_X2 _35092_ (.A(\core.keymem.prev_key1_reg[37] ),
    .B(_12434_),
    .ZN(_12435_));
 XNOR2_X1 _35093_ (.A(_12433_),
    .B(_12435_),
    .ZN(_12436_));
 AND2_X1 _35094_ (.A1(_11888_),
    .A2(_12436_),
    .ZN(_12437_));
 NOR3_X4 _35095_ (.A1(_12431_),
    .A2(_12432_),
    .A3(_12437_),
    .ZN(_12438_));
 CLKBUF_X3 _35096_ (.A(_12438_),
    .Z(_12439_));
 OAI21_X1 _35097_ (.A(_12424_),
    .B1(_12439_),
    .B2(_11954_),
    .ZN(_00895_));
 NAND2_X1 _35098_ (.A1(\core.keymem.key_mem[0][38] ),
    .A2(_12313_),
    .ZN(_12440_));
 NOR2_X1 _35099_ (.A1(\core.key[38] ),
    .A2(_12149_),
    .ZN(_12441_));
 BUF_X1 _35100_ (.A(\core.keymem.prev_key0_reg[38] ),
    .Z(_12442_));
 BUF_X1 _35101_ (.A(\core.keymem.prev_key0_reg[70] ),
    .Z(_12443_));
 INV_X1 _35102_ (.A(_12443_),
    .ZN(_12444_));
 NAND2_X1 _35103_ (.A1(_12442_),
    .A2(_12444_),
    .ZN(_12445_));
 INV_X1 _35104_ (.A(_12442_),
    .ZN(_12446_));
 NAND2_X1 _35105_ (.A1(_12446_),
    .A2(_12443_),
    .ZN(_12447_));
 AOI221_X2 _35106_ (.A(_11894_),
    .B1(_11895_),
    .B2(_11897_),
    .C1(_12445_),
    .C2(_12447_),
    .ZN(_12448_));
 INV_X1 _35107_ (.A(_11894_),
    .ZN(_12449_));
 NAND2_X1 _35108_ (.A1(_12446_),
    .A2(_12444_),
    .ZN(_12450_));
 NAND2_X1 _35109_ (.A1(_12442_),
    .A2(_12443_),
    .ZN(_12451_));
 AOI221_X2 _35110_ (.A(_12449_),
    .B1(_11895_),
    .B2(_11897_),
    .C1(_12450_),
    .C2(_12451_),
    .ZN(_12452_));
 NOR4_X4 _35111_ (.A1(_11851_),
    .A2(_07044_),
    .A3(_08916_),
    .A4(_10525_),
    .ZN(_12453_));
 NAND3_X1 _35112_ (.A1(_12446_),
    .A2(_12444_),
    .A3(_12449_),
    .ZN(_12454_));
 OR2_X1 _35113_ (.A1(_11894_),
    .A2(_12451_),
    .ZN(_12455_));
 AOI221_X2 _35114_ (.A(_12453_),
    .B1(_12454_),
    .B2(_12455_),
    .C1(_10221_),
    .C2(_11920_),
    .ZN(_12456_));
 NAND3_X1 _35115_ (.A1(_12442_),
    .A2(_12444_),
    .A3(_11894_),
    .ZN(_12457_));
 NAND3_X1 _35116_ (.A1(_12446_),
    .A2(_12443_),
    .A3(_11894_),
    .ZN(_12458_));
 AOI221_X2 _35117_ (.A(_12453_),
    .B1(_12457_),
    .B2(_12458_),
    .C1(_10221_),
    .C2(_11920_),
    .ZN(_12459_));
 NOR4_X4 _35118_ (.A1(_12448_),
    .A2(_12452_),
    .A3(_12456_),
    .A4(_12459_),
    .ZN(_12460_));
 AOI21_X1 _35119_ (.A(_12441_),
    .B1(_12460_),
    .B2(_11901_),
    .ZN(_12461_));
 NAND2_X2 _35120_ (.A1(_11936_),
    .A2(_12461_),
    .ZN(_12462_));
 NOR2_X1 _35121_ (.A1(_00047_),
    .A2(_11863_),
    .ZN(_12463_));
 CLKBUF_X2 _35122_ (.A(\core.keymem.prev_key1_reg[70] ),
    .Z(_12464_));
 XOR2_X2 _35123_ (.A(\core.keymem.prev_key1_reg[38] ),
    .B(_12464_),
    .Z(_12465_));
 XOR2_X2 _35124_ (.A(_11887_),
    .B(_12465_),
    .Z(_12466_));
 AOI21_X2 _35125_ (.A(_12463_),
    .B1(_12466_),
    .B2(_11889_),
    .ZN(_12467_));
 AND2_X1 _35126_ (.A1(_12462_),
    .A2(_12467_),
    .ZN(_12468_));
 OAI21_X1 _35127_ (.A(_12440_),
    .B1(_12468_),
    .B2(_11954_),
    .ZN(_00896_));
 NOR2_X1 _35128_ (.A1(_12339_),
    .A2(_00048_),
    .ZN(_12469_));
 MUX2_X1 _35129_ (.A(\core.keymem.key_mem[0][39] ),
    .B(_12469_),
    .S(_12222_),
    .Z(_00897_));
 INV_X2 _35130_ (.A(_00374_),
    .ZN(_12470_));
 NAND3_X1 _35131_ (.A1(_12230_),
    .A2(_12470_),
    .A3(_12236_),
    .ZN(_12471_));
 INV_X1 _35132_ (.A(\core.keymem.key_mem[0][3] ),
    .ZN(_12472_));
 OAI21_X1 _35133_ (.A(_12471_),
    .B1(_12238_),
    .B2(_12472_),
    .ZN(_00898_));
 NOR2_X1 _35134_ (.A1(_12339_),
    .A2(_00049_),
    .ZN(_12473_));
 BUF_X4 _35135_ (.A(_11877_),
    .Z(_12474_));
 MUX2_X1 _35136_ (.A(\core.keymem.key_mem[0][40] ),
    .B(_12473_),
    .S(_12474_),
    .Z(_00899_));
 NOR2_X1 _35137_ (.A1(_12339_),
    .A2(_00050_),
    .ZN(_12475_));
 MUX2_X1 _35138_ (.A(\core.keymem.key_mem[0][41] ),
    .B(_12475_),
    .S(_12474_),
    .Z(_00900_));
 INV_X1 _35139_ (.A(_00051_),
    .ZN(_12476_));
 NAND3_X1 _35140_ (.A1(_12230_),
    .A2(_12476_),
    .A3(_12236_),
    .ZN(_12477_));
 INV_X1 _35141_ (.A(\core.keymem.key_mem[0][42] ),
    .ZN(_12478_));
 OAI21_X1 _35142_ (.A(_12477_),
    .B1(_12238_),
    .B2(_12478_),
    .ZN(_00901_));
 NOR2_X1 _35143_ (.A1(_12339_),
    .A2(_00052_),
    .ZN(_12479_));
 MUX2_X1 _35144_ (.A(\core.keymem.key_mem[0][43] ),
    .B(_12479_),
    .S(_12474_),
    .Z(_00902_));
 NAND2_X1 _35145_ (.A1(\core.keymem.key_mem[0][44] ),
    .A2(_12313_),
    .ZN(_12480_));
 BUF_X2 _35146_ (.A(\core.keymem.prev_key0_reg[44] ),
    .Z(_12481_));
 BUF_X2 _35147_ (.A(\core.keymem.prev_key0_reg[76] ),
    .Z(_12482_));
 NOR3_X1 _35148_ (.A1(_12481_),
    .A2(_12482_),
    .A3(_11969_),
    .ZN(_12483_));
 INV_X1 _35149_ (.A(_12481_),
    .ZN(_12484_));
 INV_X1 _35150_ (.A(_12482_),
    .ZN(_12485_));
 NOR3_X1 _35151_ (.A1(_12484_),
    .A2(_12485_),
    .A3(_11969_),
    .ZN(_12486_));
 OAI221_X1 _35152_ (.A(_12044_),
    .B1(_11971_),
    .B2(_11972_),
    .C1(_12483_),
    .C2(_12486_),
    .ZN(_12487_));
 NOR3_X1 _35153_ (.A1(_12484_),
    .A2(_12482_),
    .A3(_11970_),
    .ZN(_12488_));
 NOR3_X1 _35154_ (.A1(_12481_),
    .A2(_12485_),
    .A3(_11970_),
    .ZN(_12489_));
 OAI221_X1 _35155_ (.A(_11925_),
    .B1(_11971_),
    .B2(_11972_),
    .C1(_12488_),
    .C2(_12489_),
    .ZN(_12490_));
 NAND2_X1 _35156_ (.A1(_12487_),
    .A2(_12490_),
    .ZN(_12491_));
 NAND3_X1 _35157_ (.A1(_12481_),
    .A2(_12485_),
    .A3(_11970_),
    .ZN(_12492_));
 NAND3_X1 _35158_ (.A1(_12484_),
    .A2(_12482_),
    .A3(_11970_),
    .ZN(_12493_));
 AOI221_X2 _35159_ (.A(_11973_),
    .B1(_12492_),
    .B2(_12493_),
    .C1(_11812_),
    .C2(_11816_),
    .ZN(_12494_));
 NAND4_X1 _35160_ (.A1(_12484_),
    .A2(_12485_),
    .A3(_11969_),
    .A4(_11860_),
    .ZN(_12495_));
 NAND4_X1 _35161_ (.A1(_12481_),
    .A2(_12482_),
    .A3(_11969_),
    .A4(_11848_),
    .ZN(_12496_));
 AOI21_X2 _35162_ (.A(_11973_),
    .B1(_12495_),
    .B2(_12496_),
    .ZN(_12497_));
 OAI21_X2 _35163_ (.A(_11823_),
    .B1(_12044_),
    .B2(\core.key[44] ),
    .ZN(_12498_));
 NOR4_X4 _35164_ (.A1(_12491_),
    .A2(_12494_),
    .A3(_12497_),
    .A4(_12498_),
    .ZN(_12499_));
 NOR2_X2 _35165_ (.A1(_00053_),
    .A2(_11885_),
    .ZN(_12500_));
 XNOR2_X1 _35166_ (.A(\core.keymem.prev_key1_reg[76] ),
    .B(\core.keymem.prev_key1_reg[108] ),
    .ZN(_12501_));
 XNOR2_X2 _35167_ (.A(_10413_),
    .B(_12501_),
    .ZN(_12502_));
 XNOR2_X2 _35168_ (.A(\core.keymem.prev_key1_reg[44] ),
    .B(_12502_),
    .ZN(_12503_));
 NOR2_X1 _35169_ (.A1(_12001_),
    .A2(_12503_),
    .ZN(_12504_));
 OR3_X4 _35170_ (.A1(_12499_),
    .A2(_12500_),
    .A3(_12504_),
    .ZN(_12505_));
 NAND2_X1 _35171_ (.A1(_16285_),
    .A2(_12505_),
    .ZN(_12506_));
 OAI21_X1 _35172_ (.A(_12480_),
    .B1(_12506_),
    .B2(_12005_),
    .ZN(_00903_));
 NOR3_X1 _35173_ (.A1(_11930_),
    .A2(_00054_),
    .A3(_11801_),
    .ZN(_12507_));
 AOI21_X1 _35174_ (.A(_12507_),
    .B1(_11933_),
    .B2(\core.keymem.key_mem[0][45] ),
    .ZN(_12508_));
 INV_X1 _35175_ (.A(_12508_),
    .ZN(_00904_));
 NOR2_X1 _35176_ (.A1(_12339_),
    .A2(_00055_),
    .ZN(_12509_));
 MUX2_X1 _35177_ (.A(\core.keymem.key_mem[0][46] ),
    .B(_12509_),
    .S(_12474_),
    .Z(_00905_));
 NAND2_X1 _35178_ (.A1(\core.keymem.key_mem[0][47] ),
    .A2(_12313_),
    .ZN(_12510_));
 OAI21_X1 _35179_ (.A(_12098_),
    .B1(_12149_),
    .B2(\core.key[47] ),
    .ZN(_12511_));
 XNOR2_X2 _35180_ (.A(\core.keymem.prev_key0_reg[79] ),
    .B(_12013_),
    .ZN(_12512_));
 XOR2_X2 _35181_ (.A(\core.keymem.prev_key0_reg[47] ),
    .B(_12512_),
    .Z(_12513_));
 AOI21_X2 _35182_ (.A(_12511_),
    .B1(_12513_),
    .B2(_12365_),
    .ZN(_12514_));
 XNOR2_X1 _35183_ (.A(\core.keymem.prev_key1_reg[79] ),
    .B(\core.keymem.prev_key1_reg[111] ),
    .ZN(_12515_));
 XNOR2_X2 _35184_ (.A(_10565_),
    .B(_12515_),
    .ZN(_12516_));
 XNOR2_X2 _35185_ (.A(\core.keymem.prev_key1_reg[47] ),
    .B(_12516_),
    .ZN(_12517_));
 OAI22_X4 _35186_ (.A1(_00056_),
    .A2(_12184_),
    .B1(_12001_),
    .B2(_12517_),
    .ZN(_12518_));
 OAI21_X4 _35187_ (.A(_16229_),
    .B1(_12514_),
    .B2(_12518_),
    .ZN(_12519_));
 CLKBUF_X3 _35188_ (.A(_12519_),
    .Z(_12520_));
 OAI21_X1 _35189_ (.A(_12510_),
    .B1(_12520_),
    .B2(_12005_),
    .ZN(_00906_));
 NAND2_X1 _35190_ (.A1(\core.keymem.key_mem[0][48] ),
    .A2(_12313_),
    .ZN(_12521_));
 XOR2_X2 _35191_ (.A(\core.keymem.prev_key0_reg[80] ),
    .B(_12021_),
    .Z(_12522_));
 XNOR2_X1 _35192_ (.A(\core.keymem.prev_key0_reg[48] ),
    .B(_12522_),
    .ZN(_12523_));
 OR2_X1 _35193_ (.A1(_12241_),
    .A2(_12523_),
    .ZN(_12524_));
 NOR2_X2 _35194_ (.A1(_00057_),
    .A2(_11862_),
    .ZN(_12525_));
 BUF_X2 _35195_ (.A(\core.keymem.prev_key1_reg[48] ),
    .Z(_12526_));
 BUF_X2 _35196_ (.A(\core.keymem.prev_key1_reg[80] ),
    .Z(_12527_));
 XNOR2_X2 _35197_ (.A(_12527_),
    .B(_12026_),
    .ZN(_12528_));
 XNOR2_X1 _35198_ (.A(_12526_),
    .B(_12528_),
    .ZN(_12529_));
 AOI221_X2 _35199_ (.A(_12525_),
    .B1(_12529_),
    .B2(_11888_),
    .C1(_12269_),
    .C2(\core.key[48] ),
    .ZN(_12530_));
 AND2_X4 _35200_ (.A1(_12524_),
    .A2(_12530_),
    .ZN(_12531_));
 CLKBUF_X3 _35201_ (.A(_12531_),
    .Z(_12532_));
 BUF_X4 _35202_ (.A(_11953_),
    .Z(_12533_));
 OAI21_X1 _35203_ (.A(_12521_),
    .B1(_12532_),
    .B2(_12533_),
    .ZN(_00907_));
 NOR2_X1 _35204_ (.A1(_12339_),
    .A2(_00058_),
    .ZN(_12534_));
 MUX2_X1 _35205_ (.A(\core.keymem.key_mem[0][49] ),
    .B(_12534_),
    .S(_12474_),
    .Z(_00908_));
 NOR2_X1 _35206_ (.A1(_12339_),
    .A2(_00375_),
    .ZN(_12535_));
 MUX2_X1 _35207_ (.A(\core.keymem.key_mem[0][4] ),
    .B(_12535_),
    .S(_12474_),
    .Z(_00909_));
 INV_X1 _35208_ (.A(_00059_),
    .ZN(_12536_));
 NAND3_X1 _35209_ (.A1(_12230_),
    .A2(_12536_),
    .A3(_12236_),
    .ZN(_12537_));
 INV_X1 _35210_ (.A(\core.keymem.key_mem[0][50] ),
    .ZN(_12538_));
 OAI21_X1 _35211_ (.A(_12537_),
    .B1(_12238_),
    .B2(_12538_),
    .ZN(_00910_));
 NOR2_X1 _35212_ (.A1(_12339_),
    .A2(_00060_),
    .ZN(_12539_));
 MUX2_X1 _35213_ (.A(\core.keymem.key_mem[0][51] ),
    .B(_12539_),
    .S(_12474_),
    .Z(_00911_));
 BUF_X4 _35214_ (.A(_11801_),
    .Z(_12540_));
 NAND2_X1 _35215_ (.A1(\core.keymem.key_mem[0][52] ),
    .A2(_12540_),
    .ZN(_12541_));
 NOR2_X1 _35216_ (.A1(_00061_),
    .A2(_11862_),
    .ZN(_12542_));
 AOI21_X1 _35217_ (.A(_12542_),
    .B1(_12269_),
    .B2(\core.key[52] ),
    .ZN(_12543_));
 XOR2_X2 _35218_ (.A(\core.keymem.prev_key1_reg[84] ),
    .B(\core.keymem.prev_key1_reg[116] ),
    .Z(_12544_));
 XNOR2_X2 _35219_ (.A(_12073_),
    .B(_12544_),
    .ZN(_12545_));
 XNOR2_X2 _35220_ (.A(\core.keymem.prev_key1_reg[52] ),
    .B(_12545_),
    .ZN(_12546_));
 OAI21_X2 _35221_ (.A(_12543_),
    .B1(_12546_),
    .B2(_12001_),
    .ZN(_12547_));
 CLKBUF_X2 _35222_ (.A(\core.keymem.prev_key0_reg[52] ),
    .Z(_12548_));
 CLKBUF_X2 _35223_ (.A(\core.keymem.prev_key0_reg[84] ),
    .Z(_12549_));
 INV_X1 _35224_ (.A(_12549_),
    .ZN(_12550_));
 NAND2_X1 _35225_ (.A1(_12548_),
    .A2(_12550_),
    .ZN(_12551_));
 INV_X1 _35226_ (.A(_12548_),
    .ZN(_12552_));
 NAND2_X1 _35227_ (.A1(_12552_),
    .A2(_12549_),
    .ZN(_12553_));
 AOI221_X2 _35228_ (.A(_12061_),
    .B1(_12066_),
    .B2(_12067_),
    .C1(_12551_),
    .C2(_12553_),
    .ZN(_12554_));
 NAND2_X1 _35229_ (.A1(_12552_),
    .A2(_12550_),
    .ZN(_12555_));
 NAND2_X1 _35230_ (.A1(_12548_),
    .A2(_12549_),
    .ZN(_12556_));
 AOI221_X2 _35231_ (.A(_12062_),
    .B1(_12066_),
    .B2(_12067_),
    .C1(_12555_),
    .C2(_12556_),
    .ZN(_12557_));
 NOR3_X2 _35232_ (.A1(_12063_),
    .A2(_07828_),
    .A3(_07891_),
    .ZN(_12558_));
 NAND3_X1 _35233_ (.A1(_12552_),
    .A2(_12550_),
    .A3(_12062_),
    .ZN(_12559_));
 OR2_X1 _35234_ (.A1(_12061_),
    .A2(_12556_),
    .ZN(_12560_));
 NOR2_X1 _35235_ (.A1(_09027_),
    .A2(_09058_),
    .ZN(_12561_));
 AOI221_X2 _35236_ (.A(_12558_),
    .B1(_12559_),
    .B2(_12560_),
    .C1(_12561_),
    .C2(_12040_),
    .ZN(_12562_));
 NAND3_X1 _35237_ (.A1(_12548_),
    .A2(_12550_),
    .A3(_12061_),
    .ZN(_12563_));
 NAND3_X1 _35238_ (.A1(_12552_),
    .A2(_12549_),
    .A3(_12061_),
    .ZN(_12564_));
 AOI221_X2 _35239_ (.A(_12558_),
    .B1(_12563_),
    .B2(_12564_),
    .C1(_12561_),
    .C2(_12040_),
    .ZN(_12565_));
 OR4_X4 _35240_ (.A1(_12554_),
    .A2(_12557_),
    .A3(_12562_),
    .A4(_12565_),
    .ZN(_12566_));
 AOI21_X4 _35241_ (.A(_12547_),
    .B1(_12566_),
    .B2(_12311_),
    .ZN(_12567_));
 CLKBUF_X3 _35242_ (.A(_12567_),
    .Z(_12568_));
 OAI21_X1 _35243_ (.A(_12541_),
    .B1(_12568_),
    .B2(_12533_),
    .ZN(_00912_));
 NAND2_X1 _35244_ (.A1(\core.keymem.key_mem[0][53] ),
    .A2(_12540_),
    .ZN(_12569_));
 OAI21_X2 _35245_ (.A(_11823_),
    .B1(_11900_),
    .B2(\core.key[53] ),
    .ZN(_12570_));
 MUX2_X2 _35246_ (.A(_08036_),
    .B(_09123_),
    .S(_12040_),
    .Z(_12571_));
 XNOR2_X2 _35247_ (.A(\core.keymem.prev_key0_reg[85] ),
    .B(\core.keymem.prev_key0_reg[117] ),
    .ZN(_12572_));
 XOR2_X2 _35248_ (.A(_12571_),
    .B(_12572_),
    .Z(_12573_));
 XOR2_X2 _35249_ (.A(\core.keymem.prev_key0_reg[53] ),
    .B(_12573_),
    .Z(_12574_));
 AOI21_X4 _35250_ (.A(_12570_),
    .B1(_12574_),
    .B2(_12333_),
    .ZN(_12575_));
 NOR2_X2 _35251_ (.A1(_00062_),
    .A2(_11863_),
    .ZN(_12576_));
 NOR3_X4 _35252_ (.A1(_07974_),
    .A2(_07982_),
    .A3(_08035_),
    .ZN(_12577_));
 XNOR2_X2 _35253_ (.A(\core.keymem.prev_key1_reg[117] ),
    .B(_12577_),
    .ZN(_12578_));
 BUF_X2 _35254_ (.A(\core.keymem.prev_key1_reg[85] ),
    .Z(_12579_));
 XNOR2_X1 _35255_ (.A(\core.keymem.prev_key1_reg[53] ),
    .B(_12579_),
    .ZN(_12580_));
 XNOR2_X2 _35256_ (.A(_12578_),
    .B(_12580_),
    .ZN(_12581_));
 AND2_X1 _35257_ (.A1(_11888_),
    .A2(_12581_),
    .ZN(_12582_));
 NOR3_X4 _35258_ (.A1(_12575_),
    .A2(_12576_),
    .A3(_12582_),
    .ZN(_12583_));
 BUF_X4 _35259_ (.A(_12583_),
    .Z(_12584_));
 OAI21_X1 _35260_ (.A(_12569_),
    .B1(_12584_),
    .B2(_12533_),
    .ZN(_00913_));
 NOR2_X1 _35261_ (.A1(_12339_),
    .A2(_00063_),
    .ZN(_12585_));
 MUX2_X1 _35262_ (.A(\core.keymem.key_mem[0][54] ),
    .B(_12585_),
    .S(_12474_),
    .Z(_00914_));
 BUF_X4 _35263_ (.A(_11805_),
    .Z(_12586_));
 NOR2_X1 _35264_ (.A1(_12586_),
    .A2(_00064_),
    .ZN(_12587_));
 MUX2_X1 _35265_ (.A(\core.keymem.key_mem[0][55] ),
    .B(_12587_),
    .S(_12474_),
    .Z(_00915_));
 INV_X1 _35266_ (.A(_00065_),
    .ZN(_12588_));
 NAND3_X1 _35267_ (.A1(_12230_),
    .A2(_12588_),
    .A3(_12236_),
    .ZN(_12589_));
 INV_X1 _35268_ (.A(\core.keymem.key_mem[0][56] ),
    .ZN(_12590_));
 OAI21_X1 _35269_ (.A(_12589_),
    .B1(_12238_),
    .B2(_12590_),
    .ZN(_00916_));
 NOR2_X1 _35270_ (.A1(_12586_),
    .A2(_00067_),
    .ZN(_12591_));
 MUX2_X1 _35271_ (.A(\core.keymem.key_mem[0][57] ),
    .B(_12591_),
    .S(_12474_),
    .Z(_00917_));
 NOR2_X1 _35272_ (.A1(_12586_),
    .A2(_00069_),
    .ZN(_12592_));
 BUF_X4 _35273_ (.A(_11877_),
    .Z(_12593_));
 MUX2_X1 _35274_ (.A(\core.keymem.key_mem[0][58] ),
    .B(_12592_),
    .S(_12593_),
    .Z(_00918_));
 NOR2_X1 _35275_ (.A1(_12586_),
    .A2(_00071_),
    .ZN(_12594_));
 MUX2_X1 _35276_ (.A(\core.keymem.key_mem[0][59] ),
    .B(_12594_),
    .S(_12593_),
    .Z(_00919_));
 XNOR2_X1 _35277_ (.A(\core.keymem.prev_key1_reg[5] ),
    .B(_00377_),
    .ZN(_12595_));
 XNOR2_X1 _35278_ (.A(_12435_),
    .B(_12595_),
    .ZN(_12596_));
 XNOR2_X1 _35279_ (.A(_10075_),
    .B(_12596_),
    .ZN(_12597_));
 AND2_X1 _35280_ (.A1(_11888_),
    .A2(_12597_),
    .ZN(_12598_));
 AOI21_X1 _35281_ (.A(_11987_),
    .B1(_12092_),
    .B2(\core.key[5] ),
    .ZN(_12599_));
 XNOR2_X1 _35282_ (.A(\core.keymem.prev_key0_reg[69] ),
    .B(\core.keymem.prev_key0_reg[101] ),
    .ZN(_12600_));
 XNOR2_X1 _35283_ (.A(\core.keymem.prev_key0_reg[5] ),
    .B(\core.keymem.prev_key0_reg[37] ),
    .ZN(_12601_));
 XNOR2_X1 _35284_ (.A(_12600_),
    .B(_12601_),
    .ZN(_12602_));
 XNOR2_X1 _35285_ (.A(net10),
    .B(_12602_),
    .ZN(_12603_));
 OR2_X1 _35286_ (.A1(_11988_),
    .A2(_12603_),
    .ZN(_12604_));
 AOI221_X2 _35287_ (.A(_12598_),
    .B1(_12599_),
    .B2(_12604_),
    .C1(_00376_),
    .C2(_11842_),
    .ZN(_12605_));
 BUF_X2 _35288_ (.A(_12605_),
    .Z(_12606_));
 AOI22_X1 _35289_ (.A1(\core.keymem.key_mem[0][5] ),
    .A2(_11802_),
    .B1(_11806_),
    .B2(_12606_),
    .ZN(_12607_));
 INV_X1 _35290_ (.A(_12607_),
    .ZN(_00920_));
 NOR2_X1 _35291_ (.A1(_12586_),
    .A2(_00073_),
    .ZN(_12608_));
 MUX2_X1 _35292_ (.A(\core.keymem.key_mem[0][60] ),
    .B(_12608_),
    .S(_12593_),
    .Z(_00921_));
 NOR2_X1 _35293_ (.A1(_12586_),
    .A2(_00075_),
    .ZN(_12609_));
 MUX2_X1 _35294_ (.A(\core.keymem.key_mem[0][61] ),
    .B(_12609_),
    .S(_12593_),
    .Z(_00922_));
 INV_X1 _35295_ (.A(_00077_),
    .ZN(_12610_));
 NAND3_X1 _35296_ (.A1(_12230_),
    .A2(_12610_),
    .A3(_12236_),
    .ZN(_12611_));
 INV_X1 _35297_ (.A(\core.keymem.key_mem[0][62] ),
    .ZN(_12612_));
 OAI21_X1 _35298_ (.A(_12611_),
    .B1(_12238_),
    .B2(_12612_),
    .ZN(_00923_));
 NOR2_X1 _35299_ (.A1(_12586_),
    .A2(_00079_),
    .ZN(_12613_));
 MUX2_X1 _35300_ (.A(\core.keymem.key_mem[0][63] ),
    .B(_12613_),
    .S(_12593_),
    .Z(_00924_));
 AND2_X1 _35301_ (.A1(_00081_),
    .A2(_11841_),
    .ZN(_12614_));
 INV_X1 _35302_ (.A(\core.keymem.prev_key1_reg[64] ),
    .ZN(_12615_));
 XNOR2_X1 _35303_ (.A(_12615_),
    .B(_12351_),
    .ZN(_12616_));
 NOR2_X1 _35304_ (.A1(_11841_),
    .A2(_12616_),
    .ZN(_12617_));
 OR2_X1 _35305_ (.A1(\core.key[64] ),
    .A2(_12044_),
    .ZN(_12618_));
 XOR2_X1 _35306_ (.A(\core.keymem.prev_key0_reg[64] ),
    .B(_11835_),
    .Z(_12619_));
 OAI21_X1 _35307_ (.A(_12618_),
    .B1(_12619_),
    .B2(_12101_),
    .ZN(_12620_));
 AOI221_X2 _35308_ (.A(_12614_),
    .B1(_12617_),
    .B2(_11916_),
    .C1(_12620_),
    .C2(_12098_),
    .ZN(_12621_));
 BUF_X2 _35309_ (.A(_12621_),
    .Z(_12622_));
 AOI22_X1 _35310_ (.A1(\core.keymem.key_mem[0][64] ),
    .A2(_11802_),
    .B1(_11806_),
    .B2(_12622_),
    .ZN(_12623_));
 INV_X1 _35311_ (.A(_12623_),
    .ZN(_00925_));
 NOR2_X1 _35312_ (.A1(_12586_),
    .A2(_00082_),
    .ZN(_12624_));
 MUX2_X1 _35313_ (.A(\core.keymem.key_mem[0][65] ),
    .B(_12624_),
    .S(_12593_),
    .Z(_00926_));
 NOR2_X1 _35314_ (.A1(_12586_),
    .A2(_00083_),
    .ZN(_12625_));
 MUX2_X1 _35315_ (.A(\core.keymem.key_mem[0][66] ),
    .B(_12625_),
    .S(_12593_),
    .Z(_00927_));
 NOR2_X1 _35316_ (.A1(_12586_),
    .A2(_00084_),
    .ZN(_12626_));
 MUX2_X1 _35317_ (.A(\core.keymem.key_mem[0][67] ),
    .B(_12626_),
    .S(_12593_),
    .Z(_00928_));
 NAND2_X1 _35318_ (.A1(\core.keymem.key_mem[0][68] ),
    .A2(_12540_),
    .ZN(_12627_));
 AOI22_X2 _35319_ (.A1(_00085_),
    .A2(_12193_),
    .B1(_11889_),
    .B2(_12416_),
    .ZN(_12628_));
 BUF_X4 _35320_ (.A(_11892_),
    .Z(_12629_));
 NAND2_X1 _35321_ (.A1(\core.key[68] ),
    .A2(_12629_),
    .ZN(_12630_));
 NAND2_X1 _35322_ (.A1(_11936_),
    .A2(_12630_),
    .ZN(_12631_));
 XNOR2_X2 _35323_ (.A(_11858_),
    .B(_12418_),
    .ZN(_12632_));
 NOR2_X2 _35324_ (.A1(_12172_),
    .A2(_12632_),
    .ZN(_12633_));
 OAI21_X4 _35325_ (.A(_12628_),
    .B1(_12631_),
    .B2(_12633_),
    .ZN(_12634_));
 CLKBUF_X3 _35326_ (.A(_12634_),
    .Z(_12635_));
 OAI21_X1 _35327_ (.A(_12627_),
    .B1(_12635_),
    .B2(_12533_),
    .ZN(_00929_));
 BUF_X4 _35328_ (.A(_11805_),
    .Z(_12636_));
 NOR2_X1 _35329_ (.A1(_12636_),
    .A2(_00086_),
    .ZN(_12637_));
 MUX2_X1 _35330_ (.A(\core.keymem.key_mem[0][69] ),
    .B(_12637_),
    .S(_12593_),
    .Z(_00930_));
 CLKBUF_X3 _35331_ (.A(_11805_),
    .Z(_12638_));
 NAND2_X1 _35332_ (.A1(_12638_),
    .A2(_11877_),
    .ZN(_12639_));
 OAI21_X1 _35333_ (.A(_12639_),
    .B1(_11878_),
    .B2(\core.keymem.key_mem[0][6] ),
    .ZN(_12640_));
 AOI21_X1 _35334_ (.A(_12640_),
    .B1(_11883_),
    .B2(_00378_),
    .ZN(_00931_));
 NAND2_X1 _35335_ (.A1(\core.keymem.key_mem[0][70] ),
    .A2(_12540_),
    .ZN(_12641_));
 NOR2_X1 _35336_ (.A1(_00087_),
    .A2(_11862_),
    .ZN(_12642_));
 XOR2_X2 _35337_ (.A(_12464_),
    .B(_11887_),
    .Z(_12643_));
 AND2_X1 _35338_ (.A1(\core.key[70] ),
    .A2(_11820_),
    .ZN(_12644_));
 AOI221_X2 _35339_ (.A(_12642_),
    .B1(_12643_),
    .B2(_11888_),
    .C1(_12098_),
    .C2(_12644_),
    .ZN(_12645_));
 XNOR2_X2 _35340_ (.A(_12444_),
    .B(_11899_),
    .ZN(_12646_));
 NAND2_X1 _35341_ (.A1(_12311_),
    .A2(_12646_),
    .ZN(_12647_));
 AND2_X1 _35342_ (.A1(_12645_),
    .A2(_12647_),
    .ZN(_12648_));
 OAI21_X1 _35343_ (.A(_12641_),
    .B1(_12648_),
    .B2(_12533_),
    .ZN(_00932_));
 NAND2_X1 _35344_ (.A1(\core.keymem.key_mem[0][71] ),
    .A2(_12540_),
    .ZN(_12649_));
 NAND2_X1 _35345_ (.A1(_00088_),
    .A2(_12193_),
    .ZN(_12650_));
 NAND2_X1 _35346_ (.A1(\core.key[71] ),
    .A2(_12092_),
    .ZN(_12651_));
 NAND2_X1 _35347_ (.A1(_12098_),
    .A2(_12651_),
    .ZN(_12652_));
 BUF_X2 _35348_ (.A(\core.keymem.prev_key0_reg[71] ),
    .Z(_12653_));
 XNOR2_X2 _35349_ (.A(_12653_),
    .B(_11924_),
    .ZN(_12654_));
 NOR2_X1 _35350_ (.A1(_12629_),
    .A2(_12654_),
    .ZN(_12655_));
 XNOR2_X1 _35351_ (.A(\core.keymem.prev_key1_reg[71] ),
    .B(\core.keymem.prev_key1_reg[103] ),
    .ZN(_12656_));
 XNOR2_X2 _35352_ (.A(_11910_),
    .B(_12656_),
    .ZN(_12657_));
 OAI221_X2 _35353_ (.A(_12650_),
    .B1(_12652_),
    .B2(_12655_),
    .C1(_12263_),
    .C2(_12657_),
    .ZN(_12658_));
 CLKBUF_X3 _35354_ (.A(_12658_),
    .Z(_12659_));
 OAI21_X1 _35355_ (.A(_12649_),
    .B1(_12659_),
    .B2(_12533_),
    .ZN(_00933_));
 NAND2_X1 _35356_ (.A1(\core.keymem.key_mem[0][72] ),
    .A2(_12540_),
    .ZN(_12660_));
 NOR2_X1 _35357_ (.A1(_00089_),
    .A2(_11862_),
    .ZN(_12661_));
 AOI21_X1 _35358_ (.A(_12661_),
    .B1(_12269_),
    .B2(\core.key[72] ),
    .ZN(_12662_));
 XNOR2_X2 _35359_ (.A(\core.keymem.prev_key1_reg[104] ),
    .B(_07222_),
    .ZN(_12663_));
 XNOR2_X2 _35360_ (.A(\core.keymem.prev_key1_reg[72] ),
    .B(_12663_),
    .ZN(_12664_));
 OAI21_X2 _35361_ (.A(_12662_),
    .B1(_12664_),
    .B2(_12001_),
    .ZN(_12665_));
 CLKBUF_X3 _35362_ (.A(\core.keymem.prev_key0_reg[72] ),
    .Z(_12666_));
 BUF_X2 _35363_ (.A(\core.keymem.prev_key0_reg[104] ),
    .Z(_12667_));
 NOR2_X1 _35364_ (.A1(_07974_),
    .A2(_07982_),
    .ZN(_12668_));
 NOR2_X1 _35365_ (.A1(_11857_),
    .A2(_10612_),
    .ZN(_12669_));
 AOI22_X4 _35366_ (.A1(_11920_),
    .A2(_07222_),
    .B1(_12668_),
    .B2(_12669_),
    .ZN(_12670_));
 XNOR2_X2 _35367_ (.A(_12667_),
    .B(_12670_),
    .ZN(_12671_));
 XNOR2_X2 _35368_ (.A(_12666_),
    .B(_12671_),
    .ZN(_12672_));
 AOI21_X4 _35369_ (.A(_12665_),
    .B1(_12672_),
    .B2(_12311_),
    .ZN(_12673_));
 OR2_X1 _35370_ (.A1(_12183_),
    .A2(_12673_),
    .ZN(_12674_));
 OAI21_X1 _35371_ (.A(_12660_),
    .B1(_12674_),
    .B2(_12005_),
    .ZN(_00934_));
 NAND2_X1 _35372_ (.A1(\core.keymem.key_mem[0][73] ),
    .A2(_12540_),
    .ZN(_12675_));
 OR4_X1 _35373_ (.A1(_11830_),
    .A2(_08946_),
    .A3(_08966_),
    .A4(_08994_),
    .ZN(_12676_));
 OAI33_X1 _35374_ (.A1(_11857_),
    .A2(_07974_),
    .A3(_10668_),
    .B1(_12676_),
    .B2(_08916_),
    .B3(_07044_),
    .ZN(_12677_));
 XOR2_X2 _35375_ (.A(\core.keymem.prev_key0_reg[105] ),
    .B(net9),
    .Z(_12678_));
 XNOR2_X2 _35376_ (.A(\core.keymem.prev_key0_reg[73] ),
    .B(_12678_),
    .ZN(_12679_));
 BUF_X8 _35377_ (.A(_11798_),
    .Z(_12680_));
 NAND2_X1 _35378_ (.A1(_00090_),
    .A2(_12680_),
    .ZN(_12681_));
 NAND2_X1 _35379_ (.A1(_11908_),
    .A2(\core.key[73] ),
    .ZN(_12682_));
 BUF_X1 _35380_ (.A(\core.keymem.prev_key1_reg[73] ),
    .Z(_12683_));
 XOR2_X2 _35381_ (.A(\core.keymem.prev_key1_reg[105] ),
    .B(_08996_),
    .Z(_12684_));
 XNOR2_X1 _35382_ (.A(_12683_),
    .B(_12684_),
    .ZN(_12685_));
 OAI221_X2 _35383_ (.A(_11917_),
    .B1(_12099_),
    .B2(_12682_),
    .C1(_12685_),
    .C2(_12349_),
    .ZN(_12686_));
 AOI22_X4 _35384_ (.A1(_12311_),
    .A2(_12679_),
    .B1(_12681_),
    .B2(_12686_),
    .ZN(_12687_));
 CLKBUF_X3 _35385_ (.A(_12687_),
    .Z(_12688_));
 OAI21_X1 _35386_ (.A(_12675_),
    .B1(_12688_),
    .B2(_12533_),
    .ZN(_00935_));
 INV_X1 _35387_ (.A(_00091_),
    .ZN(_12689_));
 NAND3_X1 _35388_ (.A1(_12230_),
    .A2(_12689_),
    .A3(_12236_),
    .ZN(_12690_));
 INV_X1 _35389_ (.A(\core.keymem.key_mem[0][74] ),
    .ZN(_12691_));
 OAI21_X1 _35390_ (.A(_12690_),
    .B1(_12238_),
    .B2(_12691_),
    .ZN(_00936_));
 NOR2_X1 _35391_ (.A1(_12636_),
    .A2(_00092_),
    .ZN(_12692_));
 MUX2_X1 _35392_ (.A(\core.keymem.key_mem[0][75] ),
    .B(_12692_),
    .S(_12593_),
    .Z(_00937_));
 NOR2_X1 _35393_ (.A1(_12636_),
    .A2(_00093_),
    .ZN(_12693_));
 BUF_X4 _35394_ (.A(_11877_),
    .Z(_12694_));
 MUX2_X1 _35395_ (.A(\core.keymem.key_mem[0][76] ),
    .B(_12693_),
    .S(_12694_),
    .Z(_00938_));
 NOR2_X1 _35396_ (.A1(_12636_),
    .A2(_00094_),
    .ZN(_12695_));
 MUX2_X1 _35397_ (.A(\core.keymem.key_mem[0][77] ),
    .B(_12695_),
    .S(_12694_),
    .Z(_00939_));
 NAND2_X1 _35398_ (.A1(\core.keymem.key_mem[0][78] ),
    .A2(_12540_),
    .ZN(_12696_));
 AOI21_X1 _35399_ (.A(_11987_),
    .B1(_12629_),
    .B2(\core.key[78] ),
    .ZN(_12697_));
 BUF_X2 _35400_ (.A(\core.keymem.prev_key0_reg[78] ),
    .Z(_12698_));
 XNOR2_X1 _35401_ (.A(_12698_),
    .B(_11996_),
    .ZN(_12699_));
 OAI21_X1 _35402_ (.A(_12697_),
    .B1(_12699_),
    .B2(_12172_),
    .ZN(_12700_));
 BUF_X2 _35403_ (.A(\core.keymem.prev_key1_reg[78] ),
    .Z(_12701_));
 INV_X2 _35404_ (.A(_12701_),
    .ZN(_12702_));
 XNOR2_X2 _35405_ (.A(_11999_),
    .B(_10526_),
    .ZN(_12703_));
 XNOR2_X2 _35406_ (.A(_12702_),
    .B(_12703_),
    .ZN(_12704_));
 BUF_X8 _35407_ (.A(_11814_),
    .Z(_12705_));
 INV_X1 _35408_ (.A(_00095_),
    .ZN(_12706_));
 OAI221_X2 _35409_ (.A(_12700_),
    .B1(_12704_),
    .B2(_12705_),
    .C1(_12706_),
    .C2(_12035_),
    .ZN(_12707_));
 CLKBUF_X3 _35410_ (.A(_12707_),
    .Z(_12708_));
 OAI21_X1 _35411_ (.A(_12696_),
    .B1(_12708_),
    .B2(_12533_),
    .ZN(_00940_));
 NOR2_X1 _35412_ (.A1(_12636_),
    .A2(_00096_),
    .ZN(_12709_));
 MUX2_X1 _35413_ (.A(\core.keymem.key_mem[0][79] ),
    .B(_12709_),
    .S(_12694_),
    .Z(_00941_));
 NOR2_X1 _35414_ (.A1(_12636_),
    .A2(_00380_),
    .ZN(_12710_));
 MUX2_X1 _35415_ (.A(\core.keymem.key_mem[0][7] ),
    .B(_12710_),
    .S(_12694_),
    .Z(_00942_));
 NAND2_X1 _35416_ (.A1(\core.keymem.key_mem[0][80] ),
    .A2(_12540_),
    .ZN(_12711_));
 OAI22_X4 _35417_ (.A1(_00097_),
    .A2(_11917_),
    .B1(_12001_),
    .B2(_12528_),
    .ZN(_12712_));
 NAND2_X1 _35418_ (.A1(_12311_),
    .A2(_12522_),
    .ZN(_12713_));
 NAND3_X1 _35419_ (.A1(\core.key[80] ),
    .A2(_12101_),
    .A3(_11823_),
    .ZN(_12714_));
 NAND2_X2 _35420_ (.A1(_12713_),
    .A2(_12714_),
    .ZN(_12715_));
 NOR2_X4 _35421_ (.A1(_12712_),
    .A2(_12715_),
    .ZN(_12716_));
 OAI21_X1 _35422_ (.A(_12711_),
    .B1(_12716_),
    .B2(_12533_),
    .ZN(_00943_));
 NOR2_X1 _35423_ (.A1(_12636_),
    .A2(_00098_),
    .ZN(_12717_));
 MUX2_X1 _35424_ (.A(\core.keymem.key_mem[0][81] ),
    .B(_12717_),
    .S(_12694_),
    .Z(_00944_));
 NOR2_X1 _35425_ (.A1(_12636_),
    .A2(_00099_),
    .ZN(_12718_));
 MUX2_X1 _35426_ (.A(\core.keymem.key_mem[0][82] ),
    .B(_12718_),
    .S(_12694_),
    .Z(_00945_));
 NOR2_X1 _35427_ (.A1(_12636_),
    .A2(_00100_),
    .ZN(_12719_));
 MUX2_X1 _35428_ (.A(\core.keymem.key_mem[0][83] ),
    .B(_12719_),
    .S(_12694_),
    .Z(_00946_));
 NAND2_X1 _35429_ (.A1(\core.keymem.key_mem[0][84] ),
    .A2(_12540_),
    .ZN(_12720_));
 NOR2_X2 _35430_ (.A1(_00101_),
    .A2(_11863_),
    .ZN(_12721_));
 XNOR2_X1 _35431_ (.A(_12549_),
    .B(_12069_),
    .ZN(_12722_));
 MUX2_X1 _35432_ (.A(\core.key[84] ),
    .B(_12722_),
    .S(_11900_),
    .Z(_12723_));
 AOI221_X2 _35433_ (.A(_12721_),
    .B1(_12545_),
    .B2(_12027_),
    .C1(_11936_),
    .C2(_12723_),
    .ZN(_12724_));
 CLKBUF_X3 _35434_ (.A(_12724_),
    .Z(_12725_));
 OAI21_X1 _35435_ (.A(_12720_),
    .B1(_12725_),
    .B2(_12533_),
    .ZN(_00947_));
 NOR2_X1 _35436_ (.A1(_12636_),
    .A2(_00102_),
    .ZN(_12726_));
 MUX2_X1 _35437_ (.A(\core.keymem.key_mem[0][85] ),
    .B(_12726_),
    .S(_12694_),
    .Z(_00948_));
 BUF_X2 _35438_ (.A(\core.keymem.prev_key1_reg[86] ),
    .Z(_12727_));
 XOR2_X2 _35439_ (.A(\core.keymem.prev_key1_reg[118] ),
    .B(_08101_),
    .Z(_12728_));
 XOR2_X2 _35440_ (.A(_12727_),
    .B(_12728_),
    .Z(_12729_));
 NOR2_X1 _35441_ (.A1(_11814_),
    .A2(_12729_),
    .ZN(_12730_));
 AOI21_X1 _35442_ (.A(_11987_),
    .B1(_12092_),
    .B2(\core.key[86] ),
    .ZN(_12731_));
 CLKBUF_X3 _35443_ (.A(\core.keymem.prev_key0_reg[86] ),
    .Z(_12732_));
 INV_X1 _35444_ (.A(\core.keymem.prev_key0_reg[118] ),
    .ZN(_12733_));
 NAND3_X1 _35445_ (.A1(_11850_),
    .A2(_08085_),
    .A3(_08099_),
    .ZN(_12734_));
 NAND2_X1 _35446_ (.A1(_08070_),
    .A2(_08078_),
    .ZN(_12735_));
 OAI33_X1 _35447_ (.A1(_11856_),
    .A2(_08483_),
    .A3(_09170_),
    .B1(_12734_),
    .B2(_12735_),
    .B3(_07974_),
    .ZN(_12736_));
 XNOR2_X2 _35448_ (.A(_12733_),
    .B(_12736_),
    .ZN(_12737_));
 XOR2_X2 _35449_ (.A(_12732_),
    .B(_12737_),
    .Z(_12738_));
 OR2_X1 _35450_ (.A1(_11988_),
    .A2(_12738_),
    .ZN(_12739_));
 AOI221_X2 _35451_ (.A(_12730_),
    .B1(_12731_),
    .B2(_12739_),
    .C1(_00103_),
    .C2(_11842_),
    .ZN(_12740_));
 BUF_X4 _35452_ (.A(_12740_),
    .Z(_12741_));
 AOI22_X1 _35453_ (.A1(\core.keymem.key_mem[0][86] ),
    .A2(_11802_),
    .B1(_11806_),
    .B2(_12741_),
    .ZN(_12742_));
 INV_X1 _35454_ (.A(_12742_),
    .ZN(_00949_));
 NOR2_X1 _35455_ (.A1(_12638_),
    .A2(_00104_),
    .ZN(_12743_));
 MUX2_X1 _35456_ (.A(\core.keymem.key_mem[0][87] ),
    .B(_12743_),
    .S(_12694_),
    .Z(_00950_));
 NOR2_X1 _35457_ (.A1(_12638_),
    .A2(_00105_),
    .ZN(_12744_));
 MUX2_X1 _35458_ (.A(\core.keymem.key_mem[0][88] ),
    .B(_12744_),
    .S(_12694_),
    .Z(_00951_));
 NOR2_X1 _35459_ (.A1(_12638_),
    .A2(_00107_),
    .ZN(_12745_));
 MUX2_X1 _35460_ (.A(\core.keymem.key_mem[0][89] ),
    .B(_12745_),
    .S(_11882_),
    .Z(_00952_));
 INV_X1 _35461_ (.A(_00381_),
    .ZN(_12746_));
 NAND3_X1 _35462_ (.A1(_12230_),
    .A2(_12746_),
    .A3(_12236_),
    .ZN(_12747_));
 INV_X1 _35463_ (.A(\core.keymem.key_mem[0][8] ),
    .ZN(_12748_));
 OAI21_X1 _35464_ (.A(_12747_),
    .B1(_12238_),
    .B2(_12748_),
    .ZN(_00953_));
 NOR2_X1 _35465_ (.A1(_12638_),
    .A2(_00109_),
    .ZN(_12749_));
 MUX2_X1 _35466_ (.A(\core.keymem.key_mem[0][90] ),
    .B(_12749_),
    .S(_11882_),
    .Z(_00954_));
 NOR2_X1 _35467_ (.A1(_12638_),
    .A2(_00111_),
    .ZN(_12750_));
 MUX2_X1 _35468_ (.A(\core.keymem.key_mem[0][91] ),
    .B(_12750_),
    .S(_11882_),
    .Z(_00955_));
 BUF_X4 _35469_ (.A(_11952_),
    .Z(_12751_));
 INV_X1 _35470_ (.A(_00113_),
    .ZN(_12752_));
 NAND3_X1 _35471_ (.A1(_12751_),
    .A2(_12752_),
    .A3(_12236_),
    .ZN(_12753_));
 INV_X1 _35472_ (.A(\core.keymem.key_mem[0][92] ),
    .ZN(_12754_));
 OAI21_X1 _35473_ (.A(_12753_),
    .B1(_12238_),
    .B2(_12754_),
    .ZN(_00956_));
 NOR2_X1 _35474_ (.A1(_12638_),
    .A2(_00115_),
    .ZN(_12755_));
 MUX2_X1 _35475_ (.A(\core.keymem.key_mem[0][93] ),
    .B(_12755_),
    .S(_11882_),
    .Z(_00957_));
 NOR2_X1 _35476_ (.A1(_12638_),
    .A2(_00117_),
    .ZN(_12756_));
 MUX2_X1 _35477_ (.A(\core.keymem.key_mem[0][94] ),
    .B(_12756_),
    .S(_11882_),
    .Z(_00958_));
 NOR2_X1 _35478_ (.A1(_12638_),
    .A2(_00119_),
    .ZN(_12757_));
 MUX2_X1 _35479_ (.A(\core.keymem.key_mem[0][95] ),
    .B(_12757_),
    .S(_11882_),
    .Z(_00959_));
 INV_X1 _35480_ (.A(_00121_),
    .ZN(_12758_));
 NAND3_X1 _35481_ (.A1(_12751_),
    .A2(_12758_),
    .A3(_11878_),
    .ZN(_12759_));
 INV_X1 _35482_ (.A(\core.keymem.key_mem[0][96] ),
    .ZN(_12760_));
 OAI21_X1 _35483_ (.A(_12759_),
    .B1(_11880_),
    .B2(_12760_),
    .ZN(_00960_));
 NAND2_X1 _35484_ (.A1(\core.keymem.key_mem[0][97] ),
    .A2(_11802_),
    .ZN(_12761_));
 NOR2_X2 _35485_ (.A1(_00122_),
    .A2(_11868_),
    .ZN(_12762_));
 AND2_X1 _35486_ (.A1(_11868_),
    .A2(_12358_),
    .ZN(_12763_));
 OR3_X1 _35487_ (.A1(_11908_),
    .A2(_12762_),
    .A3(_12763_),
    .ZN(_12764_));
 AND2_X1 _35488_ (.A1(_16229_),
    .A2(_12764_),
    .ZN(_12765_));
 NAND2_X2 _35489_ (.A1(_09707_),
    .A2(_09706_),
    .ZN(_12766_));
 NOR2_X1 _35490_ (.A1(_11829_),
    .A2(_09705_),
    .ZN(_12767_));
 AND4_X1 _35491_ (.A1(_09734_),
    .A2(_09753_),
    .A3(_09775_),
    .A4(_12767_),
    .ZN(_12768_));
 OR2_X1 _35492_ (.A1(_11850_),
    .A2(_08916_),
    .ZN(_12769_));
 NOR4_X4 _35493_ (.A1(_08946_),
    .A2(_08966_),
    .A3(_08994_),
    .A4(_12769_),
    .ZN(_12770_));
 AOI22_X4 _35494_ (.A1(_12766_),
    .A2(_12768_),
    .B1(_12770_),
    .B2(_08907_),
    .ZN(_12771_));
 XNOR2_X2 _35495_ (.A(\core.keymem.prev_key0_reg[97] ),
    .B(_12771_),
    .ZN(_12772_));
 NOR2_X1 _35496_ (.A1(_11988_),
    .A2(_12772_),
    .ZN(_12773_));
 AOI21_X1 _35497_ (.A(_12773_),
    .B1(_12101_),
    .B2(\core.key[97] ),
    .ZN(_12774_));
 OAI21_X2 _35498_ (.A(_12156_),
    .B1(_11842_),
    .B2(_12774_),
    .ZN(_12775_));
 OAI21_X4 _35499_ (.A(_12765_),
    .B1(_12775_),
    .B2(_12762_),
    .ZN(_12776_));
 CLKBUF_X3 _35500_ (.A(_12776_),
    .Z(_12777_));
 OAI21_X1 _35501_ (.A(_12761_),
    .B1(_12777_),
    .B2(_12005_),
    .ZN(_00961_));
 NAND2_X1 _35502_ (.A1(\core.keymem.key_mem[0][98] ),
    .A2(_11802_),
    .ZN(_12778_));
 BUF_X4 _35503_ (.A(_11799_),
    .Z(_12779_));
 NAND2_X2 _35504_ (.A1(_09808_),
    .A2(_09858_),
    .ZN(_12780_));
 XNOR2_X1 _35505_ (.A(_00124_),
    .B(_12780_),
    .ZN(_12781_));
 NOR2_X1 _35506_ (.A1(_11799_),
    .A2(_12781_),
    .ZN(_12782_));
 AOI22_X2 _35507_ (.A1(_00123_),
    .A2(_12779_),
    .B1(_12782_),
    .B2(_11847_),
    .ZN(_12783_));
 NAND2_X1 _35508_ (.A1(\core.key[98] ),
    .A2(_11989_),
    .ZN(_12784_));
 OAI21_X2 _35509_ (.A(_12784_),
    .B1(_12324_),
    .B2(_11997_),
    .ZN(_12785_));
 BUF_X4 _35510_ (.A(_11904_),
    .Z(_12786_));
 OAI21_X4 _35511_ (.A(_12783_),
    .B1(_12785_),
    .B2(_12786_),
    .ZN(_12787_));
 OR2_X1 _35512_ (.A1(_12183_),
    .A2(_12787_),
    .ZN(_12788_));
 OAI21_X1 _35513_ (.A(_12778_),
    .B1(_12788_),
    .B2(_12005_),
    .ZN(_00962_));
 XOR2_X1 _35514_ (.A(_00126_),
    .B(_09949_),
    .Z(_12789_));
 NOR2_X1 _35515_ (.A1(_11798_),
    .A2(_12789_),
    .ZN(_12790_));
 AOI21_X2 _35516_ (.A(_12790_),
    .B1(_11841_),
    .B2(_00125_),
    .ZN(_12791_));
 OAI21_X2 _35517_ (.A(_16228_),
    .B1(_11909_),
    .B2(_12791_),
    .ZN(_12792_));
 OR2_X1 _35518_ (.A1(_00125_),
    .A2(_11885_),
    .ZN(_12793_));
 NOR3_X1 _35519_ (.A1(_12385_),
    .A2(_12390_),
    .A3(_12391_),
    .ZN(_12794_));
 AOI21_X1 _35520_ (.A(_12393_),
    .B1(_12378_),
    .B2(_12381_),
    .ZN(_12795_));
 OR2_X1 _35521_ (.A1(_12794_),
    .A2(_12795_),
    .ZN(_12796_));
 MUX2_X1 _35522_ (.A(\core.key[99] ),
    .B(_12796_),
    .S(_11925_),
    .Z(_12797_));
 AOI21_X2 _35523_ (.A(_11916_),
    .B1(_11917_),
    .B2(_12797_),
    .ZN(_12798_));
 AOI21_X4 _35524_ (.A(_12792_),
    .B1(_12793_),
    .B2(_12798_),
    .ZN(_12799_));
 BUF_X2 _35525_ (.A(_12799_),
    .Z(_12800_));
 MUX2_X1 _35526_ (.A(\core.keymem.key_mem[0][99] ),
    .B(_12800_),
    .S(_11882_),
    .Z(_00963_));
 NOR2_X1 _35527_ (.A1(_12638_),
    .A2(_00404_),
    .ZN(_12801_));
 MUX2_X1 _35528_ (.A(\core.keymem.key_mem[0][9] ),
    .B(_12801_),
    .S(_11882_),
    .Z(_00964_));
 INV_X2 _35529_ (.A(_16218_),
    .ZN(_12802_));
 NAND2_X4 _35530_ (.A1(_11794_),
    .A2(_12802_),
    .ZN(_12803_));
 NAND2_X4 _35531_ (.A1(_16222_),
    .A2(_16216_),
    .ZN(_12804_));
 NOR2_X4 _35532_ (.A1(_12803_),
    .A2(_12804_),
    .ZN(_12805_));
 BUF_X4 _35533_ (.A(_12805_),
    .Z(_12806_));
 BUF_X4 _35534_ (.A(_12806_),
    .Z(_12807_));
 MUX2_X1 _35535_ (.A(\core.keymem.key_mem[10][0] ),
    .B(_11844_),
    .S(_12807_),
    .Z(_00965_));
 MUX2_X1 _35536_ (.A(\core.keymem.key_mem[10][100] ),
    .B(_11873_),
    .S(_12807_),
    .Z(_00966_));
 BUF_X4 _35537_ (.A(_11916_),
    .Z(_12808_));
 AOI21_X2 _35538_ (.A(_12779_),
    .B1(_12433_),
    .B2(_12808_),
    .ZN(_12809_));
 MUX2_X1 _35539_ (.A(\core.key[101] ),
    .B(_12428_),
    .S(_11828_),
    .Z(_12810_));
 INV_X1 _35540_ (.A(_12810_),
    .ZN(_12811_));
 OAI21_X4 _35541_ (.A(_12809_),
    .B1(_12811_),
    .B2(_12292_),
    .ZN(_12812_));
 BUF_X2 _35542_ (.A(_12812_),
    .Z(_12813_));
 MUX2_X1 _35543_ (.A(\core.keymem.key_mem[10][101] ),
    .B(_12813_),
    .S(_12807_),
    .Z(_00967_));
 MUX2_X1 _35544_ (.A(\core.keymem.key_mem[10][102] ),
    .B(_11906_),
    .S(_12807_),
    .Z(_00968_));
 MUX2_X1 _35545_ (.A(\core.keymem.key_mem[10][103] ),
    .B(_11929_),
    .S(_12807_),
    .Z(_00969_));
 OR2_X1 _35546_ (.A1(_12803_),
    .A2(_12804_),
    .ZN(_12814_));
 CLKBUF_X3 _35547_ (.A(_12814_),
    .Z(_12815_));
 BUF_X4 _35548_ (.A(_12815_),
    .Z(_12816_));
 NAND2_X1 _35549_ (.A1(\core.keymem.key_mem[10][104] ),
    .A2(_12816_),
    .ZN(_12817_));
 AND2_X1 _35550_ (.A1(_11846_),
    .A2(_12663_),
    .ZN(_12818_));
 NOR2_X1 _35551_ (.A1(\core.key[104] ),
    .A2(_11945_),
    .ZN(_12819_));
 AOI21_X2 _35552_ (.A(_12819_),
    .B1(_12671_),
    .B2(_12149_),
    .ZN(_12820_));
 AOI221_X2 _35553_ (.A(_12818_),
    .B1(_11812_),
    .B2(_11793_),
    .C1(_12156_),
    .C2(_12820_),
    .ZN(_12821_));
 BUF_X2 _35554_ (.A(_12821_),
    .Z(_12822_));
 BUF_X4 _35555_ (.A(_12815_),
    .Z(_12823_));
 BUF_X4 _35556_ (.A(_12823_),
    .Z(_12824_));
 OAI21_X1 _35557_ (.A(_12817_),
    .B1(_12822_),
    .B2(_12824_),
    .ZN(_00970_));
 AOI21_X2 _35558_ (.A(_12779_),
    .B1(_12684_),
    .B2(_11847_),
    .ZN(_12825_));
 XNOR2_X2 _35559_ (.A(\core.keymem.prev_key0_reg[105] ),
    .B(net9),
    .ZN(_12826_));
 MUX2_X1 _35560_ (.A(\core.key[105] ),
    .B(_12826_),
    .S(_11900_),
    .Z(_12827_));
 INV_X1 _35561_ (.A(_12827_),
    .ZN(_12828_));
 OAI21_X4 _35562_ (.A(_12825_),
    .B1(_12828_),
    .B2(_12292_),
    .ZN(_12829_));
 BUF_X2 _35563_ (.A(_12829_),
    .Z(_12830_));
 MUX2_X1 _35564_ (.A(\core.keymem.key_mem[10][105] ),
    .B(_12830_),
    .S(_12807_),
    .Z(_00971_));
 NAND2_X1 _35565_ (.A1(_11935_),
    .A2(_11950_),
    .ZN(_12831_));
 CLKBUF_X2 _35566_ (.A(_12831_),
    .Z(_12832_));
 BUF_X4 _35567_ (.A(_12806_),
    .Z(_12833_));
 MUX2_X1 _35568_ (.A(\core.keymem.key_mem[10][106] ),
    .B(_12832_),
    .S(_12833_),
    .Z(_00972_));
 MUX2_X1 _35569_ (.A(\core.keymem.key_mem[10][107] ),
    .B(_11967_),
    .S(_12833_),
    .Z(_00973_));
 MUX2_X1 _35570_ (.A(\core.keymem.key_mem[10][108] ),
    .B(_11981_),
    .S(_12833_),
    .Z(_00974_));
 BUF_X4 _35571_ (.A(_12347_),
    .Z(_12834_));
 BUF_X2 _35572_ (.A(\core.keymem.prev_key0_reg[109] ),
    .Z(_12835_));
 MUX2_X2 _35573_ (.A(_12577_),
    .B(_10469_),
    .S(_11920_),
    .Z(_12836_));
 XNOR2_X1 _35574_ (.A(_12835_),
    .B(_12836_),
    .ZN(_12837_));
 NOR2_X1 _35575_ (.A1(_12629_),
    .A2(_12837_),
    .ZN(_12838_));
 OAI21_X1 _35576_ (.A(_06677_),
    .B1(\core.key[109] ),
    .B2(_12333_),
    .ZN(_12839_));
 XOR2_X2 _35577_ (.A(\core.keymem.prev_key1_reg[109] ),
    .B(_10469_),
    .Z(_12840_));
 OAI221_X2 _35578_ (.A(_12834_),
    .B1(_12838_),
    .B2(_12839_),
    .C1(_12840_),
    .C2(_12301_),
    .ZN(_12841_));
 BUF_X2 _35579_ (.A(_12841_),
    .Z(_12842_));
 MUX2_X1 _35580_ (.A(\core.keymem.key_mem[10][109] ),
    .B(_12842_),
    .S(_12833_),
    .Z(_00975_));
 NAND2_X1 _35581_ (.A1(\core.keymem.key_mem[10][10] ),
    .A2(_12816_),
    .ZN(_12843_));
 BUF_X4 _35582_ (.A(_12333_),
    .Z(_12844_));
 BUF_X2 _35583_ (.A(\core.keymem.prev_key0_reg[42] ),
    .Z(_12845_));
 BUF_X2 _35584_ (.A(\core.keymem.prev_key0_reg[74] ),
    .Z(_12846_));
 XNOR2_X1 _35585_ (.A(_12845_),
    .B(_12846_),
    .ZN(_12847_));
 XNOR2_X1 _35586_ (.A(\core.keymem.prev_key0_reg[10] ),
    .B(_12847_),
    .ZN(_12848_));
 XOR2_X2 _35587_ (.A(_11944_),
    .B(_12848_),
    .Z(_12849_));
 AND2_X2 _35588_ (.A1(_12844_),
    .A2(_12849_),
    .ZN(_12850_));
 NAND2_X1 _35589_ (.A1(\core.key[10] ),
    .A2(_11997_),
    .ZN(_12851_));
 NAND2_X1 _35590_ (.A1(_12335_),
    .A2(_12851_),
    .ZN(_12852_));
 XNOR2_X1 _35591_ (.A(\core.keymem.prev_key1_reg[74] ),
    .B(\core.keymem.prev_key1_reg[106] ),
    .ZN(_12853_));
 XNOR2_X2 _35592_ (.A(_11947_),
    .B(_12853_),
    .ZN(_12854_));
 XOR2_X2 _35593_ (.A(\core.keymem.prev_key1_reg[42] ),
    .B(_12854_),
    .Z(_12855_));
 XNOR2_X2 _35594_ (.A(\core.keymem.prev_key1_reg[10] ),
    .B(_12855_),
    .ZN(_12856_));
 OAI22_X4 _35595_ (.A1(_12850_),
    .A2(_12852_),
    .B1(_12856_),
    .B2(_12263_),
    .ZN(_12857_));
 CLKBUF_X3 _35596_ (.A(_12857_),
    .Z(_12858_));
 OAI21_X1 _35597_ (.A(_12843_),
    .B1(_12858_),
    .B2(_12824_),
    .ZN(_00976_));
 CLKBUF_X2 _35598_ (.A(_12003_),
    .Z(_12859_));
 MUX2_X1 _35599_ (.A(\core.keymem.key_mem[10][110] ),
    .B(_12859_),
    .S(_12833_),
    .Z(_00977_));
 MUX2_X1 _35600_ (.A(\core.keymem.key_mem[10][111] ),
    .B(_12017_),
    .S(_12833_),
    .Z(_00978_));
 MUX2_X1 _35601_ (.A(\core.keymem.key_mem[10][112] ),
    .B(_12031_),
    .S(_12833_),
    .Z(_00979_));
 BUF_X4 _35602_ (.A(_11842_),
    .Z(_12860_));
 NOR2_X1 _35603_ (.A1(_08705_),
    .A2(_08715_),
    .ZN(_12861_));
 MUX2_X2 _35604_ (.A(_12861_),
    .B(_10669_),
    .S(_11920_),
    .Z(_12862_));
 XNOR2_X1 _35605_ (.A(\core.keymem.prev_key0_reg[113] ),
    .B(_12862_),
    .ZN(_12863_));
 MUX2_X1 _35606_ (.A(\core.key[113] ),
    .B(_12863_),
    .S(_11860_),
    .Z(_12864_));
 XNOR2_X2 _35607_ (.A(\core.keymem.prev_key1_reg[113] ),
    .B(_10669_),
    .ZN(_12865_));
 MUX2_X1 _35608_ (.A(_12864_),
    .B(_12865_),
    .S(_11846_),
    .Z(_12866_));
 OR2_X1 _35609_ (.A1(_12860_),
    .A2(_12866_),
    .ZN(_12867_));
 CLKBUF_X2 _35610_ (.A(_12867_),
    .Z(_12868_));
 MUX2_X1 _35611_ (.A(\core.keymem.key_mem[10][113] ),
    .B(_12868_),
    .S(_12833_),
    .Z(_00980_));
 CLKBUF_X2 _35612_ (.A(_12048_),
    .Z(_12869_));
 MUX2_X1 _35613_ (.A(\core.keymem.key_mem[10][114] ),
    .B(_12869_),
    .S(_12833_),
    .Z(_00981_));
 MUX2_X1 _35614_ (.A(\core.keymem.key_mem[10][115] ),
    .B(_12059_),
    .S(_12833_),
    .Z(_00982_));
 BUF_X4 _35615_ (.A(_12806_),
    .Z(_12870_));
 MUX2_X1 _35616_ (.A(\core.keymem.key_mem[10][116] ),
    .B(_12077_),
    .S(_12870_),
    .Z(_00983_));
 BUF_X8 _35617_ (.A(_12035_),
    .Z(_12871_));
 XOR2_X1 _35618_ (.A(\core.keymem.prev_key0_reg[117] ),
    .B(_12571_),
    .Z(_12872_));
 MUX2_X2 _35619_ (.A(\core.key[117] ),
    .B(_12872_),
    .S(_11828_),
    .Z(_12873_));
 NAND2_X2 _35620_ (.A1(_06678_),
    .A2(_12873_),
    .ZN(_12874_));
 NAND2_X2 _35621_ (.A1(_12292_),
    .A2(_12578_),
    .ZN(_12875_));
 NAND3_X4 _35622_ (.A1(_12871_),
    .A2(_12874_),
    .A3(_12875_),
    .ZN(_12876_));
 BUF_X2 _35623_ (.A(_12876_),
    .Z(_12877_));
 MUX2_X1 _35624_ (.A(\core.keymem.key_mem[10][117] ),
    .B(_12877_),
    .S(_12870_),
    .Z(_00984_));
 AOI21_X2 _35625_ (.A(_12779_),
    .B1(_12728_),
    .B2(_12808_),
    .ZN(_12878_));
 NAND2_X1 _35626_ (.A1(_11901_),
    .A2(_12737_),
    .ZN(_12879_));
 OAI21_X2 _35627_ (.A(_12879_),
    .B1(_12170_),
    .B2(\core.key[118] ),
    .ZN(_12880_));
 OAI21_X4 _35628_ (.A(_12878_),
    .B1(_12880_),
    .B2(_12292_),
    .ZN(_12881_));
 BUF_X2 _35629_ (.A(_12881_),
    .Z(_12882_));
 MUX2_X1 _35630_ (.A(\core.keymem.key_mem[10][118] ),
    .B(_12882_),
    .S(_12870_),
    .Z(_00985_));
 MUX2_X1 _35631_ (.A(\core.keymem.key_mem[10][119] ),
    .B(_12096_),
    .S(_12870_),
    .Z(_00986_));
 NAND2_X1 _35632_ (.A1(\core.keymem.key_mem[10][11] ),
    .A2(_12816_),
    .ZN(_12883_));
 BUF_X4 _35633_ (.A(_12705_),
    .Z(_12884_));
 XNOR2_X1 _35634_ (.A(\core.keymem.prev_key1_reg[75] ),
    .B(\core.keymem.prev_key1_reg[107] ),
    .ZN(_12885_));
 XNOR2_X2 _35635_ (.A(_10352_),
    .B(_12885_),
    .ZN(_12886_));
 XOR2_X2 _35636_ (.A(\core.keymem.prev_key1_reg[43] ),
    .B(_12886_),
    .Z(_12887_));
 XNOR2_X2 _35637_ (.A(\core.keymem.prev_key1_reg[11] ),
    .B(_12887_),
    .ZN(_12888_));
 XNOR2_X2 _35638_ (.A(\core.keymem.prev_key0_reg[75] ),
    .B(\core.keymem.prev_key0_reg[107] ),
    .ZN(_12889_));
 XNOR2_X1 _35639_ (.A(\core.keymem.prev_key0_reg[43] ),
    .B(_12889_),
    .ZN(_12890_));
 XOR2_X1 _35640_ (.A(\core.keymem.prev_key0_reg[11] ),
    .B(_12890_),
    .Z(_12891_));
 XNOR2_X1 _35641_ (.A(_11962_),
    .B(_12891_),
    .ZN(_12892_));
 MUX2_X2 _35642_ (.A(\core.key[11] ),
    .B(_12892_),
    .S(_12099_),
    .Z(_12893_));
 OAI22_X4 _35643_ (.A1(_12884_),
    .A2(_12888_),
    .B1(_12893_),
    .B2(_12786_),
    .ZN(_12894_));
 CLKBUF_X3 _35644_ (.A(_12894_),
    .Z(_12895_));
 BUF_X4 _35645_ (.A(_12823_),
    .Z(_12896_));
 OAI21_X1 _35646_ (.A(_12883_),
    .B1(_12895_),
    .B2(_12896_),
    .ZN(_00987_));
 MUX2_X1 _35647_ (.A(\core.keymem.key_mem[10][120] ),
    .B(_12124_),
    .S(_12870_),
    .Z(_00988_));
 MUX2_X1 _35648_ (.A(\core.keymem.key_mem[10][121] ),
    .B(_12160_),
    .S(_12870_),
    .Z(_00989_));
 NAND2_X1 _35649_ (.A1(_12162_),
    .A2(_11842_),
    .ZN(_12897_));
 MUX2_X2 _35650_ (.A(_12780_),
    .B(_12278_),
    .S(_12175_),
    .Z(_12898_));
 XNOR2_X1 _35651_ (.A(\core.keymem.prev_key0_reg[122] ),
    .B(_12898_),
    .ZN(_12899_));
 MUX2_X1 _35652_ (.A(_00162_),
    .B(_12899_),
    .S(_11945_),
    .Z(_12900_));
 XNOR2_X2 _35653_ (.A(\core.keymem.prev_key1_reg[122] ),
    .B(_12278_),
    .ZN(_12901_));
 OAI221_X2 _35654_ (.A(_12897_),
    .B1(_12900_),
    .B2(_11904_),
    .C1(_12901_),
    .C2(_12705_),
    .ZN(_12902_));
 BUF_X2 _35655_ (.A(_12902_),
    .Z(_12903_));
 MUX2_X1 _35656_ (.A(\core.keymem.key_mem[10][122] ),
    .B(_12903_),
    .S(_12870_),
    .Z(_00990_));
 NAND2_X1 _35657_ (.A1(\core.keymem.key_mem[10][123] ),
    .A2(_12816_),
    .ZN(_12904_));
 BUF_X4 _35658_ (.A(_12823_),
    .Z(_12905_));
 OAI21_X1 _35659_ (.A(_12904_),
    .B1(_12905_),
    .B2(_12182_),
    .ZN(_00991_));
 NAND2_X1 _35660_ (.A1(\core.keymem.key_mem[10][124] ),
    .A2(_12816_),
    .ZN(_12906_));
 NAND2_X1 _35661_ (.A1(_00165_),
    .A2(_12779_),
    .ZN(_12907_));
 BUF_X2 _35662_ (.A(\core.keymem.rcon_logic.tmp_rcon[5] ),
    .Z(_12908_));
 OAI21_X1 _35663_ (.A(_12908_),
    .B1(_09027_),
    .B2(_09058_),
    .ZN(_12909_));
 OR3_X1 _35664_ (.A1(_12908_),
    .A2(_09027_),
    .A3(_09058_),
    .ZN(_12910_));
 AND2_X2 _35665_ (.A1(_12909_),
    .A2(_12910_),
    .ZN(_12911_));
 XNOR2_X2 _35666_ (.A(\core.keymem.prev_key1_reg[124] ),
    .B(_12911_),
    .ZN(_12912_));
 NAND2_X1 _35667_ (.A1(_11875_),
    .A2(_12912_),
    .ZN(_12913_));
 INV_X1 _35668_ (.A(_00166_),
    .ZN(_12914_));
 INV_X2 _35669_ (.A(\core.keymem.prev_key0_reg[124] ),
    .ZN(_12915_));
 NAND4_X1 _35670_ (.A1(_12176_),
    .A2(_12915_),
    .A3(_12909_),
    .A4(_12910_),
    .ZN(_12916_));
 BUF_X4 _35671_ (.A(_11832_),
    .Z(_12917_));
 NAND2_X1 _35672_ (.A1(_12917_),
    .A2(_12915_),
    .ZN(_12918_));
 BUF_X2 _35673_ (.A(\core.keymem.prev_key0_reg[124] ),
    .Z(_12919_));
 NAND2_X1 _35674_ (.A1(_12917_),
    .A2(_12919_),
    .ZN(_12920_));
 MUX2_X1 _35675_ (.A(_12918_),
    .B(_12920_),
    .S(_10009_),
    .Z(_12921_));
 NAND2_X1 _35676_ (.A1(_12176_),
    .A2(_12919_),
    .ZN(_12922_));
 OAI211_X2 _35677_ (.A(_12916_),
    .B(_12921_),
    .C1(_12911_),
    .C2(_12922_),
    .ZN(_12923_));
 MUX2_X1 _35678_ (.A(_12914_),
    .B(_12923_),
    .S(_11900_),
    .Z(_12924_));
 OAI221_X2 _35679_ (.A(_12907_),
    .B1(_12913_),
    .B2(_12156_),
    .C1(_11904_),
    .C2(_12924_),
    .ZN(_12925_));
 BUF_X2 _35680_ (.A(_12925_),
    .Z(_12926_));
 OAI21_X1 _35681_ (.A(_12906_),
    .B1(_12905_),
    .B2(_12926_),
    .ZN(_00992_));
 NOR2_X1 _35682_ (.A1(_00168_),
    .A2(_11826_),
    .ZN(_12927_));
 OR2_X1 _35683_ (.A1(_11903_),
    .A2(_12927_),
    .ZN(_12928_));
 AOI21_X1 _35684_ (.A(_12928_),
    .B1(_12306_),
    .B2(_11828_),
    .ZN(_12929_));
 XNOR2_X2 _35685_ (.A(\core.keymem.prev_key1_reg[125] ),
    .B(_12293_),
    .ZN(_12930_));
 AOI221_X2 _35686_ (.A(_12929_),
    .B1(_12930_),
    .B2(_12027_),
    .C1(_12189_),
    .C2(_12680_),
    .ZN(_12931_));
 BUF_X2 _35687_ (.A(_12931_),
    .Z(_12932_));
 MUX2_X1 _35688_ (.A(\core.keymem.key_mem[10][125] ),
    .B(_12932_),
    .S(_12870_),
    .Z(_00993_));
 NAND2_X1 _35689_ (.A1(\core.keymem.key_mem[10][126] ),
    .A2(_12816_),
    .ZN(_12933_));
 OAI21_X1 _35690_ (.A(_12933_),
    .B1(_12905_),
    .B2(_12207_),
    .ZN(_00994_));
 NAND2_X1 _35691_ (.A1(_12208_),
    .A2(_11842_),
    .ZN(_12934_));
 NOR2_X1 _35692_ (.A1(_00172_),
    .A2(_11945_),
    .ZN(_12935_));
 BUF_X2 _35693_ (.A(\core.keymem.prev_key0_reg[127] ),
    .Z(_12936_));
 CLKBUF_X3 _35694_ (.A(\core.keymem.rcon_logic.tmp_rcon[0] ),
    .Z(_12937_));
 XNOR2_X1 _35695_ (.A(_12937_),
    .B(_09209_),
    .ZN(_12938_));
 MUX2_X1 _35696_ (.A(_10260_),
    .B(_12938_),
    .S(_11920_),
    .Z(_12939_));
 XNOR2_X2 _35697_ (.A(_12936_),
    .B(_12939_),
    .ZN(_12940_));
 AOI21_X2 _35698_ (.A(_12935_),
    .B1(_12940_),
    .B2(_12099_),
    .ZN(_12941_));
 XOR2_X2 _35699_ (.A(_12937_),
    .B(_09209_),
    .Z(_12942_));
 XNOR2_X2 _35700_ (.A(\core.keymem.prev_key1_reg[127] ),
    .B(_12942_),
    .ZN(_12943_));
 OAI221_X2 _35701_ (.A(_12934_),
    .B1(_12941_),
    .B2(_11904_),
    .C1(_12943_),
    .C2(_12705_),
    .ZN(_12944_));
 BUF_X2 _35702_ (.A(_12944_),
    .Z(_12945_));
 MUX2_X1 _35703_ (.A(\core.keymem.key_mem[10][127] ),
    .B(_12945_),
    .S(_12870_),
    .Z(_00995_));
 NOR2_X4 _35704_ (.A1(_11840_),
    .A2(_11848_),
    .ZN(_12946_));
 AND3_X1 _35705_ (.A1(_12148_),
    .A2(\core.key[12] ),
    .A3(_12946_),
    .ZN(_12947_));
 NOR2_X1 _35706_ (.A1(_00407_),
    .A2(_11917_),
    .ZN(_12948_));
 AOI21_X2 _35707_ (.A(_12947_),
    .B1(_12948_),
    .B2(_12808_),
    .ZN(_12949_));
 XNOR2_X1 _35708_ (.A(_07313_),
    .B(_12503_),
    .ZN(_12950_));
 BUF_X4 _35709_ (.A(_12349_),
    .Z(_12951_));
 OAI21_X2 _35710_ (.A(_12002_),
    .B1(_12950_),
    .B2(_12951_),
    .ZN(_12952_));
 XNOR2_X1 _35711_ (.A(_12481_),
    .B(_12482_),
    .ZN(_12953_));
 XNOR2_X2 _35712_ (.A(\core.keymem.prev_key0_reg[12] ),
    .B(_12953_),
    .ZN(_12954_));
 XNOR2_X2 _35713_ (.A(_11974_),
    .B(_12954_),
    .ZN(_12955_));
 AOI21_X2 _35714_ (.A(_11847_),
    .B1(_12844_),
    .B2(_12955_),
    .ZN(_12956_));
 OAI21_X4 _35715_ (.A(_12949_),
    .B1(_12952_),
    .B2(_12956_),
    .ZN(_12957_));
 CLKBUF_X2 _35716_ (.A(_12957_),
    .Z(_12958_));
 MUX2_X1 _35717_ (.A(\core.keymem.key_mem[10][12] ),
    .B(_12958_),
    .S(_12870_),
    .Z(_00996_));
 NAND2_X4 _35718_ (.A1(_16219_),
    .A2(_11826_),
    .ZN(_12959_));
 BUF_X1 _35719_ (.A(\core.keymem.prev_key0_reg[77] ),
    .Z(_12960_));
 XNOR2_X1 _35720_ (.A(_12960_),
    .B(_12835_),
    .ZN(_12961_));
 CLKBUF_X2 _35721_ (.A(\core.keymem.prev_key0_reg[45] ),
    .Z(_12962_));
 XOR2_X1 _35722_ (.A(\core.keymem.prev_key0_reg[13] ),
    .B(_12962_),
    .Z(_12963_));
 XNOR2_X1 _35723_ (.A(_12961_),
    .B(_12963_),
    .ZN(_12964_));
 XNOR2_X2 _35724_ (.A(_12836_),
    .B(_12964_),
    .ZN(_12965_));
 NAND2_X4 _35725_ (.A1(_16219_),
    .A2(_11820_),
    .ZN(_12966_));
 OAI22_X4 _35726_ (.A1(_12959_),
    .A2(_12965_),
    .B1(_12966_),
    .B2(\core.key[13] ),
    .ZN(_12967_));
 XNOR2_X2 _35727_ (.A(\core.keymem.prev_key1_reg[77] ),
    .B(_12840_),
    .ZN(_12968_));
 XOR2_X2 _35728_ (.A(\core.keymem.prev_key1_reg[45] ),
    .B(_12968_),
    .Z(_12969_));
 XNOR2_X1 _35729_ (.A(\core.keymem.prev_key1_reg[13] ),
    .B(_12969_),
    .ZN(_12970_));
 BUF_X4 _35730_ (.A(_11846_),
    .Z(_12971_));
 BUF_X4 _35731_ (.A(_12971_),
    .Z(_12972_));
 AOI21_X2 _35732_ (.A(_12967_),
    .B1(_12970_),
    .B2(_12972_),
    .ZN(_12973_));
 CLKBUF_X2 _35733_ (.A(_12973_),
    .Z(_12974_));
 BUF_X4 _35734_ (.A(_12805_),
    .Z(_12975_));
 MUX2_X1 _35735_ (.A(\core.keymem.key_mem[10][13] ),
    .B(_12974_),
    .S(_12975_),
    .Z(_00997_));
 NOR2_X1 _35736_ (.A1(\core.keymem.key_mem[10][14] ),
    .A2(_12807_),
    .ZN(_12976_));
 AND2_X1 _35737_ (.A1(\core.key[14] ),
    .A2(_11891_),
    .ZN(_12977_));
 BUF_X1 _35738_ (.A(\core.keymem.prev_key0_reg[14] ),
    .Z(_12978_));
 BUF_X1 _35739_ (.A(\core.keymem.prev_key0_reg[46] ),
    .Z(_12979_));
 XOR2_X2 _35740_ (.A(_12979_),
    .B(_12698_),
    .Z(_12980_));
 XNOR2_X1 _35741_ (.A(_12978_),
    .B(_12980_),
    .ZN(_12981_));
 XNOR2_X1 _35742_ (.A(_11996_),
    .B(_12981_),
    .ZN(_12982_));
 AOI21_X2 _35743_ (.A(_12977_),
    .B1(_12982_),
    .B2(_12365_),
    .ZN(_12983_));
 NOR2_X2 _35744_ (.A1(_12786_),
    .A2(_12983_),
    .ZN(_12984_));
 NOR3_X1 _35745_ (.A1(_12349_),
    .A2(_07466_),
    .A3(_11841_),
    .ZN(_12985_));
 NOR3_X1 _35746_ (.A1(_12349_),
    .A2(_07349_),
    .A3(_11841_),
    .ZN(_12986_));
 CLKBUF_X3 _35747_ (.A(\core.keymem.prev_key1_reg[46] ),
    .Z(_12987_));
 INV_X2 _35748_ (.A(_12987_),
    .ZN(_12988_));
 XNOR2_X2 _35749_ (.A(_12988_),
    .B(_12704_),
    .ZN(_12989_));
 MUX2_X1 _35750_ (.A(_12985_),
    .B(_12986_),
    .S(_12989_),
    .Z(_12990_));
 NOR4_X1 _35751_ (.A1(_07349_),
    .A2(_12987_),
    .A3(_12701_),
    .A4(_11840_),
    .ZN(_12991_));
 NAND2_X1 _35752_ (.A1(_07349_),
    .A2(_12987_),
    .ZN(_12992_));
 NOR3_X1 _35753_ (.A1(_12701_),
    .A2(_11840_),
    .A3(_12992_),
    .ZN(_12993_));
 OAI21_X1 _35754_ (.A(_12000_),
    .B1(_12991_),
    .B2(_12993_),
    .ZN(_12994_));
 NOR4_X1 _35755_ (.A1(_07466_),
    .A2(_12987_),
    .A3(_12702_),
    .A4(_11840_),
    .ZN(_12995_));
 NOR4_X1 _35756_ (.A1(_07349_),
    .A2(_12988_),
    .A3(_12702_),
    .A4(_11797_),
    .ZN(_12996_));
 OAI21_X1 _35757_ (.A(_12000_),
    .B1(_12995_),
    .B2(_12996_),
    .ZN(_12997_));
 NOR4_X1 _35758_ (.A1(_07466_),
    .A2(_12987_),
    .A3(_12701_),
    .A4(_11840_),
    .ZN(_12998_));
 NOR4_X2 _35759_ (.A1(_07349_),
    .A2(_12988_),
    .A3(_12701_),
    .A4(_11797_),
    .ZN(_12999_));
 OAI21_X2 _35760_ (.A(_12703_),
    .B1(_12998_),
    .B2(_12999_),
    .ZN(_13000_));
 NOR4_X1 _35761_ (.A1(_07349_),
    .A2(_12987_),
    .A3(_12702_),
    .A4(_11840_),
    .ZN(_13001_));
 NOR3_X1 _35762_ (.A1(_12702_),
    .A2(_11840_),
    .A3(_12992_),
    .ZN(_13002_));
 OAI21_X2 _35763_ (.A(_12703_),
    .B1(_13001_),
    .B2(_13002_),
    .ZN(_13003_));
 NAND4_X4 _35764_ (.A1(_12994_),
    .A2(_12997_),
    .A3(_13000_),
    .A4(_13003_),
    .ZN(_13004_));
 NOR3_X2 _35765_ (.A1(_12301_),
    .A2(_00409_),
    .A3(_13004_),
    .ZN(_13005_));
 NOR3_X4 _35766_ (.A1(_12984_),
    .A2(_12990_),
    .A3(_13005_),
    .ZN(_13006_));
 CLKBUF_X3 _35767_ (.A(_13006_),
    .Z(_13007_));
 AOI21_X1 _35768_ (.A(_12976_),
    .B1(_13007_),
    .B2(_12807_),
    .ZN(_00998_));
 XOR2_X1 _35769_ (.A(\core.keymem.prev_key0_reg[47] ),
    .B(\core.keymem.prev_key0_reg[79] ),
    .Z(_13008_));
 XNOR2_X1 _35770_ (.A(\core.keymem.prev_key0_reg[15] ),
    .B(_13008_),
    .ZN(_13009_));
 XNOR2_X2 _35771_ (.A(_12013_),
    .B(_13009_),
    .ZN(_13010_));
 NOR2_X4 _35772_ (.A1(_11797_),
    .A2(_11818_),
    .ZN(_13011_));
 AOI221_X2 _35773_ (.A(_11846_),
    .B1(\core.key[15] ),
    .B2(_12946_),
    .C1(_13010_),
    .C2(_13011_),
    .ZN(_13012_));
 NAND2_X1 _35774_ (.A1(_00410_),
    .A2(_11799_),
    .ZN(_13013_));
 XNOR2_X1 _35775_ (.A(_07357_),
    .B(_12517_),
    .ZN(_13014_));
 OAI221_X2 _35776_ (.A(_16228_),
    .B1(_11909_),
    .B2(_13013_),
    .C1(_13014_),
    .C2(_12705_),
    .ZN(_13015_));
 NOR2_X2 _35777_ (.A1(_13012_),
    .A2(_13015_),
    .ZN(_13016_));
 CLKBUF_X2 _35778_ (.A(_13016_),
    .Z(_13017_));
 MUX2_X1 _35779_ (.A(\core.keymem.key_mem[10][15] ),
    .B(_13017_),
    .S(_12975_),
    .Z(_00999_));
 XOR2_X1 _35780_ (.A(\core.keymem.prev_key0_reg[80] ),
    .B(\core.keymem.prev_key0_reg[112] ),
    .Z(_13018_));
 XNOR2_X1 _35781_ (.A(\core.keymem.prev_key0_reg[16] ),
    .B(\core.keymem.prev_key0_reg[48] ),
    .ZN(_13019_));
 XNOR2_X1 _35782_ (.A(_13018_),
    .B(_13019_),
    .ZN(_13020_));
 XNOR2_X1 _35783_ (.A(net13),
    .B(_13020_),
    .ZN(_13021_));
 NOR2_X1 _35784_ (.A1(_12241_),
    .A2(_13021_),
    .ZN(_13022_));
 INV_X1 _35785_ (.A(_12526_),
    .ZN(_13023_));
 XNOR2_X2 _35786_ (.A(_08195_),
    .B(_12527_),
    .ZN(_13024_));
 XNOR2_X2 _35787_ (.A(_13023_),
    .B(_13024_),
    .ZN(_13025_));
 XOR2_X2 _35788_ (.A(_12026_),
    .B(_13025_),
    .Z(_13026_));
 INV_X1 _35789_ (.A(\core.key[16] ),
    .ZN(_13027_));
 AOI221_X2 _35790_ (.A(_13022_),
    .B1(_13026_),
    .B2(_12027_),
    .C1(_13027_),
    .C2(_12269_),
    .ZN(_13028_));
 BUF_X2 _35791_ (.A(_13028_),
    .Z(_13029_));
 MUX2_X1 _35792_ (.A(\core.keymem.key_mem[10][16] ),
    .B(_13029_),
    .S(_12975_),
    .Z(_01000_));
 NAND2_X1 _35793_ (.A1(\core.keymem.key_mem[10][17] ),
    .A2(_12816_),
    .ZN(_13030_));
 XNOR2_X2 _35794_ (.A(\core.keymem.prev_key0_reg[81] ),
    .B(\core.keymem.prev_key0_reg[113] ),
    .ZN(_13031_));
 XOR2_X1 _35795_ (.A(\core.keymem.prev_key0_reg[17] ),
    .B(\core.keymem.prev_key0_reg[49] ),
    .Z(_13032_));
 XNOR2_X1 _35796_ (.A(_13031_),
    .B(_13032_),
    .ZN(_13033_));
 XNOR2_X2 _35797_ (.A(_12862_),
    .B(_13033_),
    .ZN(_13034_));
 AND2_X1 _35798_ (.A1(_12365_),
    .A2(_13034_),
    .ZN(_13035_));
 NAND2_X1 _35799_ (.A1(\core.key[17] ),
    .A2(_12345_),
    .ZN(_13036_));
 NAND2_X1 _35800_ (.A1(_12335_),
    .A2(_13036_),
    .ZN(_13037_));
 XNOR2_X2 _35801_ (.A(\core.keymem.prev_key1_reg[81] ),
    .B(_12865_),
    .ZN(_13038_));
 XOR2_X2 _35802_ (.A(\core.keymem.prev_key1_reg[49] ),
    .B(\core.keymem.prev_key1_reg[17] ),
    .Z(_13039_));
 XNOR2_X2 _35803_ (.A(_13038_),
    .B(_13039_),
    .ZN(_13040_));
 OAI22_X4 _35804_ (.A1(_13035_),
    .A2(_13037_),
    .B1(_13040_),
    .B2(_12263_),
    .ZN(_13041_));
 CLKBUF_X3 _35805_ (.A(_13041_),
    .Z(_13042_));
 OAI21_X1 _35806_ (.A(_13030_),
    .B1(_13042_),
    .B2(_12896_),
    .ZN(_01001_));
 BUF_X4 _35807_ (.A(_12039_),
    .Z(_13043_));
 BUF_X2 _35808_ (.A(\core.keymem.prev_key0_reg[18] ),
    .Z(_13044_));
 INV_X1 _35809_ (.A(_13044_),
    .ZN(_13045_));
 BUF_X2 _35810_ (.A(\core.keymem.prev_key0_reg[50] ),
    .Z(_13046_));
 NOR2_X1 _35811_ (.A1(_13045_),
    .A2(_13046_),
    .ZN(_13047_));
 CLKBUF_X3 _35812_ (.A(\core.keymem.prev_key0_reg[82] ),
    .Z(_13048_));
 NOR2_X1 _35813_ (.A1(_13048_),
    .A2(_12037_),
    .ZN(_13049_));
 AND2_X1 _35814_ (.A1(_13047_),
    .A2(_13049_),
    .ZN(_13050_));
 INV_X1 _35815_ (.A(\core.keymem.prev_key0_reg[50] ),
    .ZN(_13051_));
 NOR2_X1 _35816_ (.A1(_13044_),
    .A2(_13051_),
    .ZN(_13052_));
 AND2_X1 _35817_ (.A1(_13052_),
    .A2(_13049_),
    .ZN(_13053_));
 OAI221_X2 _35818_ (.A(_12044_),
    .B1(_13043_),
    .B2(_12041_),
    .C1(_13050_),
    .C2(_13053_),
    .ZN(_13054_));
 NOR2_X1 _35819_ (.A1(_13044_),
    .A2(_13046_),
    .ZN(_13055_));
 INV_X2 _35820_ (.A(\core.keymem.prev_key0_reg[82] ),
    .ZN(_13056_));
 NOR2_X1 _35821_ (.A1(_13056_),
    .A2(_12037_),
    .ZN(_13057_));
 AND2_X1 _35822_ (.A1(_13055_),
    .A2(_13057_),
    .ZN(_13058_));
 NAND2_X1 _35823_ (.A1(_13044_),
    .A2(_13046_),
    .ZN(_13059_));
 NOR3_X1 _35824_ (.A1(_13056_),
    .A2(_12037_),
    .A3(_13059_),
    .ZN(_13060_));
 OAI221_X2 _35825_ (.A(_11925_),
    .B1(_13043_),
    .B2(_12041_),
    .C1(_13058_),
    .C2(_13060_),
    .ZN(_13061_));
 NOR2_X1 _35826_ (.A1(_13048_),
    .A2(_12038_),
    .ZN(_13062_));
 AND2_X1 _35827_ (.A1(_13055_),
    .A2(_13062_),
    .ZN(_13063_));
 NOR3_X1 _35828_ (.A1(_13048_),
    .A2(_12038_),
    .A3(_13059_),
    .ZN(_13064_));
 OAI221_X2 _35829_ (.A(_11925_),
    .B1(_13043_),
    .B2(_12041_),
    .C1(_13063_),
    .C2(_13064_),
    .ZN(_13065_));
 NAND2_X1 _35830_ (.A1(_13048_),
    .A2(_12037_),
    .ZN(_13066_));
 NOR3_X1 _35831_ (.A1(_13045_),
    .A2(_13046_),
    .A3(_13066_),
    .ZN(_13067_));
 NOR3_X1 _35832_ (.A1(_13044_),
    .A2(_13051_),
    .A3(_13066_),
    .ZN(_13068_));
 OAI221_X2 _35833_ (.A(_11925_),
    .B1(_13043_),
    .B2(_12041_),
    .C1(_13067_),
    .C2(_13068_),
    .ZN(_13069_));
 NAND4_X2 _35834_ (.A1(_13054_),
    .A2(_13061_),
    .A3(_13065_),
    .A4(_13069_),
    .ZN(_13070_));
 NAND3_X1 _35835_ (.A1(_11825_),
    .A2(_13049_),
    .A3(_13055_),
    .ZN(_13071_));
 NAND4_X1 _35836_ (.A1(_13044_),
    .A2(_13046_),
    .A3(_11825_),
    .A4(_13049_),
    .ZN(_13072_));
 AOI221_X1 _35837_ (.A(_13043_),
    .B1(_13071_),
    .B2(_13072_),
    .C1(_12046_),
    .C2(_12175_),
    .ZN(_13073_));
 NAND3_X1 _35838_ (.A1(_11825_),
    .A2(_13047_),
    .A3(_13057_),
    .ZN(_13074_));
 NAND3_X1 _35839_ (.A1(_11825_),
    .A2(_13052_),
    .A3(_13057_),
    .ZN(_13075_));
 AOI221_X1 _35840_ (.A(_13043_),
    .B1(_13074_),
    .B2(_13075_),
    .C1(_12046_),
    .C2(_12175_),
    .ZN(_13076_));
 OR2_X1 _35841_ (.A1(_13073_),
    .A2(_13076_),
    .ZN(_13077_));
 NAND3_X1 _35842_ (.A1(_11925_),
    .A2(_13047_),
    .A3(_13062_),
    .ZN(_13078_));
 NAND3_X1 _35843_ (.A1(_11827_),
    .A2(_13052_),
    .A3(_13062_),
    .ZN(_13079_));
 AOI21_X2 _35844_ (.A(_12042_),
    .B1(_13078_),
    .B2(_13079_),
    .ZN(_13080_));
 NAND4_X1 _35845_ (.A1(_13048_),
    .A2(_12037_),
    .A3(_11860_),
    .A4(_13055_),
    .ZN(_13081_));
 OR3_X1 _35846_ (.A1(_11819_),
    .A2(_13059_),
    .A3(_13066_),
    .ZN(_13082_));
 AOI21_X2 _35847_ (.A(_12042_),
    .B1(_13081_),
    .B2(_13082_),
    .ZN(_13083_));
 NOR4_X4 _35848_ (.A1(_13070_),
    .A2(_13077_),
    .A3(_13080_),
    .A4(_13083_),
    .ZN(_13084_));
 NAND2_X1 _35849_ (.A1(\core.key[18] ),
    .A2(_12101_),
    .ZN(_13085_));
 AND2_X1 _35850_ (.A1(_12098_),
    .A2(_13085_),
    .ZN(_13086_));
 INV_X1 _35851_ (.A(\core.keymem.prev_key1_reg[18] ),
    .ZN(_13087_));
 INV_X1 _35852_ (.A(\core.keymem.prev_key1_reg[50] ),
    .ZN(_13088_));
 XNOR2_X1 _35853_ (.A(\core.keymem.prev_key1_reg[82] ),
    .B(\core.keymem.prev_key1_reg[114] ),
    .ZN(_13089_));
 XNOR2_X2 _35854_ (.A(_12046_),
    .B(_13089_),
    .ZN(_13090_));
 XNOR2_X2 _35855_ (.A(_13088_),
    .B(_13090_),
    .ZN(_13091_));
 XNOR2_X2 _35856_ (.A(_13087_),
    .B(_13091_),
    .ZN(_13092_));
 AOI22_X4 _35857_ (.A1(_13084_),
    .A2(_13086_),
    .B1(_13092_),
    .B2(_12028_),
    .ZN(_13093_));
 BUF_X2 _35858_ (.A(_13093_),
    .Z(_13094_));
 MUX2_X1 _35859_ (.A(\core.keymem.key_mem[10][18] ),
    .B(_13094_),
    .S(_12975_),
    .Z(_01002_));
 BUF_X4 _35860_ (.A(_12815_),
    .Z(_13095_));
 NAND2_X1 _35861_ (.A1(\core.keymem.key_mem[10][19] ),
    .A2(_13095_),
    .ZN(_13096_));
 NOR3_X1 _35862_ (.A1(_06677_),
    .A2(_00436_),
    .A3(_11875_),
    .ZN(_13097_));
 AND2_X1 _35863_ (.A1(_12148_),
    .A2(\core.key[19] ),
    .ZN(_13098_));
 XNOR2_X1 _35864_ (.A(\core.keymem.prev_key1_reg[83] ),
    .B(\core.keymem.prev_key1_reg[115] ),
    .ZN(_13099_));
 XNOR2_X2 _35865_ (.A(_11961_),
    .B(_13099_),
    .ZN(_13100_));
 XNOR2_X2 _35866_ (.A(\core.keymem.prev_key1_reg[51] ),
    .B(_13100_),
    .ZN(_13101_));
 XNOR2_X2 _35867_ (.A(\core.keymem.prev_key1_reg[19] ),
    .B(_13101_),
    .ZN(_13102_));
 AOI21_X4 _35868_ (.A(_12680_),
    .B1(_13102_),
    .B2(_11866_),
    .ZN(_13103_));
 XNOR2_X2 _35869_ (.A(\core.keymem.prev_key0_reg[51] ),
    .B(\core.keymem.prev_key0_reg[83] ),
    .ZN(_13104_));
 XOR2_X2 _35870_ (.A(\core.keymem.prev_key0_reg[19] ),
    .B(_13104_),
    .Z(_13105_));
 XNOR2_X2 _35871_ (.A(_12052_),
    .B(_13105_),
    .ZN(_13106_));
 OAI21_X1 _35872_ (.A(_12156_),
    .B1(_12345_),
    .B2(_13106_),
    .ZN(_13107_));
 AOI221_X2 _35873_ (.A(_13097_),
    .B1(_13098_),
    .B2(_12946_),
    .C1(_13103_),
    .C2(_13107_),
    .ZN(_13108_));
 CLKBUF_X3 _35874_ (.A(_13108_),
    .Z(_13109_));
 OAI21_X1 _35875_ (.A(_13096_),
    .B1(_13109_),
    .B2(_12896_),
    .ZN(_01003_));
 AOI21_X1 _35876_ (.A(_06676_),
    .B1(_12227_),
    .B2(_11798_),
    .ZN(_13110_));
 XOR2_X1 _35877_ (.A(\core.keymem.prev_key1_reg[1] ),
    .B(_00372_),
    .Z(_13111_));
 XNOR2_X1 _35878_ (.A(_12359_),
    .B(_13111_),
    .ZN(_13112_));
 XOR2_X1 _35879_ (.A(_09777_),
    .B(_13112_),
    .Z(_13113_));
 OAI21_X1 _35880_ (.A(_13110_),
    .B1(_13113_),
    .B2(_11799_),
    .ZN(_13114_));
 NAND2_X2 _35881_ (.A1(_16228_),
    .A2(_13114_),
    .ZN(_13115_));
 INV_X1 _35882_ (.A(\core.keymem.prev_key0_reg[1] ),
    .ZN(_13116_));
 CLKBUF_X2 _35883_ (.A(\core.keymem.prev_key0_reg[33] ),
    .Z(_13117_));
 BUF_X2 _35884_ (.A(\core.keymem.prev_key0_reg[65] ),
    .Z(_13118_));
 XNOR2_X1 _35885_ (.A(_13117_),
    .B(_13118_),
    .ZN(_13119_));
 XNOR2_X1 _35886_ (.A(_13116_),
    .B(_13119_),
    .ZN(_13120_));
 XNOR2_X2 _35887_ (.A(_12772_),
    .B(_13120_),
    .ZN(_13121_));
 NOR2_X1 _35888_ (.A1(_11997_),
    .A2(_13121_),
    .ZN(_13122_));
 INV_X1 _35889_ (.A(\core.key[1] ),
    .ZN(_13123_));
 NOR2_X1 _35890_ (.A1(\core.keymem.prev_key0_reg[1] ),
    .A2(_13117_),
    .ZN(_13124_));
 AND4_X1 _35891_ (.A1(_13118_),
    .A2(\core.keymem.prev_key0_reg[97] ),
    .A3(_12771_),
    .A4(_13124_),
    .ZN(_13125_));
 NOR3_X1 _35892_ (.A1(_13116_),
    .A2(_13117_),
    .A3(_13118_),
    .ZN(_13126_));
 INV_X1 _35893_ (.A(_13118_),
    .ZN(_13127_));
 AND4_X1 _35894_ (.A1(_13116_),
    .A2(_13117_),
    .A3(_13127_),
    .A4(\core.keymem.prev_key0_reg[97] ),
    .ZN(_13128_));
 AOI221_X1 _35895_ (.A(_13125_),
    .B1(_13126_),
    .B2(_12772_),
    .C1(_12771_),
    .C2(_13128_),
    .ZN(_13129_));
 AOI21_X1 _35896_ (.A(_13123_),
    .B1(_12333_),
    .B2(_13129_),
    .ZN(_13130_));
 OAI21_X2 _35897_ (.A(_12002_),
    .B1(_13122_),
    .B2(_13130_),
    .ZN(_13131_));
 BUF_X4 _35898_ (.A(_11909_),
    .Z(_13132_));
 AOI21_X4 _35899_ (.A(_13115_),
    .B1(_13131_),
    .B2(_13132_),
    .ZN(_13133_));
 BUF_X2 _35900_ (.A(_13133_),
    .Z(_13134_));
 MUX2_X1 _35901_ (.A(\core.keymem.key_mem[10][1] ),
    .B(_13134_),
    .S(_12975_),
    .Z(_01004_));
 AND2_X1 _35902_ (.A1(\core.keymem.prev_key0_reg[20] ),
    .A2(_13011_),
    .ZN(_13135_));
 NAND2_X4 _35903_ (.A1(_11813_),
    .A2(_11848_),
    .ZN(_13136_));
 NOR2_X1 _35904_ (.A1(\core.keymem.prev_key0_reg[20] ),
    .A2(_13136_),
    .ZN(_13137_));
 MUX2_X2 _35905_ (.A(_13135_),
    .B(_13137_),
    .S(_12566_),
    .Z(_13138_));
 NAND2_X1 _35906_ (.A1(\core.key[20] ),
    .A2(_12946_),
    .ZN(_13139_));
 NAND2_X1 _35907_ (.A1(_12156_),
    .A2(_13139_),
    .ZN(_13140_));
 NOR2_X4 _35908_ (.A1(_13138_),
    .A2(_13140_),
    .ZN(_13141_));
 NAND2_X1 _35909_ (.A1(_00437_),
    .A2(_11799_),
    .ZN(_13142_));
 XNOR2_X1 _35910_ (.A(_08233_),
    .B(_12546_),
    .ZN(_13143_));
 OAI221_X2 _35911_ (.A(_16228_),
    .B1(_11909_),
    .B2(_13142_),
    .C1(_13143_),
    .C2(_12001_),
    .ZN(_13144_));
 NOR2_X2 _35912_ (.A1(_13141_),
    .A2(_13144_),
    .ZN(_13145_));
 BUF_X2 _35913_ (.A(_13145_),
    .Z(_13146_));
 MUX2_X1 _35914_ (.A(\core.keymem.key_mem[10][20] ),
    .B(_13146_),
    .S(_12975_),
    .Z(_01005_));
 XNOR2_X1 _35915_ (.A(\core.keymem.prev_key0_reg[21] ),
    .B(\core.keymem.prev_key0_reg[53] ),
    .ZN(_13147_));
 XNOR2_X1 _35916_ (.A(_12572_),
    .B(_13147_),
    .ZN(_13148_));
 XNOR2_X1 _35917_ (.A(_12571_),
    .B(_13148_),
    .ZN(_13149_));
 NAND2_X1 _35918_ (.A1(_12149_),
    .A2(_13149_),
    .ZN(_13150_));
 NAND2_X1 _35919_ (.A1(\core.key[21] ),
    .A2(_11989_),
    .ZN(_13151_));
 AND2_X1 _35920_ (.A1(_13150_),
    .A2(_13151_),
    .ZN(_13152_));
 XNOR2_X2 _35921_ (.A(\core.keymem.prev_key1_reg[21] ),
    .B(_12581_),
    .ZN(_13153_));
 AOI22_X4 _35922_ (.A1(_12335_),
    .A2(_13152_),
    .B1(_13153_),
    .B2(_12028_),
    .ZN(_13154_));
 CLKBUF_X2 _35923_ (.A(_13154_),
    .Z(_13155_));
 MUX2_X1 _35924_ (.A(\core.keymem.key_mem[10][21] ),
    .B(_13155_),
    .S(_12975_),
    .Z(_01006_));
 NOR2_X1 _35925_ (.A1(\core.keymem.key_mem[10][22] ),
    .A2(_12807_),
    .ZN(_13156_));
 OAI21_X1 _35926_ (.A(_11874_),
    .B1(_12966_),
    .B2(\core.key[22] ),
    .ZN(_13157_));
 BUF_X2 _35927_ (.A(\core.keymem.prev_key1_reg[54] ),
    .Z(_13158_));
 XOR2_X2 _35928_ (.A(_08298_),
    .B(_13158_),
    .Z(_13159_));
 NOR3_X1 _35929_ (.A1(_16219_),
    .A2(_12727_),
    .A3(_13159_),
    .ZN(_13160_));
 OR4_X1 _35930_ (.A1(_16219_),
    .A2(_08299_),
    .A3(_13158_),
    .A4(_12727_),
    .ZN(_13161_));
 NAND2_X1 _35931_ (.A1(_11811_),
    .A2(_12727_),
    .ZN(_13162_));
 OAI21_X1 _35932_ (.A(_13161_),
    .B1(_13162_),
    .B2(_13159_),
    .ZN(_13163_));
 MUX2_X1 _35933_ (.A(_13160_),
    .B(_13163_),
    .S(_12728_),
    .Z(_13164_));
 AND2_X1 _35934_ (.A1(_12727_),
    .A2(_13159_),
    .ZN(_13165_));
 INV_X1 _35935_ (.A(_13158_),
    .ZN(_13166_));
 NOR3_X1 _35936_ (.A1(_08298_),
    .A2(_13166_),
    .A3(_12727_),
    .ZN(_13167_));
 MUX2_X1 _35937_ (.A(_13165_),
    .B(_13167_),
    .S(_12728_),
    .Z(_13168_));
 AOI211_X2 _35938_ (.A(_13157_),
    .B(_13164_),
    .C1(_11866_),
    .C2(_13168_),
    .ZN(_13169_));
 OR2_X2 _35939_ (.A1(_08483_),
    .A2(_09170_),
    .ZN(_13170_));
 MUX2_X2 _35940_ (.A(_08101_),
    .B(_13170_),
    .S(_12917_),
    .Z(_13171_));
 CLKBUF_X2 _35941_ (.A(\core.keymem.prev_key0_reg[54] ),
    .Z(_13172_));
 XOR2_X2 _35942_ (.A(\core.keymem.prev_key0_reg[22] ),
    .B(_13172_),
    .Z(_13173_));
 NOR3_X1 _35943_ (.A1(_12732_),
    .A2(_12959_),
    .A3(_13173_),
    .ZN(_13174_));
 INV_X1 _35944_ (.A(_13172_),
    .ZN(_13175_));
 NOR2_X4 _35945_ (.A1(_11811_),
    .A2(_11818_),
    .ZN(_13176_));
 AND4_X1 _35946_ (.A1(\core.keymem.prev_key0_reg[22] ),
    .A2(_13175_),
    .A3(_12732_),
    .A4(_13176_),
    .ZN(_13177_));
 NOR2_X1 _35947_ (.A1(_13174_),
    .A2(_13177_),
    .ZN(_13178_));
 NOR3_X1 _35948_ (.A1(\core.keymem.prev_key0_reg[118] ),
    .A2(_13171_),
    .A3(_13178_),
    .ZN(_13179_));
 AND4_X1 _35949_ (.A1(_12732_),
    .A2(\core.keymem.prev_key0_reg[118] ),
    .A3(_13176_),
    .A4(_13173_),
    .ZN(_13180_));
 AOI21_X2 _35950_ (.A(_13179_),
    .B1(_13180_),
    .B2(_13171_),
    .ZN(_13181_));
 XNOR2_X1 _35951_ (.A(_12732_),
    .B(_13173_),
    .ZN(_13182_));
 NOR2_X1 _35952_ (.A1(_12737_),
    .A2(_13182_),
    .ZN(_13183_));
 INV_X1 _35953_ (.A(\core.keymem.prev_key0_reg[22] ),
    .ZN(_13184_));
 NOR4_X2 _35954_ (.A1(_13184_),
    .A2(_13175_),
    .A3(_12732_),
    .A4(_12733_),
    .ZN(_13185_));
 NOR3_X1 _35955_ (.A1(_13172_),
    .A2(_12732_),
    .A3(_12733_),
    .ZN(_13186_));
 AND3_X1 _35956_ (.A1(_13172_),
    .A2(_12732_),
    .A3(_12733_),
    .ZN(_13187_));
 MUX2_X1 _35957_ (.A(_13186_),
    .B(_13187_),
    .S(_12736_),
    .Z(_13188_));
 AOI221_X2 _35958_ (.A(_13183_),
    .B1(_13185_),
    .B2(_13171_),
    .C1(_13184_),
    .C2(_13188_),
    .ZN(_13189_));
 OAI211_X4 _35959_ (.A(_13169_),
    .B(_13181_),
    .C1(_12959_),
    .C2(_13189_),
    .ZN(_13190_));
 CLKBUF_X3 _35960_ (.A(_13190_),
    .Z(_13191_));
 AOI21_X1 _35961_ (.A(_13156_),
    .B1(_13191_),
    .B2(_12807_),
    .ZN(_01007_));
 AOI21_X1 _35962_ (.A(_06676_),
    .B1(_00016_),
    .B2(_11798_),
    .ZN(_13192_));
 INV_X1 _35963_ (.A(_13192_),
    .ZN(_13193_));
 AOI21_X1 _35964_ (.A(_13193_),
    .B1(_12267_),
    .B2(_11875_),
    .ZN(_13194_));
 OR3_X2 _35965_ (.A1(_12261_),
    .A2(_12271_),
    .A3(_13194_),
    .ZN(_13195_));
 BUF_X2 _35966_ (.A(_13195_),
    .Z(_13196_));
 MUX2_X1 _35967_ (.A(\core.keymem.key_mem[10][23] ),
    .B(_13196_),
    .S(_12975_),
    .Z(_01008_));
 NAND2_X1 _35968_ (.A1(\core.keymem.key_mem[10][24] ),
    .A2(_13095_),
    .ZN(_13197_));
 AOI21_X1 _35969_ (.A(_11903_),
    .B1(_11892_),
    .B2(_00019_),
    .ZN(_13198_));
 INV_X1 _35970_ (.A(_13198_),
    .ZN(_13199_));
 XOR2_X2 _35971_ (.A(\core.keymem.prev_key0_reg[24] ),
    .B(\core.keymem.prev_key0_reg[56] ),
    .Z(_13200_));
 XNOR2_X2 _35972_ (.A(\core.keymem.prev_key0_reg[88] ),
    .B(_12118_),
    .ZN(_13201_));
 XNOR2_X2 _35973_ (.A(_13200_),
    .B(_13201_),
    .ZN(_13202_));
 AOI21_X4 _35974_ (.A(_13199_),
    .B1(_13202_),
    .B2(_12365_),
    .ZN(_13203_));
 BUF_X2 _35975_ (.A(\core.keymem.prev_key1_reg[88] ),
    .Z(_13204_));
 XNOR2_X2 _35976_ (.A(\core.keymem.prev_key1_reg[56] ),
    .B(_13204_),
    .ZN(_13205_));
 XNOR2_X1 _35977_ (.A(_09318_),
    .B(_00018_),
    .ZN(_13206_));
 XNOR2_X1 _35978_ (.A(_13205_),
    .B(_13206_),
    .ZN(_13207_));
 XNOR2_X1 _35979_ (.A(_12121_),
    .B(_13207_),
    .ZN(_13208_));
 NOR2_X2 _35980_ (.A1(_12705_),
    .A2(_13208_),
    .ZN(_13209_));
 NOR2_X4 _35981_ (.A1(_00017_),
    .A2(_12347_),
    .ZN(_13210_));
 NOR3_X4 _35982_ (.A1(_13203_),
    .A2(_13209_),
    .A3(_13210_),
    .ZN(_13211_));
 CLKBUF_X3 _35983_ (.A(_13211_),
    .Z(_13212_));
 OAI21_X1 _35984_ (.A(_13197_),
    .B1(_13212_),
    .B2(_12896_),
    .ZN(_01009_));
 CLKBUF_X2 _35985_ (.A(\core.keymem.prev_key1_reg[89] ),
    .Z(_13213_));
 XNOR2_X2 _35986_ (.A(\core.keymem.prev_key1_reg[57] ),
    .B(_13213_),
    .ZN(_13214_));
 XOR2_X1 _35987_ (.A(\core.keymem.prev_key1_reg[25] ),
    .B(_00021_),
    .Z(_13215_));
 XNOR2_X1 _35988_ (.A(_13214_),
    .B(_13215_),
    .ZN(_13216_));
 XNOR2_X1 _35989_ (.A(_12154_),
    .B(_13216_),
    .ZN(_13217_));
 AOI21_X2 _35990_ (.A(_12779_),
    .B1(_13217_),
    .B2(_11847_),
    .ZN(_13218_));
 AND2_X1 _35991_ (.A1(_00022_),
    .A2(_11892_),
    .ZN(_13219_));
 OR2_X1 _35992_ (.A1(_11866_),
    .A2(_13219_),
    .ZN(_13220_));
 BUF_X1 _35993_ (.A(\core.keymem.prev_key0_reg[57] ),
    .Z(_13221_));
 XNOR2_X1 _35994_ (.A(\core.keymem.prev_key0_reg[25] ),
    .B(_13221_),
    .ZN(_13222_));
 CLKBUF_X2 _35995_ (.A(\core.keymem.prev_key0_reg[89] ),
    .Z(_13223_));
 XNOR2_X1 _35996_ (.A(_13223_),
    .B(_12126_),
    .ZN(_13224_));
 XNOR2_X1 _35997_ (.A(_13222_),
    .B(_13224_),
    .ZN(_13225_));
 INV_X1 _35998_ (.A(_13225_),
    .ZN(_13226_));
 NOR3_X2 _35999_ (.A1(_12917_),
    .A2(_12152_),
    .A3(_12153_),
    .ZN(_13227_));
 AOI21_X2 _36000_ (.A(_12176_),
    .B1(_09708_),
    .B2(_09776_),
    .ZN(_13228_));
 OAI21_X2 _36001_ (.A(_13226_),
    .B1(_13227_),
    .B2(_13228_),
    .ZN(_13229_));
 OR3_X2 _36002_ (.A1(_13228_),
    .A2(_13227_),
    .A3(_13226_),
    .ZN(_13230_));
 AOI21_X4 _36003_ (.A(_11997_),
    .B1(_13229_),
    .B2(_13230_),
    .ZN(_13231_));
 OAI21_X4 _36004_ (.A(_13218_),
    .B1(_13220_),
    .B2(_13231_),
    .ZN(_13232_));
 BUF_X2 _36005_ (.A(_13232_),
    .Z(_13233_));
 MUX2_X1 _36006_ (.A(\core.keymem.key_mem[10][25] ),
    .B(_13233_),
    .S(_12975_),
    .Z(_01010_));
 AOI21_X1 _36007_ (.A(_11987_),
    .B1(_12629_),
    .B2(_00025_),
    .ZN(_13234_));
 XNOR2_X2 _36008_ (.A(\core.keymem.prev_key0_reg[90] ),
    .B(\core.keymem.prev_key0_reg[122] ),
    .ZN(_13235_));
 XNOR2_X1 _36009_ (.A(\core.keymem.prev_key0_reg[26] ),
    .B(\core.keymem.prev_key0_reg[58] ),
    .ZN(_13236_));
 XNOR2_X1 _36010_ (.A(_13235_),
    .B(_13236_),
    .ZN(_13237_));
 XNOR2_X1 _36011_ (.A(_12898_),
    .B(_13237_),
    .ZN(_13238_));
 OAI21_X2 _36012_ (.A(_13234_),
    .B1(_13238_),
    .B2(_12172_),
    .ZN(_13239_));
 NAND2_X2 _36013_ (.A1(_12285_),
    .A2(_13239_),
    .ZN(_13240_));
 CLKBUF_X2 _36014_ (.A(_13240_),
    .Z(_13241_));
 MUX2_X1 _36015_ (.A(\core.keymem.key_mem[10][26] ),
    .B(_13241_),
    .S(_12975_),
    .Z(_01011_));
 CLKBUF_X2 _36016_ (.A(\core.keymem.prev_key0_reg[59] ),
    .Z(_13242_));
 INV_X1 _36017_ (.A(_13242_),
    .ZN(_13243_));
 BUF_X2 _36018_ (.A(\core.keymem.prev_key0_reg[91] ),
    .Z(_13244_));
 NAND3_X1 _36019_ (.A1(_11831_),
    .A2(_13244_),
    .A3(_12174_),
    .ZN(_13245_));
 INV_X1 _36020_ (.A(_13244_),
    .ZN(_13246_));
 NAND3_X1 _36021_ (.A1(_11831_),
    .A2(_13246_),
    .A3(_12173_),
    .ZN(_13247_));
 AOI22_X1 _36022_ (.A1(_12379_),
    .A2(_12380_),
    .B1(_13245_),
    .B2(_13247_),
    .ZN(_13248_));
 NAND3_X1 _36023_ (.A1(_11830_),
    .A2(_13246_),
    .A3(_12174_),
    .ZN(_13249_));
 NAND3_X1 _36024_ (.A1(_11830_),
    .A2(_13244_),
    .A3(_12173_),
    .ZN(_13250_));
 AOI211_X2 _36025_ (.A(_09934_),
    .B(_09948_),
    .C1(_13249_),
    .C2(_13250_),
    .ZN(_13251_));
 NAND4_X1 _36026_ (.A1(_11850_),
    .A2(_12166_),
    .A3(_13246_),
    .A4(_12174_),
    .ZN(_13252_));
 NOR2_X1 _36027_ (.A1(_11829_),
    .A2(_12166_),
    .ZN(_13253_));
 NAND3_X1 _36028_ (.A1(_13244_),
    .A2(_12174_),
    .A3(_13253_),
    .ZN(_13254_));
 AOI22_X1 _36029_ (.A1(_08827_),
    .A2(_08885_),
    .B1(_13252_),
    .B2(_13254_),
    .ZN(_13255_));
 NAND3_X1 _36030_ (.A1(_13246_),
    .A2(_12173_),
    .A3(_13253_),
    .ZN(_13256_));
 NAND4_X1 _36031_ (.A1(_11850_),
    .A2(_12166_),
    .A3(_13244_),
    .A4(_12173_),
    .ZN(_13257_));
 AOI22_X1 _36032_ (.A1(_08827_),
    .A2(_08885_),
    .B1(_13256_),
    .B2(_13257_),
    .ZN(_13258_));
 NOR4_X1 _36033_ (.A1(_13248_),
    .A2(_13251_),
    .A3(_13255_),
    .A4(_13258_),
    .ZN(_13259_));
 NOR4_X1 _36034_ (.A1(_12040_),
    .A2(_12166_),
    .A3(_13244_),
    .A4(_12173_),
    .ZN(_13260_));
 NAND2_X1 _36035_ (.A1(_11851_),
    .A2(_12166_),
    .ZN(_13261_));
 NOR3_X1 _36036_ (.A1(_13246_),
    .A2(_12173_),
    .A3(_13261_),
    .ZN(_13262_));
 OAI21_X1 _36037_ (.A(_08886_),
    .B1(_13260_),
    .B2(_13262_),
    .ZN(_13263_));
 NOR3_X1 _36038_ (.A1(_13244_),
    .A2(_12174_),
    .A3(_13261_),
    .ZN(_13264_));
 AND3_X1 _36039_ (.A1(_13244_),
    .A2(_12173_),
    .A3(_13253_),
    .ZN(_13265_));
 OAI21_X1 _36040_ (.A(_08886_),
    .B1(_13264_),
    .B2(_13265_),
    .ZN(_13266_));
 AND3_X2 _36041_ (.A1(_13259_),
    .A2(_13263_),
    .A3(_13266_),
    .ZN(_13267_));
 AND4_X1 _36042_ (.A1(\core.keymem.prev_key0_reg[27] ),
    .A2(_13243_),
    .A3(_11827_),
    .A4(_13267_),
    .ZN(_13268_));
 INV_X1 _36043_ (.A(\core.keymem.prev_key0_reg[27] ),
    .ZN(_13269_));
 AND4_X1 _36044_ (.A1(_13269_),
    .A2(_13242_),
    .A3(_11860_),
    .A4(_13267_),
    .ZN(_13270_));
 NAND3_X1 _36045_ (.A1(_13269_),
    .A2(_13243_),
    .A3(_11860_),
    .ZN(_13271_));
 NAND3_X1 _36046_ (.A1(\core.keymem.prev_key0_reg[27] ),
    .A2(_13242_),
    .A3(_11860_),
    .ZN(_13272_));
 AOI21_X2 _36047_ (.A(_13267_),
    .B1(_13271_),
    .B2(_13272_),
    .ZN(_13273_));
 AOI21_X1 _36048_ (.A(_11903_),
    .B1(_11891_),
    .B2(_00028_),
    .ZN(_13274_));
 INV_X1 _36049_ (.A(_13274_),
    .ZN(_13275_));
 NOR4_X4 _36050_ (.A1(_13268_),
    .A2(_13270_),
    .A3(_13273_),
    .A4(_13275_),
    .ZN(_13276_));
 BUF_X2 _36051_ (.A(\core.keymem.prev_key1_reg[91] ),
    .Z(_13277_));
 XNOR2_X2 _36052_ (.A(\core.keymem.prev_key1_reg[59] ),
    .B(_13277_),
    .ZN(_13278_));
 XNOR2_X1 _36053_ (.A(\core.keymem.prev_key1_reg[27] ),
    .B(_00027_),
    .ZN(_13279_));
 XNOR2_X1 _36054_ (.A(_13278_),
    .B(_13279_),
    .ZN(_13280_));
 XNOR2_X2 _36055_ (.A(_12167_),
    .B(_13280_),
    .ZN(_13281_));
 OAI22_X4 _36056_ (.A1(_00026_),
    .A2(_11875_),
    .B1(_11814_),
    .B2(_13281_),
    .ZN(_13282_));
 OR2_X2 _36057_ (.A1(_13276_),
    .A2(_13282_),
    .ZN(_13283_));
 CLKBUF_X2 _36058_ (.A(_13283_),
    .Z(_13284_));
 BUF_X4 _36059_ (.A(_12805_),
    .Z(_13285_));
 MUX2_X1 _36060_ (.A(\core.keymem.key_mem[10][27] ),
    .B(_13284_),
    .S(_13285_),
    .Z(_01012_));
 AOI21_X1 _36061_ (.A(_11904_),
    .B1(_12629_),
    .B2(_00031_),
    .ZN(_13286_));
 BUF_X2 _36062_ (.A(\core.keymem.prev_key0_reg[92] ),
    .Z(_13287_));
 NAND3_X1 _36063_ (.A1(_12040_),
    .A2(_13287_),
    .A3(_12915_),
    .ZN(_13288_));
 INV_X1 _36064_ (.A(_13287_),
    .ZN(_13289_));
 NAND3_X1 _36065_ (.A1(_12040_),
    .A2(_13289_),
    .A3(_12919_),
    .ZN(_13290_));
 AOI22_X1 _36066_ (.A1(_11853_),
    .A2(_11854_),
    .B1(_13288_),
    .B2(_13290_),
    .ZN(_13291_));
 NAND3_X1 _36067_ (.A1(_11830_),
    .A2(_13289_),
    .A3(_12915_),
    .ZN(_13292_));
 NAND3_X1 _36068_ (.A1(_11830_),
    .A2(_13287_),
    .A3(_12919_),
    .ZN(_13293_));
 AOI211_X2 _36069_ (.A(_09974_),
    .B(_10008_),
    .C1(_13292_),
    .C2(_13293_),
    .ZN(_13294_));
 NAND4_X1 _36070_ (.A1(_11856_),
    .A2(_12908_),
    .A3(_13289_),
    .A4(_12915_),
    .ZN(_13295_));
 NOR2_X1 _36071_ (.A1(_11830_),
    .A2(_12908_),
    .ZN(_13296_));
 NAND3_X1 _36072_ (.A1(_13287_),
    .A2(_12915_),
    .A3(_13296_),
    .ZN(_13297_));
 AOI22_X1 _36073_ (.A1(_12064_),
    .A2(_12065_),
    .B1(_13295_),
    .B2(_13297_),
    .ZN(_13298_));
 NAND3_X1 _36074_ (.A1(_13289_),
    .A2(_12919_),
    .A3(_13296_),
    .ZN(_13299_));
 NAND4_X1 _36075_ (.A1(_11856_),
    .A2(_12908_),
    .A3(_13287_),
    .A4(_12919_),
    .ZN(_13300_));
 AOI22_X1 _36076_ (.A1(_12064_),
    .A2(_12065_),
    .B1(_13299_),
    .B2(_13300_),
    .ZN(_13301_));
 OR4_X2 _36077_ (.A1(_13291_),
    .A2(_13294_),
    .A3(_13298_),
    .A4(_13301_),
    .ZN(_13302_));
 NOR4_X1 _36078_ (.A1(_11832_),
    .A2(_12908_),
    .A3(_13287_),
    .A4(_12919_),
    .ZN(_13303_));
 NAND2_X1 _36079_ (.A1(_11851_),
    .A2(_12908_),
    .ZN(_13304_));
 NOR3_X1 _36080_ (.A1(_13289_),
    .A2(_12919_),
    .A3(_13304_),
    .ZN(_13305_));
 OAI211_X2 _36081_ (.A(_12064_),
    .B(_12065_),
    .C1(_13303_),
    .C2(_13305_),
    .ZN(_13306_));
 NOR3_X1 _36082_ (.A1(_13287_),
    .A2(_12915_),
    .A3(_13304_),
    .ZN(_13307_));
 NAND3_X1 _36083_ (.A1(_12064_),
    .A2(_12065_),
    .A3(_13307_),
    .ZN(_13308_));
 AND3_X1 _36084_ (.A1(_13287_),
    .A2(_12919_),
    .A3(_13296_),
    .ZN(_13309_));
 NAND3_X1 _36085_ (.A1(_12064_),
    .A2(_12065_),
    .A3(_13309_),
    .ZN(_13310_));
 NAND3_X2 _36086_ (.A1(_13306_),
    .A2(_13308_),
    .A3(_13310_),
    .ZN(_13311_));
 NOR2_X2 _36087_ (.A1(_13302_),
    .A2(_13311_),
    .ZN(_13312_));
 XNOR2_X1 _36088_ (.A(\core.keymem.prev_key0_reg[28] ),
    .B(\core.keymem.prev_key0_reg[60] ),
    .ZN(_13313_));
 XNOR2_X1 _36089_ (.A(_13312_),
    .B(_13313_),
    .ZN(_13314_));
 OAI21_X2 _36090_ (.A(_13286_),
    .B1(_13314_),
    .B2(_12172_),
    .ZN(_13315_));
 NOR2_X2 _36091_ (.A1(_00029_),
    .A2(_11960_),
    .ZN(_13316_));
 CLKBUF_X2 _36092_ (.A(\core.keymem.prev_key1_reg[92] ),
    .Z(_13317_));
 XOR2_X2 _36093_ (.A(\core.keymem.prev_key1_reg[60] ),
    .B(_13317_),
    .Z(_13318_));
 XOR2_X1 _36094_ (.A(_09282_),
    .B(_00030_),
    .Z(_13319_));
 XNOR2_X1 _36095_ (.A(_13318_),
    .B(_13319_),
    .ZN(_13320_));
 XNOR2_X1 _36096_ (.A(_12911_),
    .B(_13320_),
    .ZN(_13321_));
 INV_X1 _36097_ (.A(_13321_),
    .ZN(_13322_));
 AOI21_X2 _36098_ (.A(_13316_),
    .B1(_13322_),
    .B2(_11889_),
    .ZN(_13323_));
 NAND2_X4 _36099_ (.A1(_13315_),
    .A2(_13323_),
    .ZN(_13324_));
 CLKBUF_X2 _36100_ (.A(_13324_),
    .Z(_13325_));
 MUX2_X1 _36101_ (.A(\core.keymem.key_mem[10][28] ),
    .B(_13325_),
    .S(_13285_),
    .Z(_01013_));
 MUX2_X1 _36102_ (.A(_12299_),
    .B(_12303_),
    .S(_12148_),
    .Z(_13326_));
 XNOR2_X2 _36103_ (.A(_12306_),
    .B(_12309_),
    .ZN(_13327_));
 OAI221_X2 _36104_ (.A(_13326_),
    .B1(_13327_),
    .B2(_12241_),
    .C1(_12158_),
    .C2(_00032_),
    .ZN(_13328_));
 BUF_X2 _36105_ (.A(_13328_),
    .Z(_13329_));
 MUX2_X1 _36106_ (.A(\core.keymem.key_mem[10][29] ),
    .B(_13329_),
    .S(_13285_),
    .Z(_01014_));
 NAND2_X1 _36107_ (.A1(\core.keymem.key_mem[10][2] ),
    .A2(_13095_),
    .ZN(_13330_));
 BUF_X8 _36108_ (.A(_12347_),
    .Z(_13331_));
 NAND2_X1 _36109_ (.A1(_13331_),
    .A2(_12318_),
    .ZN(_13332_));
 AOI21_X2 _36110_ (.A(_12951_),
    .B1(_00373_),
    .B2(_12193_),
    .ZN(_13333_));
 AOI22_X4 _36111_ (.A1(_12335_),
    .A2(_12334_),
    .B1(_13332_),
    .B2(_13333_),
    .ZN(_13334_));
 BUF_X2 _36112_ (.A(_13334_),
    .Z(_13335_));
 OAI21_X1 _36113_ (.A(_13330_),
    .B1(_13335_),
    .B2(_12896_),
    .ZN(_01015_));
 CLKBUF_X2 _36114_ (.A(\core.keymem.prev_key1_reg[94] ),
    .Z(_13336_));
 XNOR2_X2 _36115_ (.A(\core.keymem.prev_key1_reg[62] ),
    .B(_13336_),
    .ZN(_13337_));
 XNOR2_X1 _36116_ (.A(_09349_),
    .B(_00036_),
    .ZN(_13338_));
 XNOR2_X1 _36117_ (.A(_13337_),
    .B(_13338_),
    .ZN(_13339_));
 XNOR2_X2 _36118_ (.A(_12195_),
    .B(_13339_),
    .ZN(_13340_));
 OAI22_X4 _36119_ (.A1(_00035_),
    .A2(_11917_),
    .B1(_11814_),
    .B2(_13340_),
    .ZN(_13341_));
 CLKBUF_X2 _36120_ (.A(\core.keymem.prev_key0_reg[62] ),
    .Z(_13342_));
 INV_X1 _36121_ (.A(_13342_),
    .ZN(_13343_));
 BUF_X2 _36122_ (.A(\core.keymem.prev_key0_reg[94] ),
    .Z(_13344_));
 NAND2_X1 _36123_ (.A1(_11830_),
    .A2(_13344_),
    .ZN(_13345_));
 NOR2_X1 _36124_ (.A1(_12200_),
    .A2(_13345_),
    .ZN(_13346_));
 NOR3_X1 _36125_ (.A1(_11856_),
    .A2(_13344_),
    .A3(_12201_),
    .ZN(_13347_));
 OAI22_X1 _36126_ (.A1(_10179_),
    .A2(_10220_),
    .B1(_13346_),
    .B2(_13347_),
    .ZN(_13348_));
 NOR3_X1 _36127_ (.A1(_11851_),
    .A2(_13344_),
    .A3(_12200_),
    .ZN(_13349_));
 NOR2_X1 _36128_ (.A1(_12201_),
    .A2(_13345_),
    .ZN(_13350_));
 OAI211_X2 _36129_ (.A(_09708_),
    .B(_11896_),
    .C1(_13349_),
    .C2(_13350_),
    .ZN(_13351_));
 INV_X2 _36130_ (.A(_12194_),
    .ZN(_13352_));
 NOR4_X1 _36131_ (.A1(_12063_),
    .A2(_13352_),
    .A3(_13344_),
    .A4(_12200_),
    .ZN(_13353_));
 INV_X1 _36132_ (.A(_13344_),
    .ZN(_13354_));
 NOR4_X2 _36133_ (.A1(_12063_),
    .A2(_12194_),
    .A3(_13354_),
    .A4(_12200_),
    .ZN(_13355_));
 OAI22_X2 _36134_ (.A1(_08483_),
    .A2(_09170_),
    .B1(_13353_),
    .B2(_13355_),
    .ZN(_13356_));
 NOR4_X1 _36135_ (.A1(_12063_),
    .A2(_12194_),
    .A3(_13344_),
    .A4(_12201_),
    .ZN(_13357_));
 NOR4_X2 _36136_ (.A1(_12063_),
    .A2(_13352_),
    .A3(_13354_),
    .A4(_12201_),
    .ZN(_13358_));
 OAI22_X2 _36137_ (.A1(_08483_),
    .A2(_09170_),
    .B1(_13357_),
    .B2(_13358_),
    .ZN(_13359_));
 NAND4_X2 _36138_ (.A1(_13348_),
    .A2(_13351_),
    .A3(_13356_),
    .A4(_13359_),
    .ZN(_13360_));
 NAND4_X1 _36139_ (.A1(_11857_),
    .A2(_13352_),
    .A3(_13354_),
    .A4(_12201_),
    .ZN(_13361_));
 NOR2_X1 _36140_ (.A1(_12063_),
    .A2(_13352_),
    .ZN(_13362_));
 NAND3_X1 _36141_ (.A1(_13344_),
    .A2(_12201_),
    .A3(_13362_),
    .ZN(_13363_));
 AOI21_X2 _36142_ (.A(_13170_),
    .B1(_13361_),
    .B2(_13363_),
    .ZN(_13364_));
 NAND3_X1 _36143_ (.A1(_13354_),
    .A2(_12200_),
    .A3(_13362_),
    .ZN(_13365_));
 NAND4_X1 _36144_ (.A1(_11851_),
    .A2(_13352_),
    .A3(_13344_),
    .A4(_12200_),
    .ZN(_13366_));
 AOI21_X2 _36145_ (.A(_13170_),
    .B1(_13365_),
    .B2(_13366_),
    .ZN(_13367_));
 NOR3_X4 _36146_ (.A1(_13360_),
    .A2(_13364_),
    .A3(_13367_),
    .ZN(_13368_));
 AND4_X1 _36147_ (.A1(\core.keymem.prev_key0_reg[30] ),
    .A2(_13343_),
    .A3(_12044_),
    .A4(_13368_),
    .ZN(_13369_));
 INV_X1 _36148_ (.A(\core.keymem.prev_key0_reg[30] ),
    .ZN(_13370_));
 AND4_X1 _36149_ (.A1(_13370_),
    .A2(_13342_),
    .A3(_11827_),
    .A4(_13368_),
    .ZN(_13371_));
 NAND3_X1 _36150_ (.A1(_13370_),
    .A2(_13343_),
    .A3(_11827_),
    .ZN(_13372_));
 NAND3_X1 _36151_ (.A1(\core.keymem.prev_key0_reg[30] ),
    .A2(_13342_),
    .A3(_11827_),
    .ZN(_13373_));
 AOI21_X2 _36152_ (.A(_13368_),
    .B1(_13372_),
    .B2(_13373_),
    .ZN(_13374_));
 AOI21_X2 _36153_ (.A(_11903_),
    .B1(_11891_),
    .B2(_00037_),
    .ZN(_13375_));
 INV_X1 _36154_ (.A(_13375_),
    .ZN(_13376_));
 NOR4_X4 _36155_ (.A1(_13369_),
    .A2(_13371_),
    .A3(_13374_),
    .A4(_13376_),
    .ZN(_13377_));
 OR2_X2 _36156_ (.A1(_13341_),
    .A2(_13377_),
    .ZN(_13378_));
 CLKBUF_X2 _36157_ (.A(_13378_),
    .Z(_13379_));
 MUX2_X1 _36158_ (.A(\core.keymem.key_mem[10][30] ),
    .B(_13379_),
    .S(_13285_),
    .Z(_01016_));
 AOI21_X1 _36159_ (.A(_11903_),
    .B1(_11988_),
    .B2(_00040_),
    .ZN(_13380_));
 INV_X1 _36160_ (.A(_13380_),
    .ZN(_13381_));
 BUF_X2 _36161_ (.A(\core.keymem.prev_key0_reg[95] ),
    .Z(_13382_));
 XNOR2_X1 _36162_ (.A(\core.keymem.prev_key0_reg[63] ),
    .B(_13382_),
    .ZN(_13383_));
 XNOR2_X1 _36163_ (.A(\core.keymem.prev_key0_reg[31] ),
    .B(_13383_),
    .ZN(_13384_));
 XNOR2_X2 _36164_ (.A(_12940_),
    .B(_13384_),
    .ZN(_13385_));
 AOI21_X4 _36165_ (.A(_13381_),
    .B1(_13385_),
    .B2(_11901_),
    .ZN(_13386_));
 CLKBUF_X2 _36166_ (.A(\core.keymem.prev_key1_reg[95] ),
    .Z(_13387_));
 XOR2_X2 _36167_ (.A(\core.keymem.prev_key1_reg[63] ),
    .B(_13387_),
    .Z(_13388_));
 XNOR2_X1 _36168_ (.A(_09268_),
    .B(_00039_),
    .ZN(_13389_));
 XNOR2_X1 _36169_ (.A(_13388_),
    .B(_13389_),
    .ZN(_13390_));
 XNOR2_X2 _36170_ (.A(_12942_),
    .B(_13390_),
    .ZN(_13391_));
 NAND2_X1 _36171_ (.A1(_12027_),
    .A2(_13391_),
    .ZN(_13392_));
 OAI21_X2 _36172_ (.A(_13392_),
    .B1(_12347_),
    .B2(_00038_),
    .ZN(_13393_));
 OR2_X2 _36173_ (.A1(_13386_),
    .A2(_13393_),
    .ZN(_13394_));
 CLKBUF_X2 _36174_ (.A(_13394_),
    .Z(_13395_));
 MUX2_X1 _36175_ (.A(\core.keymem.key_mem[10][31] ),
    .B(_13395_),
    .S(_13285_),
    .Z(_01017_));
 CLKBUF_X2 _36176_ (.A(_12354_),
    .Z(_13396_));
 MUX2_X1 _36177_ (.A(\core.keymem.key_mem[10][32] ),
    .B(_13396_),
    .S(_13285_),
    .Z(_01018_));
 INV_X1 _36178_ (.A(\core.key[33] ),
    .ZN(_13397_));
 AOI21_X1 _36179_ (.A(_11987_),
    .B1(_12629_),
    .B2(_13397_),
    .ZN(_13398_));
 XOR2_X1 _36180_ (.A(_12772_),
    .B(_13119_),
    .Z(_13399_));
 OAI21_X2 _36181_ (.A(_13398_),
    .B1(_13399_),
    .B2(_12172_),
    .ZN(_13400_));
 NAND2_X4 _36182_ (.A1(_12361_),
    .A2(_13400_),
    .ZN(_13401_));
 BUF_X2 _36183_ (.A(_13401_),
    .Z(_13402_));
 MUX2_X1 _36184_ (.A(\core.keymem.key_mem[10][33] ),
    .B(_13402_),
    .S(_13285_),
    .Z(_01019_));
 BUF_X2 _36185_ (.A(_12375_),
    .Z(_13403_));
 MUX2_X1 _36186_ (.A(\core.keymem.key_mem[10][34] ),
    .B(_13403_),
    .S(_13285_),
    .Z(_01020_));
 NAND2_X4 _36187_ (.A1(_12407_),
    .A2(_12412_),
    .ZN(_13404_));
 BUF_X2 _36188_ (.A(_13404_),
    .Z(_13405_));
 MUX2_X1 _36189_ (.A(\core.keymem.key_mem[10][35] ),
    .B(_13405_),
    .S(_13285_),
    .Z(_01021_));
 NAND2_X1 _36190_ (.A1(\core.keymem.key_mem[10][36] ),
    .A2(_13095_),
    .ZN(_13406_));
 CLKBUF_X3 _36191_ (.A(_12422_),
    .Z(_13407_));
 OAI21_X1 _36192_ (.A(_13406_),
    .B1(_12905_),
    .B2(_13407_),
    .ZN(_01022_));
 NAND2_X1 _36193_ (.A1(\core.keymem.key_mem[10][37] ),
    .A2(_13095_),
    .ZN(_13408_));
 OAI21_X1 _36194_ (.A(_13408_),
    .B1(_12905_),
    .B2(_12439_),
    .ZN(_01023_));
 NAND2_X4 _36195_ (.A1(_12462_),
    .A2(_12467_),
    .ZN(_13409_));
 CLKBUF_X2 _36196_ (.A(_13409_),
    .Z(_13410_));
 MUX2_X1 _36197_ (.A(\core.keymem.key_mem[10][38] ),
    .B(_13410_),
    .S(_13285_),
    .Z(_01024_));
 NAND2_X1 _36198_ (.A1(\core.keymem.key_mem[10][39] ),
    .A2(_13095_),
    .ZN(_13411_));
 XNOR2_X2 _36199_ (.A(\core.keymem.prev_key1_reg[39] ),
    .B(_12657_),
    .ZN(_13412_));
 OAI21_X2 _36200_ (.A(_12035_),
    .B1(_13412_),
    .B2(_12156_),
    .ZN(_13413_));
 INV_X1 _36201_ (.A(\core.key[39] ),
    .ZN(_13414_));
 BUF_X4 _36202_ (.A(_11989_),
    .Z(_13415_));
 AOI21_X2 _36203_ (.A(_11847_),
    .B1(_13414_),
    .B2(_13415_),
    .ZN(_13416_));
 CLKBUF_X2 _36204_ (.A(\core.keymem.prev_key0_reg[39] ),
    .Z(_13417_));
 INV_X1 _36205_ (.A(_13417_),
    .ZN(_13418_));
 NOR2_X1 _36206_ (.A1(_13418_),
    .A2(_12653_),
    .ZN(_13419_));
 INV_X1 _36207_ (.A(_12653_),
    .ZN(_13420_));
 NOR2_X1 _36208_ (.A1(_13417_),
    .A2(_13420_),
    .ZN(_13421_));
 OAI221_X2 _36209_ (.A(_11919_),
    .B1(_11921_),
    .B2(_11922_),
    .C1(_13419_),
    .C2(_13421_),
    .ZN(_13422_));
 NOR2_X1 _36210_ (.A1(_13417_),
    .A2(_12653_),
    .ZN(_13423_));
 NOR2_X1 _36211_ (.A1(_13418_),
    .A2(_13420_),
    .ZN(_13424_));
 OAI221_X2 _36212_ (.A(_11918_),
    .B1(_11921_),
    .B2(_11922_),
    .C1(_13423_),
    .C2(_13424_),
    .ZN(_13425_));
 NAND2_X1 _36213_ (.A1(_11919_),
    .A2(_13423_),
    .ZN(_13426_));
 NAND2_X1 _36214_ (.A1(_11919_),
    .A2(_13424_),
    .ZN(_13427_));
 AOI221_X1 _36215_ (.A(_11921_),
    .B1(_13426_),
    .B2(_13427_),
    .C1(_10260_),
    .C2(_12176_),
    .ZN(_13428_));
 NAND3_X1 _36216_ (.A1(_13417_),
    .A2(_13420_),
    .A3(_11918_),
    .ZN(_13429_));
 NAND3_X1 _36217_ (.A1(_13418_),
    .A2(_12653_),
    .A3(_11918_),
    .ZN(_13430_));
 AOI221_X1 _36218_ (.A(_11921_),
    .B1(_13429_),
    .B2(_13430_),
    .C1(_10260_),
    .C2(_12176_),
    .ZN(_13431_));
 NOR2_X1 _36219_ (.A1(_13428_),
    .A2(_13431_),
    .ZN(_13432_));
 NAND4_X4 _36220_ (.A1(_12170_),
    .A2(_13422_),
    .A3(_13425_),
    .A4(_13432_),
    .ZN(_13433_));
 AOI21_X4 _36221_ (.A(_13413_),
    .B1(_13416_),
    .B2(_13433_),
    .ZN(_13434_));
 CLKBUF_X3 _36222_ (.A(_13434_),
    .Z(_13435_));
 OAI21_X1 _36223_ (.A(_13411_),
    .B1(_13435_),
    .B2(_12896_),
    .ZN(_01025_));
 NAND2_X1 _36224_ (.A1(\core.keymem.key_mem[10][3] ),
    .A2(_13095_),
    .ZN(_13436_));
 NAND2_X1 _36225_ (.A1(_00374_),
    .A2(_11841_),
    .ZN(_13437_));
 OAI21_X1 _36226_ (.A(_16228_),
    .B1(_06677_),
    .B2(_13437_),
    .ZN(_13438_));
 INV_X1 _36227_ (.A(_13438_),
    .ZN(_13439_));
 XOR2_X2 _36228_ (.A(\core.keymem.prev_key1_reg[3] ),
    .B(_12411_),
    .Z(_13440_));
 BUF_X4 _36229_ (.A(_12808_),
    .Z(_13441_));
 NOR2_X1 _36230_ (.A1(\core.key[3] ),
    .A2(_11945_),
    .ZN(_13442_));
 XOR2_X2 _36231_ (.A(_12383_),
    .B(_12384_),
    .Z(_13443_));
 XNOR2_X2 _36232_ (.A(\core.keymem.prev_key0_reg[3] ),
    .B(_13443_),
    .ZN(_13444_));
 XOR2_X2 _36233_ (.A(_12796_),
    .B(_13444_),
    .Z(_13445_));
 AOI221_X2 _36234_ (.A(_13442_),
    .B1(_13445_),
    .B2(_11900_),
    .C1(_11812_),
    .C2(_11793_),
    .ZN(_13446_));
 OAI221_X2 _36235_ (.A(_13439_),
    .B1(_13440_),
    .B2(_12263_),
    .C1(_13441_),
    .C2(_13446_),
    .ZN(_13447_));
 CLKBUF_X3 _36236_ (.A(_13447_),
    .Z(_13448_));
 OAI21_X1 _36237_ (.A(_13436_),
    .B1(_13448_),
    .B2(_12896_),
    .ZN(_01026_));
 NAND2_X1 _36238_ (.A1(\core.keymem.key_mem[10][40] ),
    .A2(_13095_),
    .ZN(_13449_));
 OAI21_X1 _36239_ (.A(_11908_),
    .B1(\core.key[40] ),
    .B2(_11900_),
    .ZN(_13450_));
 BUF_X2 _36240_ (.A(\core.keymem.prev_key0_reg[40] ),
    .Z(_13451_));
 XNOR2_X2 _36241_ (.A(_13451_),
    .B(_12666_),
    .ZN(_13452_));
 XNOR2_X2 _36242_ (.A(_12671_),
    .B(_13452_),
    .ZN(_13453_));
 AOI21_X1 _36243_ (.A(_13450_),
    .B1(_13453_),
    .B2(_12333_),
    .ZN(_13454_));
 XNOR2_X2 _36244_ (.A(\core.keymem.prev_key1_reg[40] ),
    .B(_12664_),
    .ZN(_13455_));
 AOI221_X2 _36245_ (.A(_13454_),
    .B1(_11812_),
    .B2(_11793_),
    .C1(_12808_),
    .C2(_13455_),
    .ZN(_13456_));
 CLKBUF_X3 _36246_ (.A(_13456_),
    .Z(_13457_));
 OAI21_X1 _36247_ (.A(_13449_),
    .B1(_13457_),
    .B2(_12896_),
    .ZN(_01027_));
 NOR2_X2 _36248_ (.A1(_00050_),
    .A2(_11960_),
    .ZN(_13458_));
 XNOR2_X1 _36249_ (.A(\core.keymem.prev_key1_reg[41] ),
    .B(_12683_),
    .ZN(_13459_));
 XNOR2_X2 _36250_ (.A(_12684_),
    .B(_13459_),
    .ZN(_13460_));
 AOI21_X2 _36251_ (.A(_13458_),
    .B1(_13460_),
    .B2(_11889_),
    .ZN(_13461_));
 OAI21_X2 _36252_ (.A(_12098_),
    .B1(_12365_),
    .B2(\core.key[41] ),
    .ZN(_13462_));
 XNOR2_X2 _36253_ (.A(\core.keymem.prev_key0_reg[41] ),
    .B(\core.keymem.prev_key0_reg[73] ),
    .ZN(_13463_));
 XNOR2_X1 _36254_ (.A(_12826_),
    .B(_13463_),
    .ZN(_13464_));
 NOR2_X2 _36255_ (.A1(_12345_),
    .A2(_13464_),
    .ZN(_13465_));
 OAI21_X4 _36256_ (.A(_13461_),
    .B1(_13462_),
    .B2(_13465_),
    .ZN(_13466_));
 BUF_X2 _36257_ (.A(_13466_),
    .Z(_13467_));
 BUF_X4 _36258_ (.A(_12805_),
    .Z(_13468_));
 MUX2_X1 _36259_ (.A(\core.keymem.key_mem[10][41] ),
    .B(_13467_),
    .S(_13468_),
    .Z(_01028_));
 INV_X1 _36260_ (.A(_12845_),
    .ZN(_13469_));
 INV_X1 _36261_ (.A(_12846_),
    .ZN(_13470_));
 INV_X1 _36262_ (.A(_11937_),
    .ZN(_13471_));
 NAND3_X1 _36263_ (.A1(_13469_),
    .A2(_13470_),
    .A3(_13471_),
    .ZN(_13472_));
 NAND3_X1 _36264_ (.A1(_12845_),
    .A2(_12846_),
    .A3(_13471_),
    .ZN(_13473_));
 AOI221_X2 _36265_ (.A(_11819_),
    .B1(_11938_),
    .B2(_11942_),
    .C1(_13472_),
    .C2(_13473_),
    .ZN(_13474_));
 NAND3_X1 _36266_ (.A1(_12845_),
    .A2(_13470_),
    .A3(_11937_),
    .ZN(_13475_));
 NAND3_X1 _36267_ (.A1(_13469_),
    .A2(_12846_),
    .A3(_11937_),
    .ZN(_13476_));
 AOI221_X2 _36268_ (.A(_11819_),
    .B1(_11938_),
    .B2(_11942_),
    .C1(_13475_),
    .C2(_13476_),
    .ZN(_13477_));
 NOR3_X2 _36269_ (.A1(_12175_),
    .A2(_07613_),
    .A3(_07641_),
    .ZN(_13478_));
 NAND4_X1 _36270_ (.A1(_12845_),
    .A2(_13470_),
    .A3(_13471_),
    .A4(_11825_),
    .ZN(_13479_));
 NAND4_X1 _36271_ (.A1(_13469_),
    .A2(_12846_),
    .A3(_13471_),
    .A4(_11825_),
    .ZN(_13480_));
 AOI221_X2 _36272_ (.A(_13478_),
    .B1(_13479_),
    .B2(_13480_),
    .C1(_11947_),
    .C2(_12175_),
    .ZN(_13481_));
 NAND4_X1 _36273_ (.A1(_13469_),
    .A2(_13470_),
    .A3(_11937_),
    .A4(_11825_),
    .ZN(_13482_));
 NAND4_X1 _36274_ (.A1(_12845_),
    .A2(_12846_),
    .A3(_11937_),
    .A4(_11825_),
    .ZN(_13483_));
 AOI221_X2 _36275_ (.A(_13478_),
    .B1(_13482_),
    .B2(_13483_),
    .C1(_11947_),
    .C2(_12175_),
    .ZN(_13484_));
 NOR4_X4 _36276_ (.A1(_13474_),
    .A2(_13477_),
    .A3(_13481_),
    .A4(_13484_),
    .ZN(_13485_));
 OR2_X1 _36277_ (.A1(\core.key[42] ),
    .A2(_12149_),
    .ZN(_13486_));
 NAND3_X2 _36278_ (.A1(_12301_),
    .A2(_13485_),
    .A3(_13486_),
    .ZN(_13487_));
 OR2_X1 _36279_ (.A1(_12156_),
    .A2(_12855_),
    .ZN(_13488_));
 NAND3_X4 _36280_ (.A1(_12262_),
    .A2(_13487_),
    .A3(_13488_),
    .ZN(_13489_));
 CLKBUF_X2 _36281_ (.A(_13489_),
    .Z(_13490_));
 MUX2_X1 _36282_ (.A(\core.keymem.key_mem[10][42] ),
    .B(_13490_),
    .S(_13468_),
    .Z(_01029_));
 NAND2_X1 _36283_ (.A1(\core.keymem.key_mem[10][43] ),
    .A2(_13095_),
    .ZN(_13491_));
 OAI21_X2 _36284_ (.A(_12184_),
    .B1(_12887_),
    .B2(_11909_),
    .ZN(_13492_));
 XNOR2_X1 _36285_ (.A(_11962_),
    .B(_12890_),
    .ZN(_13493_));
 MUX2_X2 _36286_ (.A(\core.key[43] ),
    .B(_13493_),
    .S(_12149_),
    .Z(_13494_));
 AOI21_X4 _36287_ (.A(_13492_),
    .B1(_13494_),
    .B2(_06678_),
    .ZN(_13495_));
 CLKBUF_X3 _36288_ (.A(_13495_),
    .Z(_13496_));
 OAI21_X1 _36289_ (.A(_13491_),
    .B1(_13496_),
    .B2(_12896_),
    .ZN(_01030_));
 CLKBUF_X2 _36290_ (.A(_12505_),
    .Z(_13497_));
 MUX2_X1 _36291_ (.A(\core.keymem.key_mem[10][44] ),
    .B(_13497_),
    .S(_13468_),
    .Z(_01031_));
 NAND2_X1 _36292_ (.A1(\core.keymem.key_mem[10][45] ),
    .A2(_13095_),
    .ZN(_13498_));
 XOR2_X1 _36293_ (.A(_12962_),
    .B(_12960_),
    .Z(_13499_));
 AND4_X1 _36294_ (.A1(_12835_),
    .A2(_11848_),
    .A3(_12836_),
    .A4(_13499_),
    .ZN(_13500_));
 XNOR2_X1 _36295_ (.A(_12962_),
    .B(_12960_),
    .ZN(_13501_));
 NOR4_X2 _36296_ (.A1(_12835_),
    .A2(_11891_),
    .A3(_12836_),
    .A4(_13501_),
    .ZN(_13502_));
 AND3_X1 _36297_ (.A1(_12835_),
    .A2(_11826_),
    .A3(_13501_),
    .ZN(_13503_));
 NOR3_X1 _36298_ (.A1(_12835_),
    .A2(_11818_),
    .A3(_13499_),
    .ZN(_13504_));
 MUX2_X1 _36299_ (.A(_13503_),
    .B(_13504_),
    .S(_12836_),
    .Z(_13505_));
 NOR3_X2 _36300_ (.A1(_13500_),
    .A2(_13502_),
    .A3(_13505_),
    .ZN(_13506_));
 OR2_X1 _36301_ (.A1(\core.key[45] ),
    .A2(_11848_),
    .ZN(_13507_));
 AND2_X1 _36302_ (.A1(_06676_),
    .A2(_13507_),
    .ZN(_13508_));
 AOI221_X2 _36303_ (.A(_12680_),
    .B1(_13506_),
    .B2(_13508_),
    .C1(_12969_),
    .C2(_12971_),
    .ZN(_13509_));
 CLKBUF_X3 _36304_ (.A(_13509_),
    .Z(_13510_));
 OAI21_X1 _36305_ (.A(_13498_),
    .B1(_12905_),
    .B2(_13510_),
    .ZN(_01032_));
 BUF_X4 _36306_ (.A(_12815_),
    .Z(_13511_));
 NAND2_X1 _36307_ (.A1(\core.keymem.key_mem[10][46] ),
    .A2(_13511_),
    .ZN(_13512_));
 NOR2_X1 _36308_ (.A1(\core.key[46] ),
    .A2(_11826_),
    .ZN(_13513_));
 XNOR2_X2 _36309_ (.A(_11996_),
    .B(_12980_),
    .ZN(_13514_));
 AOI211_X2 _36310_ (.A(_11811_),
    .B(_13513_),
    .C1(_13514_),
    .C2(_11827_),
    .ZN(_13515_));
 AOI221_X2 _36311_ (.A(_13515_),
    .B1(_11812_),
    .B2(_11793_),
    .C1(_12971_),
    .C2(_12989_),
    .ZN(_13516_));
 CLKBUF_X3 _36312_ (.A(_13516_),
    .Z(_13517_));
 OAI21_X1 _36313_ (.A(_13512_),
    .B1(_13517_),
    .B2(_12896_),
    .ZN(_01033_));
 NAND2_X1 _36314_ (.A1(\core.keymem.key_mem[10][47] ),
    .A2(_13511_),
    .ZN(_13518_));
 OAI21_X1 _36315_ (.A(_13518_),
    .B1(_12905_),
    .B2(_12520_),
    .ZN(_01034_));
 NAND2_X1 _36316_ (.A1(\core.keymem.key_mem[10][48] ),
    .A2(_13511_),
    .ZN(_13519_));
 OAI21_X1 _36317_ (.A(_13519_),
    .B1(_12905_),
    .B2(_12532_),
    .ZN(_01035_));
 NAND2_X1 _36318_ (.A1(\core.keymem.key_mem[10][49] ),
    .A2(_13511_),
    .ZN(_13520_));
 OAI21_X1 _36319_ (.A(_11909_),
    .B1(\core.key[49] ),
    .B2(_11901_),
    .ZN(_13521_));
 XNOR2_X2 _36320_ (.A(_12862_),
    .B(_13031_),
    .ZN(_13522_));
 XOR2_X2 _36321_ (.A(\core.keymem.prev_key0_reg[49] ),
    .B(_13522_),
    .Z(_13523_));
 AOI21_X2 _36322_ (.A(_13521_),
    .B1(_13523_),
    .B2(_12844_),
    .ZN(_13524_));
 INV_X1 _36323_ (.A(\core.keymem.prev_key1_reg[49] ),
    .ZN(_13525_));
 XNOR2_X1 _36324_ (.A(_13525_),
    .B(_13038_),
    .ZN(_13526_));
 OAI21_X2 _36325_ (.A(_12002_),
    .B1(_13526_),
    .B2(_12951_),
    .ZN(_13527_));
 NOR2_X4 _36326_ (.A1(_13524_),
    .A2(_13527_),
    .ZN(_13528_));
 CLKBUF_X3 _36327_ (.A(_13528_),
    .Z(_13529_));
 BUF_X4 _36328_ (.A(_12823_),
    .Z(_13530_));
 OAI21_X1 _36329_ (.A(_13520_),
    .B1(_13529_),
    .B2(_13530_),
    .ZN(_01036_));
 NOR2_X1 _36330_ (.A1(_11908_),
    .A2(_06775_),
    .ZN(_13531_));
 NOR2_X1 _36331_ (.A1(_11908_),
    .A2(_06776_),
    .ZN(_13532_));
 MUX2_X1 _36332_ (.A(_13531_),
    .B(_13532_),
    .S(_12417_),
    .Z(_13533_));
 XOR2_X1 _36333_ (.A(\core.keymem.prev_key0_reg[4] ),
    .B(_12419_),
    .Z(_13534_));
 XNOR2_X1 _36334_ (.A(_11858_),
    .B(_13534_),
    .ZN(_13535_));
 NAND2_X2 _36335_ (.A1(_12170_),
    .A2(_13535_),
    .ZN(_13536_));
 AOI21_X4 _36336_ (.A(_13533_),
    .B1(_13536_),
    .B2(_06678_),
    .ZN(_13537_));
 CLKBUF_X2 _36337_ (.A(_13537_),
    .Z(_13538_));
 MUX2_X1 _36338_ (.A(\core.keymem.key_mem[10][4] ),
    .B(_13538_),
    .S(_13468_),
    .Z(_01037_));
 NOR4_X1 _36339_ (.A1(_13046_),
    .A2(_13048_),
    .A3(_12037_),
    .A4(_11891_),
    .ZN(_13539_));
 NAND2_X1 _36340_ (.A1(_13046_),
    .A2(_13048_),
    .ZN(_13540_));
 NOR3_X1 _36341_ (.A1(_12037_),
    .A2(_11820_),
    .A3(_13540_),
    .ZN(_13541_));
 OAI21_X1 _36342_ (.A(_12042_),
    .B1(_13539_),
    .B2(_13541_),
    .ZN(_13542_));
 NOR3_X1 _36343_ (.A1(_13051_),
    .A2(_13048_),
    .A3(_12038_),
    .ZN(_13543_));
 NOR3_X1 _36344_ (.A1(_13046_),
    .A2(_13056_),
    .A3(_12038_),
    .ZN(_13544_));
 OAI221_X2 _36345_ (.A(_11828_),
    .B1(_13043_),
    .B2(_12041_),
    .C1(_13543_),
    .C2(_13544_),
    .ZN(_13545_));
 NAND4_X1 _36346_ (.A1(_13046_),
    .A2(_13056_),
    .A3(_12038_),
    .A4(_11826_),
    .ZN(_13546_));
 NAND4_X1 _36347_ (.A1(_13051_),
    .A2(_13048_),
    .A3(_12038_),
    .A4(_11825_),
    .ZN(_13547_));
 AOI221_X2 _36348_ (.A(_13043_),
    .B1(_13546_),
    .B2(_13547_),
    .C1(_12046_),
    .C2(_12175_),
    .ZN(_13548_));
 NAND4_X1 _36349_ (.A1(_13051_),
    .A2(_13056_),
    .A3(_12037_),
    .A4(_11826_),
    .ZN(_13549_));
 NOR3_X1 _36350_ (.A1(_13043_),
    .A2(_12041_),
    .A3(_13549_),
    .ZN(_13550_));
 OR3_X1 _36351_ (.A1(_12038_),
    .A2(_11818_),
    .A3(_13540_),
    .ZN(_13551_));
 NOR3_X1 _36352_ (.A1(_13043_),
    .A2(_12041_),
    .A3(_13551_),
    .ZN(_13552_));
 NOR3_X1 _36353_ (.A1(_13548_),
    .A2(_13550_),
    .A3(_13552_),
    .ZN(_13553_));
 NAND3_X2 _36354_ (.A1(_13542_),
    .A2(_13545_),
    .A3(_13553_),
    .ZN(_13554_));
 OAI21_X1 _36355_ (.A(_06677_),
    .B1(\core.key[50] ),
    .B2(_12333_),
    .ZN(_13555_));
 OAI221_X2 _36356_ (.A(_12185_),
    .B1(_13554_),
    .B2(_13555_),
    .C1(_13091_),
    .C2(_12301_),
    .ZN(_13556_));
 BUF_X2 _36357_ (.A(_13556_),
    .Z(_13557_));
 MUX2_X1 _36358_ (.A(\core.keymem.key_mem[10][50] ),
    .B(_13557_),
    .S(_13468_),
    .Z(_01038_));
 NOR2_X2 _36359_ (.A1(_00060_),
    .A2(_11960_),
    .ZN(_13558_));
 AOI21_X2 _36360_ (.A(_13558_),
    .B1(_13101_),
    .B2(_11889_),
    .ZN(_13559_));
 OAI21_X2 _36361_ (.A(_11936_),
    .B1(_12170_),
    .B2(\core.key[51] ),
    .ZN(_13560_));
 XOR2_X2 _36362_ (.A(_12052_),
    .B(_13104_),
    .Z(_13561_));
 NOR2_X2 _36363_ (.A1(_12172_),
    .A2(_13561_),
    .ZN(_13562_));
 OAI21_X4 _36364_ (.A(_13559_),
    .B1(_13560_),
    .B2(_13562_),
    .ZN(_13563_));
 CLKBUF_X2 _36365_ (.A(_13563_),
    .Z(_13564_));
 MUX2_X1 _36366_ (.A(\core.keymem.key_mem[10][51] ),
    .B(_13564_),
    .S(_13468_),
    .Z(_01039_));
 NAND2_X1 _36367_ (.A1(\core.keymem.key_mem[10][52] ),
    .A2(_13511_),
    .ZN(_13565_));
 OAI21_X1 _36368_ (.A(_13565_),
    .B1(_12905_),
    .B2(_12568_),
    .ZN(_01040_));
 NAND2_X1 _36369_ (.A1(\core.keymem.key_mem[10][53] ),
    .A2(_13511_),
    .ZN(_13566_));
 OAI21_X1 _36370_ (.A(_13566_),
    .B1(_12905_),
    .B2(_12584_),
    .ZN(_01041_));
 NAND2_X1 _36371_ (.A1(\core.keymem.key_mem[10][54] ),
    .A2(_13511_),
    .ZN(_13567_));
 OAI21_X1 _36372_ (.A(_11823_),
    .B1(_12149_),
    .B2(\core.key[54] ),
    .ZN(_13568_));
 XNOR2_X1 _36373_ (.A(_13175_),
    .B(_12738_),
    .ZN(_13569_));
 AOI21_X2 _36374_ (.A(_13568_),
    .B1(_13569_),
    .B2(_12365_),
    .ZN(_13570_));
 NOR2_X2 _36375_ (.A1(_00063_),
    .A2(_12347_),
    .ZN(_13571_));
 XNOR2_X2 _36376_ (.A(_13158_),
    .B(_12729_),
    .ZN(_13572_));
 NOR2_X2 _36377_ (.A1(_12001_),
    .A2(_13572_),
    .ZN(_13573_));
 NOR3_X4 _36378_ (.A1(_13570_),
    .A2(_13571_),
    .A3(_13573_),
    .ZN(_13574_));
 CLKBUF_X3 _36379_ (.A(_13574_),
    .Z(_13575_));
 OAI21_X1 _36380_ (.A(_13567_),
    .B1(_13575_),
    .B2(_13530_),
    .ZN(_01042_));
 NOR2_X1 _36381_ (.A1(_11909_),
    .A2(_12266_),
    .ZN(_13576_));
 NOR2_X1 _36382_ (.A1(_12193_),
    .A2(_13576_),
    .ZN(_13577_));
 OR2_X1 _36383_ (.A1(\core.key[55] ),
    .A2(_11828_),
    .ZN(_13578_));
 OAI21_X2 _36384_ (.A(_13578_),
    .B1(_12259_),
    .B2(_11997_),
    .ZN(_13579_));
 OAI21_X4 _36385_ (.A(_13577_),
    .B1(_13579_),
    .B2(_12292_),
    .ZN(_13580_));
 BUF_X2 _36386_ (.A(_13580_),
    .Z(_13581_));
 MUX2_X1 _36387_ (.A(\core.keymem.key_mem[10][55] ),
    .B(_13581_),
    .S(_13468_),
    .Z(_01043_));
 XNOR2_X2 _36388_ (.A(_12122_),
    .B(_13205_),
    .ZN(_13582_));
 AND2_X2 _36389_ (.A1(_12027_),
    .A2(_13582_),
    .ZN(_13583_));
 NOR2_X1 _36390_ (.A1(_00066_),
    .A2(_12044_),
    .ZN(_13584_));
 OR2_X1 _36391_ (.A1(_11987_),
    .A2(_13584_),
    .ZN(_13585_));
 XOR2_X2 _36392_ (.A(\core.keymem.prev_key0_reg[56] ),
    .B(_13201_),
    .Z(_13586_));
 AOI21_X4 _36393_ (.A(_13585_),
    .B1(_13586_),
    .B2(_12170_),
    .ZN(_13587_));
 NOR2_X4 _36394_ (.A1(_13583_),
    .A2(_13587_),
    .ZN(_13588_));
 CLKBUF_X2 _36395_ (.A(_13588_),
    .Z(_13589_));
 MUX2_X1 _36396_ (.A(\core.keymem.key_mem[10][56] ),
    .B(_13589_),
    .S(_13468_),
    .Z(_01044_));
 AND4_X1 _36397_ (.A1(_12130_),
    .A2(_12131_),
    .A3(_12137_),
    .A4(_12141_),
    .ZN(_13590_));
 AND3_X1 _36398_ (.A1(_12143_),
    .A2(_12144_),
    .A3(_12145_),
    .ZN(_13591_));
 INV_X1 _36399_ (.A(_13223_),
    .ZN(_13592_));
 NAND2_X1 _36400_ (.A1(_13221_),
    .A2(_13592_),
    .ZN(_13593_));
 INV_X1 _36401_ (.A(_13221_),
    .ZN(_13594_));
 NAND2_X1 _36402_ (.A1(_13594_),
    .A2(_13223_),
    .ZN(_13595_));
 AOI221_X2 _36403_ (.A(_11891_),
    .B1(_13590_),
    .B2(_13591_),
    .C1(_13593_),
    .C2(_13595_),
    .ZN(_13596_));
 NAND3_X1 _36404_ (.A1(_13594_),
    .A2(_13592_),
    .A3(_11848_),
    .ZN(_13597_));
 NAND3_X1 _36405_ (.A1(_13221_),
    .A2(_13223_),
    .A3(_11848_),
    .ZN(_13598_));
 AOI211_X2 _36406_ (.A(_12142_),
    .B(_12146_),
    .C1(_13597_),
    .C2(_13598_),
    .ZN(_13599_));
 NOR2_X1 _36407_ (.A1(_00068_),
    .A2(_11828_),
    .ZN(_13600_));
 NOR3_X4 _36408_ (.A1(_13596_),
    .A2(_13599_),
    .A3(_13600_),
    .ZN(_13601_));
 XOR2_X2 _36409_ (.A(_12155_),
    .B(_13214_),
    .Z(_13602_));
 AOI22_X4 _36410_ (.A1(_12335_),
    .A2(_13601_),
    .B1(_13602_),
    .B2(_12028_),
    .ZN(_13603_));
 CLKBUF_X2 _36411_ (.A(_13603_),
    .Z(_13604_));
 MUX2_X1 _36412_ (.A(\core.keymem.key_mem[10][57] ),
    .B(_13604_),
    .S(_13468_),
    .Z(_01045_));
 INV_X1 _36413_ (.A(_00070_),
    .ZN(_13605_));
 XNOR2_X1 _36414_ (.A(_12280_),
    .B(_12901_),
    .ZN(_13606_));
 OAI221_X2 _36415_ (.A(_12184_),
    .B1(_12966_),
    .B2(_13605_),
    .C1(_13606_),
    .C2(_11909_),
    .ZN(_13607_));
 XNOR2_X2 _36416_ (.A(_12898_),
    .B(_13235_),
    .ZN(_13608_));
 XNOR2_X2 _36417_ (.A(\core.keymem.prev_key0_reg[58] ),
    .B(_13608_),
    .ZN(_13609_));
 AOI21_X4 _36418_ (.A(_13607_),
    .B1(_13609_),
    .B2(_13176_),
    .ZN(_13610_));
 BUF_X2 _36419_ (.A(_13610_),
    .Z(_13611_));
 MUX2_X1 _36420_ (.A(\core.keymem.key_mem[10][58] ),
    .B(_13611_),
    .S(_13468_),
    .Z(_01046_));
 AND3_X1 _36421_ (.A1(_06676_),
    .A2(_00072_),
    .A3(_11988_),
    .ZN(_13612_));
 XNOR2_X2 _36422_ (.A(_13242_),
    .B(_13267_),
    .ZN(_13613_));
 XNOR2_X2 _36423_ (.A(_12168_),
    .B(_13278_),
    .ZN(_13614_));
 AOI221_X2 _36424_ (.A(_13612_),
    .B1(_13613_),
    .B2(_13176_),
    .C1(_12971_),
    .C2(_13614_),
    .ZN(_13615_));
 CLKBUF_X2 _36425_ (.A(_13615_),
    .Z(_13616_));
 BUF_X4 _36426_ (.A(_12805_),
    .Z(_13617_));
 MUX2_X1 _36427_ (.A(\core.keymem.key_mem[10][59] ),
    .B(_13616_),
    .S(_13617_),
    .Z(_01047_));
 MUX2_X1 _36428_ (.A(\core.keymem.key_mem[10][5] ),
    .B(_12606_),
    .S(_13617_),
    .Z(_01048_));
 AND3_X1 _36429_ (.A1(_06676_),
    .A2(_00074_),
    .A3(_11988_),
    .ZN(_13618_));
 XNOR2_X1 _36430_ (.A(\core.keymem.prev_key0_reg[60] ),
    .B(_13312_),
    .ZN(_13619_));
 XOR2_X2 _36431_ (.A(_12912_),
    .B(_13318_),
    .Z(_13620_));
 AOI221_X2 _36432_ (.A(_13618_),
    .B1(_13619_),
    .B2(_13176_),
    .C1(_12971_),
    .C2(_13620_),
    .ZN(_13621_));
 BUF_X2 _36433_ (.A(_13621_),
    .Z(_13622_));
 MUX2_X1 _36434_ (.A(\core.keymem.key_mem[10][60] ),
    .B(_13622_),
    .S(_13617_),
    .Z(_01049_));
 XNOR2_X2 _36435_ (.A(_12930_),
    .B(_12295_),
    .ZN(_13623_));
 NOR2_X2 _36436_ (.A1(_12705_),
    .A2(_13623_),
    .ZN(_13624_));
 OAI21_X2 _36437_ (.A(_11822_),
    .B1(_11827_),
    .B2(_00076_),
    .ZN(_13625_));
 NOR2_X1 _36438_ (.A1(_12308_),
    .A2(_13625_),
    .ZN(_13626_));
 AND2_X1 _36439_ (.A1(_12306_),
    .A2(_13626_),
    .ZN(_13627_));
 INV_X1 _36440_ (.A(_12308_),
    .ZN(_13628_));
 NOR3_X4 _36441_ (.A1(_12306_),
    .A2(_13628_),
    .A3(_13625_),
    .ZN(_13629_));
 NOR2_X2 _36442_ (.A1(_11901_),
    .A2(_13625_),
    .ZN(_13630_));
 NOR4_X4 _36443_ (.A1(_13624_),
    .A2(_13627_),
    .A3(_13629_),
    .A4(_13630_),
    .ZN(_13631_));
 CLKBUF_X2 _36444_ (.A(_13631_),
    .Z(_13632_));
 MUX2_X1 _36445_ (.A(\core.keymem.key_mem[10][61] ),
    .B(_13632_),
    .S(_13617_),
    .Z(_01050_));
 XNOR2_X1 _36446_ (.A(_13342_),
    .B(_13368_),
    .ZN(_13633_));
 MUX2_X1 _36447_ (.A(_00078_),
    .B(_13633_),
    .S(_11945_),
    .Z(_13634_));
 XNOR2_X2 _36448_ (.A(_12196_),
    .B(_13337_),
    .ZN(_13635_));
 OAI222_X2 _36449_ (.A1(_00077_),
    .A2(_12002_),
    .B1(_11904_),
    .B2(_13634_),
    .C1(_13635_),
    .C2(_12705_),
    .ZN(_13636_));
 BUF_X2 _36450_ (.A(_13636_),
    .Z(_13637_));
 MUX2_X1 _36451_ (.A(\core.keymem.key_mem[10][62] ),
    .B(_13637_),
    .S(_13617_),
    .Z(_01051_));
 NAND2_X1 _36452_ (.A1(_12148_),
    .A2(_00080_),
    .ZN(_13638_));
 XNOR2_X2 _36453_ (.A(_12943_),
    .B(_13388_),
    .ZN(_13639_));
 OAI221_X2 _36454_ (.A(_12184_),
    .B1(_11901_),
    .B2(_13638_),
    .C1(_13639_),
    .C2(_11909_),
    .ZN(_13640_));
 INV_X1 _36455_ (.A(_12936_),
    .ZN(_13641_));
 NAND3_X1 _36456_ (.A1(_12175_),
    .A2(_13382_),
    .A3(_13641_),
    .ZN(_13642_));
 NOR2_X1 _36457_ (.A1(_11832_),
    .A2(_13382_),
    .ZN(_13643_));
 NAND2_X1 _36458_ (.A1(_12936_),
    .A2(_13643_),
    .ZN(_13644_));
 AOI21_X2 _36459_ (.A(_12942_),
    .B1(_13642_),
    .B2(_13644_),
    .ZN(_13645_));
 NAND2_X1 _36460_ (.A1(_13641_),
    .A2(_13643_),
    .ZN(_13646_));
 NAND3_X1 _36461_ (.A1(_12175_),
    .A2(_13382_),
    .A3(_12936_),
    .ZN(_13647_));
 AOI21_X2 _36462_ (.A(_12938_),
    .B1(_13646_),
    .B2(_13647_),
    .ZN(_13648_));
 INV_X1 _36463_ (.A(_13382_),
    .ZN(_13649_));
 NAND3_X1 _36464_ (.A1(_12917_),
    .A2(_13649_),
    .A3(_13641_),
    .ZN(_13650_));
 NAND3_X1 _36465_ (.A1(_12917_),
    .A2(_13382_),
    .A3(_12936_),
    .ZN(_13651_));
 AOI21_X2 _36466_ (.A(_10260_),
    .B1(_13650_),
    .B2(_13651_),
    .ZN(_13652_));
 NAND3_X1 _36467_ (.A1(_12917_),
    .A2(_13382_),
    .A3(_13641_),
    .ZN(_13653_));
 NAND3_X1 _36468_ (.A1(_12917_),
    .A2(_13649_),
    .A3(_12936_),
    .ZN(_13654_));
 AOI21_X2 _36469_ (.A(_11910_),
    .B1(_13653_),
    .B2(_13654_),
    .ZN(_13655_));
 NOR4_X4 _36470_ (.A1(_13645_),
    .A2(_13648_),
    .A3(_13652_),
    .A4(_13655_),
    .ZN(_13656_));
 XOR2_X2 _36471_ (.A(\core.keymem.prev_key0_reg[63] ),
    .B(_13656_),
    .Z(_13657_));
 AOI21_X4 _36472_ (.A(_13640_),
    .B1(_13657_),
    .B2(_13176_),
    .ZN(_13658_));
 BUF_X2 _36473_ (.A(_13658_),
    .Z(_13659_));
 MUX2_X1 _36474_ (.A(\core.keymem.key_mem[10][63] ),
    .B(_13659_),
    .S(_13617_),
    .Z(_01052_));
 MUX2_X1 _36475_ (.A(\core.keymem.key_mem[10][64] ),
    .B(_12622_),
    .S(_13617_),
    .Z(_01053_));
 NAND2_X1 _36476_ (.A1(\core.keymem.key_mem[10][65] ),
    .A2(_13511_),
    .ZN(_13660_));
 AOI21_X1 _36477_ (.A(_12148_),
    .B1(_00082_),
    .B2(_11799_),
    .ZN(_13661_));
 INV_X1 _36478_ (.A(\core.keymem.prev_key1_reg[65] ),
    .ZN(_13662_));
 XNOR2_X1 _36479_ (.A(_13662_),
    .B(_12358_),
    .ZN(_13663_));
 OAI21_X1 _36480_ (.A(_13661_),
    .B1(_13663_),
    .B2(_12680_),
    .ZN(_13664_));
 INV_X1 _36481_ (.A(_13664_),
    .ZN(_13665_));
 INV_X1 _36482_ (.A(_00082_),
    .ZN(_13666_));
 OAI21_X1 _36483_ (.A(_12349_),
    .B1(_13666_),
    .B2(_11885_),
    .ZN(_13667_));
 AND2_X1 _36484_ (.A1(\core.key[65] ),
    .A2(_11988_),
    .ZN(_13668_));
 XNOR2_X1 _36485_ (.A(_13118_),
    .B(_12772_),
    .ZN(_13669_));
 AOI21_X2 _36486_ (.A(_13668_),
    .B1(_13669_),
    .B2(_12333_),
    .ZN(_13670_));
 AOI21_X2 _36487_ (.A(_13667_),
    .B1(_13670_),
    .B2(_12035_),
    .ZN(_13671_));
 OAI21_X4 _36488_ (.A(_16229_),
    .B1(_13665_),
    .B2(_13671_),
    .ZN(_13672_));
 CLKBUF_X3 _36489_ (.A(_13672_),
    .Z(_13673_));
 OAI21_X1 _36490_ (.A(_13660_),
    .B1(_13673_),
    .B2(_13530_),
    .ZN(_01054_));
 NAND2_X1 _36491_ (.A1(\core.key[66] ),
    .A2(_11892_),
    .ZN(_13674_));
 NAND2_X1 _36492_ (.A1(_12148_),
    .A2(_13674_),
    .ZN(_13675_));
 XNOR2_X2 _36493_ (.A(_12325_),
    .B(_12324_),
    .ZN(_13676_));
 AOI21_X4 _36494_ (.A(_13675_),
    .B1(_13676_),
    .B2(_12365_),
    .ZN(_13677_));
 NAND2_X1 _36495_ (.A1(_11916_),
    .A2(_12316_),
    .ZN(_13678_));
 NAND2_X2 _36496_ (.A1(_12184_),
    .A2(_13678_),
    .ZN(_13679_));
 OAI22_X4 _36497_ (.A1(_00083_),
    .A2(_13331_),
    .B1(_13677_),
    .B2(_13679_),
    .ZN(_13680_));
 CLKBUF_X2 _36498_ (.A(_13680_),
    .Z(_13681_));
 MUX2_X1 _36499_ (.A(\core.keymem.key_mem[10][66] ),
    .B(_13681_),
    .S(_13617_),
    .Z(_01055_));
 NAND2_X1 _36500_ (.A1(\core.keymem.key_mem[10][67] ),
    .A2(_13511_),
    .ZN(_13682_));
 NAND2_X1 _36501_ (.A1(\core.key[67] ),
    .A2(_12345_),
    .ZN(_13683_));
 OAI21_X1 _36502_ (.A(_12384_),
    .B1(_12794_),
    .B2(_12795_),
    .ZN(_13684_));
 OR3_X1 _36503_ (.A1(_12384_),
    .A2(_12794_),
    .A3(_12795_),
    .ZN(_13685_));
 NAND3_X2 _36504_ (.A1(_11901_),
    .A2(_13684_),
    .A3(_13685_),
    .ZN(_13686_));
 AOI21_X4 _36505_ (.A(_11904_),
    .B1(_13683_),
    .B2(_13686_),
    .ZN(_13687_));
 OAI22_X4 _36506_ (.A1(_00084_),
    .A2(_12035_),
    .B1(_12705_),
    .B2(_12410_),
    .ZN(_13688_));
 NOR2_X2 _36507_ (.A1(_13687_),
    .A2(_13688_),
    .ZN(_13689_));
 CLKBUF_X3 _36508_ (.A(_13689_),
    .Z(_13690_));
 OAI21_X1 _36509_ (.A(_13682_),
    .B1(_13690_),
    .B2(_13530_),
    .ZN(_01056_));
 NAND2_X1 _36510_ (.A1(\core.keymem.key_mem[10][68] ),
    .A2(_13511_),
    .ZN(_13691_));
 OAI21_X1 _36511_ (.A(_13691_),
    .B1(_12824_),
    .B2(_12635_),
    .ZN(_01057_));
 BUF_X4 _36512_ (.A(_12815_),
    .Z(_13692_));
 NAND2_X1 _36513_ (.A1(\core.keymem.key_mem[10][69] ),
    .A2(_13692_),
    .ZN(_13693_));
 NAND2_X1 _36514_ (.A1(_00086_),
    .A2(_11800_),
    .ZN(_13694_));
 INV_X1 _36515_ (.A(\core.key[69] ),
    .ZN(_13695_));
 OAI21_X1 _36516_ (.A(_12098_),
    .B1(_11901_),
    .B2(_13695_),
    .ZN(_13696_));
 AND2_X1 _36517_ (.A1(_12099_),
    .A2(_12429_),
    .ZN(_13697_));
 XOR2_X2 _36518_ (.A(_12434_),
    .B(_12433_),
    .Z(_13698_));
 OAI221_X2 _36519_ (.A(_13694_),
    .B1(_13696_),
    .B2(_13697_),
    .C1(_12263_),
    .C2(_13698_),
    .ZN(_13699_));
 CLKBUF_X3 _36520_ (.A(_13699_),
    .Z(_13700_));
 OAI21_X1 _36521_ (.A(_13693_),
    .B1(_13700_),
    .B2(_13530_),
    .ZN(_01058_));
 OR3_X1 _36522_ (.A1(\core.keymem.prev_key0_reg[6] ),
    .A2(_11820_),
    .A3(_11903_),
    .ZN(_13701_));
 NAND3_X1 _36523_ (.A1(\core.keymem.prev_key0_reg[6] ),
    .A2(_11900_),
    .A3(_11823_),
    .ZN(_13702_));
 MUX2_X2 _36524_ (.A(_13701_),
    .B(_13702_),
    .S(_12460_),
    .Z(_13703_));
 AND3_X1 _36525_ (.A1(\core.key[6] ),
    .A2(_11892_),
    .A3(_11823_),
    .ZN(_13704_));
 XOR2_X1 _36526_ (.A(_06823_),
    .B(_00379_),
    .Z(_13705_));
 XNOR2_X1 _36527_ (.A(_12465_),
    .B(_13705_),
    .ZN(_13706_));
 XNOR2_X1 _36528_ (.A(_10221_),
    .B(_13706_),
    .ZN(_13707_));
 AOI21_X2 _36529_ (.A(_13704_),
    .B1(_13707_),
    .B2(_12027_),
    .ZN(_13708_));
 OR2_X2 _36530_ (.A1(_00378_),
    .A2(_11875_),
    .ZN(_13709_));
 NAND3_X4 _36531_ (.A1(_13703_),
    .A2(_13708_),
    .A3(_13709_),
    .ZN(_13710_));
 BUF_X2 _36532_ (.A(_13710_),
    .Z(_13711_));
 MUX2_X1 _36533_ (.A(\core.keymem.key_mem[10][6] ),
    .B(_13711_),
    .S(_13617_),
    .Z(_01059_));
 NAND2_X2 _36534_ (.A1(_12645_),
    .A2(_12647_),
    .ZN(_13712_));
 CLKBUF_X2 _36535_ (.A(_13712_),
    .Z(_13713_));
 MUX2_X1 _36536_ (.A(\core.keymem.key_mem[10][70] ),
    .B(_13713_),
    .S(_13617_),
    .Z(_01060_));
 NAND2_X1 _36537_ (.A1(\core.keymem.key_mem[10][71] ),
    .A2(_13692_),
    .ZN(_13714_));
 OAI21_X1 _36538_ (.A(_13714_),
    .B1(_12824_),
    .B2(_12659_),
    .ZN(_01061_));
 NAND2_X1 _36539_ (.A1(\core.keymem.key_mem[10][72] ),
    .A2(_13692_),
    .ZN(_13715_));
 CLKBUF_X3 _36540_ (.A(_12673_),
    .Z(_13716_));
 OAI21_X1 _36541_ (.A(_13715_),
    .B1(_12824_),
    .B2(_13716_),
    .ZN(_01062_));
 NAND2_X1 _36542_ (.A1(\core.keymem.key_mem[10][73] ),
    .A2(_13692_),
    .ZN(_13717_));
 OAI21_X1 _36543_ (.A(_13717_),
    .B1(_12824_),
    .B2(_12688_),
    .ZN(_01063_));
 NAND2_X1 _36544_ (.A1(\core.keymem.key_mem[10][74] ),
    .A2(_13692_),
    .ZN(_13718_));
 OAI21_X1 _36545_ (.A(_12971_),
    .B1(_12689_),
    .B2(_12347_),
    .ZN(_13719_));
 BUF_X4 _36546_ (.A(_11875_),
    .Z(_13720_));
 AOI21_X2 _36547_ (.A(_13719_),
    .B1(_12854_),
    .B2(_13720_),
    .ZN(_13721_));
 NAND2_X1 _36548_ (.A1(\core.key[74] ),
    .A2(_12172_),
    .ZN(_13722_));
 XNOR2_X2 _36549_ (.A(_12846_),
    .B(_11944_),
    .ZN(_13723_));
 OAI21_X2 _36550_ (.A(_13722_),
    .B1(_13723_),
    .B2(_13415_),
    .ZN(_13724_));
 AOI21_X4 _36551_ (.A(_13721_),
    .B1(_13724_),
    .B2(_12335_),
    .ZN(_13725_));
 CLKBUF_X3 _36552_ (.A(_13725_),
    .Z(_13726_));
 OAI21_X1 _36553_ (.A(_13718_),
    .B1(_13726_),
    .B2(_13530_),
    .ZN(_01064_));
 NAND2_X1 _36554_ (.A1(\core.keymem.key_mem[10][75] ),
    .A2(_13692_),
    .ZN(_13727_));
 NAND2_X1 _36555_ (.A1(_12971_),
    .A2(_12886_),
    .ZN(_13728_));
 XOR2_X1 _36556_ (.A(_11962_),
    .B(_12889_),
    .Z(_13729_));
 MUX2_X1 _36557_ (.A(\core.key[75] ),
    .B(_13729_),
    .S(_11945_),
    .Z(_13730_));
 OAI21_X1 _36558_ (.A(_13728_),
    .B1(_13730_),
    .B2(_11847_),
    .ZN(_13731_));
 MUX2_X2 _36559_ (.A(_00092_),
    .B(_13731_),
    .S(_12002_),
    .Z(_13732_));
 CLKBUF_X3 _36560_ (.A(_13732_),
    .Z(_13733_));
 OAI21_X1 _36561_ (.A(_13727_),
    .B1(_13733_),
    .B2(_13530_),
    .ZN(_01065_));
 NAND2_X1 _36562_ (.A1(_00093_),
    .A2(_12680_),
    .ZN(_13734_));
 NOR2_X1 _36563_ (.A1(_11908_),
    .A2(_12502_),
    .ZN(_13735_));
 NAND2_X1 _36564_ (.A1(\core.key[76] ),
    .A2(_12092_),
    .ZN(_13736_));
 AOI21_X1 _36565_ (.A(_13735_),
    .B1(_13736_),
    .B2(_12349_),
    .ZN(_13737_));
 OAI21_X2 _36566_ (.A(_13734_),
    .B1(_13737_),
    .B2(_12779_),
    .ZN(_13738_));
 XNOR2_X2 _36567_ (.A(_12485_),
    .B(_11974_),
    .ZN(_13739_));
 OAI21_X4 _36568_ (.A(_13738_),
    .B1(_13739_),
    .B2(_12241_),
    .ZN(_13740_));
 BUF_X2 _36569_ (.A(_13740_),
    .Z(_13741_));
 BUF_X4 _36570_ (.A(_12805_),
    .Z(_13742_));
 MUX2_X1 _36571_ (.A(\core.keymem.key_mem[10][76] ),
    .B(_13741_),
    .S(_13742_),
    .Z(_01066_));
 NOR2_X2 _36572_ (.A1(_00094_),
    .A2(_12347_),
    .ZN(_13743_));
 INV_X1 _36573_ (.A(_13743_),
    .ZN(_13744_));
 XNOR2_X1 _36574_ (.A(_12836_),
    .B(_12961_),
    .ZN(_13745_));
 NOR2_X2 _36575_ (.A1(_11989_),
    .A2(_13745_),
    .ZN(_13746_));
 INV_X1 _36576_ (.A(\core.key[77] ),
    .ZN(_13747_));
 OAI21_X2 _36577_ (.A(_12349_),
    .B1(_13747_),
    .B2(_12099_),
    .ZN(_13748_));
 OAI22_X4 _36578_ (.A1(_12951_),
    .A2(_12968_),
    .B1(_13746_),
    .B2(_13748_),
    .ZN(_13749_));
 NAND2_X2 _36579_ (.A1(_13744_),
    .A2(_13749_),
    .ZN(_13750_));
 CLKBUF_X2 _36580_ (.A(_13750_),
    .Z(_13751_));
 MUX2_X1 _36581_ (.A(\core.keymem.key_mem[10][77] ),
    .B(_13751_),
    .S(_13742_),
    .Z(_01067_));
 NAND2_X1 _36582_ (.A1(\core.keymem.key_mem[10][78] ),
    .A2(_13692_),
    .ZN(_13752_));
 OAI21_X1 _36583_ (.A(_13752_),
    .B1(_12824_),
    .B2(_12708_),
    .ZN(_01068_));
 AOI21_X1 _36584_ (.A(_11916_),
    .B1(\core.key[79] ),
    .B2(_11989_),
    .ZN(_13753_));
 OAI21_X2 _36585_ (.A(_13753_),
    .B1(_12512_),
    .B2(_11997_),
    .ZN(_13754_));
 NOR2_X1 _36586_ (.A1(_12349_),
    .A2(_12516_),
    .ZN(_13755_));
 NOR2_X2 _36587_ (.A1(_11842_),
    .A2(_13755_),
    .ZN(_13756_));
 AND3_X2 _36588_ (.A1(_16229_),
    .A2(_13754_),
    .A3(_13756_),
    .ZN(_13757_));
 CLKBUF_X2 _36589_ (.A(_13757_),
    .Z(_13758_));
 MUX2_X1 _36590_ (.A(\core.keymem.key_mem[10][79] ),
    .B(_13758_),
    .S(_13742_),
    .Z(_01069_));
 NAND2_X1 _36591_ (.A1(\core.keymem.key_mem[10][7] ),
    .A2(_13692_),
    .ZN(_13759_));
 XNOR2_X1 _36592_ (.A(_06756_),
    .B(_13412_),
    .ZN(_13760_));
 OAI22_X2 _36593_ (.A1(_00380_),
    .A2(_12035_),
    .B1(_12705_),
    .B2(_13760_),
    .ZN(_13761_));
 XOR2_X1 _36594_ (.A(_13417_),
    .B(_12653_),
    .Z(_13762_));
 XNOR2_X1 _36595_ (.A(\core.keymem.prev_key0_reg[7] ),
    .B(_13762_),
    .ZN(_13763_));
 XNOR2_X1 _36596_ (.A(_11924_),
    .B(_13763_),
    .ZN(_13764_));
 MUX2_X2 _36597_ (.A(\core.key[7] ),
    .B(_13764_),
    .S(_12099_),
    .Z(_13765_));
 AOI21_X4 _36598_ (.A(_13761_),
    .B1(_13765_),
    .B2(_12335_),
    .ZN(_13766_));
 CLKBUF_X3 _36599_ (.A(_13766_),
    .Z(_13767_));
 OAI21_X1 _36600_ (.A(_13759_),
    .B1(_13767_),
    .B2(_13530_),
    .ZN(_01070_));
 OR2_X2 _36601_ (.A1(_12712_),
    .A2(_12715_),
    .ZN(_13768_));
 CLKBUF_X2 _36602_ (.A(_13768_),
    .Z(_13769_));
 MUX2_X1 _36603_ (.A(\core.keymem.key_mem[10][80] ),
    .B(_13769_),
    .S(_13742_),
    .Z(_01071_));
 NAND2_X1 _36604_ (.A1(\core.keymem.key_mem[10][81] ),
    .A2(_13692_),
    .ZN(_13770_));
 INV_X1 _36605_ (.A(\core.key[81] ),
    .ZN(_13771_));
 MUX2_X1 _36606_ (.A(_13771_),
    .B(_13522_),
    .S(_11925_),
    .Z(_13772_));
 MUX2_X1 _36607_ (.A(_13038_),
    .B(_13772_),
    .S(_12349_),
    .Z(_13773_));
 MUX2_X2 _36608_ (.A(_00098_),
    .B(_13773_),
    .S(_12002_),
    .Z(_13774_));
 CLKBUF_X3 _36609_ (.A(_13774_),
    .Z(_13775_));
 OAI21_X1 _36610_ (.A(_13770_),
    .B1(_13775_),
    .B2(_13530_),
    .ZN(_01072_));
 NAND2_X1 _36611_ (.A1(\core.keymem.key_mem[10][82] ),
    .A2(_13692_),
    .ZN(_13776_));
 AOI22_X2 _36612_ (.A1(_00099_),
    .A2(_11800_),
    .B1(_12028_),
    .B2(_13090_),
    .ZN(_13777_));
 NAND2_X1 _36613_ (.A1(\core.key[82] ),
    .A2(_11997_),
    .ZN(_13778_));
 NAND2_X1 _36614_ (.A1(_11936_),
    .A2(_13778_),
    .ZN(_13779_));
 XNOR2_X2 _36615_ (.A(_13056_),
    .B(_12043_),
    .ZN(_13780_));
 NOR2_X1 _36616_ (.A1(_13415_),
    .A2(_13780_),
    .ZN(_13781_));
 OAI21_X4 _36617_ (.A(_13777_),
    .B1(_13779_),
    .B2(_13781_),
    .ZN(_13782_));
 CLKBUF_X3 _36618_ (.A(_13782_),
    .Z(_13783_));
 OAI21_X1 _36619_ (.A(_13776_),
    .B1(_13783_),
    .B2(_13530_),
    .ZN(_01073_));
 NAND2_X1 _36620_ (.A1(\core.keymem.key_mem[10][83] ),
    .A2(_12823_),
    .ZN(_13784_));
 NOR2_X2 _36621_ (.A1(_00100_),
    .A2(_12184_),
    .ZN(_13785_));
 AOI21_X1 _36622_ (.A(_11866_),
    .B1(\core.key[83] ),
    .B2(_12629_),
    .ZN(_13786_));
 XOR2_X2 _36623_ (.A(\core.keymem.prev_key0_reg[83] ),
    .B(_12052_),
    .Z(_13787_));
 OAI21_X2 _36624_ (.A(_13786_),
    .B1(_13787_),
    .B2(_13415_),
    .ZN(_13788_));
 AOI21_X2 _36625_ (.A(_11842_),
    .B1(_13100_),
    .B2(_11847_),
    .ZN(_13789_));
 AOI21_X4 _36626_ (.A(_13785_),
    .B1(_13788_),
    .B2(_13789_),
    .ZN(_13790_));
 CLKBUF_X3 _36627_ (.A(_13790_),
    .Z(_13791_));
 OAI21_X1 _36628_ (.A(_13784_),
    .B1(_13791_),
    .B2(_12816_),
    .ZN(_01074_));
 NAND2_X1 _36629_ (.A1(\core.keymem.key_mem[10][84] ),
    .A2(_12823_),
    .ZN(_13792_));
 OAI21_X1 _36630_ (.A(_13792_),
    .B1(_12824_),
    .B2(_12725_),
    .ZN(_01075_));
 NOR2_X4 _36631_ (.A1(_00102_),
    .A2(_11917_),
    .ZN(_13793_));
 NAND3_X1 _36632_ (.A1(_12148_),
    .A2(\core.key[85] ),
    .A3(_12101_),
    .ZN(_13794_));
 XNOR2_X1 _36633_ (.A(_12579_),
    .B(_12578_),
    .ZN(_13795_));
 OAI221_X2 _36634_ (.A(_13794_),
    .B1(_12959_),
    .B2(_12573_),
    .C1(_06677_),
    .C2(_13795_),
    .ZN(_13796_));
 OR2_X2 _36635_ (.A1(_13793_),
    .A2(_13796_),
    .ZN(_13797_));
 BUF_X2 _36636_ (.A(_13797_),
    .Z(_13798_));
 MUX2_X1 _36637_ (.A(\core.keymem.key_mem[10][85] ),
    .B(_13798_),
    .S(_13742_),
    .Z(_01076_));
 MUX2_X1 _36638_ (.A(\core.keymem.key_mem[10][86] ),
    .B(_12741_),
    .S(_13742_),
    .Z(_01077_));
 NOR2_X1 _36639_ (.A1(_12951_),
    .A2(_12265_),
    .ZN(_13799_));
 AND2_X1 _36640_ (.A1(\core.key[87] ),
    .A2(_12092_),
    .ZN(_13800_));
 XNOR2_X2 _36641_ (.A(_12244_),
    .B(_12091_),
    .ZN(_13801_));
 AOI21_X4 _36642_ (.A(_13800_),
    .B1(_13801_),
    .B2(_12170_),
    .ZN(_13802_));
 AOI21_X4 _36643_ (.A(_13799_),
    .B1(_13802_),
    .B2(_06678_),
    .ZN(_13803_));
 CLKBUF_X2 _36644_ (.A(_13803_),
    .Z(_13804_));
 MUX2_X1 _36645_ (.A(\core.keymem.key_mem[10][87] ),
    .B(_13804_),
    .S(_13742_),
    .Z(_01078_));
 NOR2_X1 _36646_ (.A1(_11997_),
    .A2(_13201_),
    .ZN(_13805_));
 NAND2_X1 _36647_ (.A1(_00106_),
    .A2(_12101_),
    .ZN(_13806_));
 NAND2_X1 _36648_ (.A1(_06677_),
    .A2(_13806_),
    .ZN(_13807_));
 XOR2_X2 _36649_ (.A(_13204_),
    .B(_12122_),
    .Z(_13808_));
 OAI221_X2 _36650_ (.A(_12834_),
    .B1(_13805_),
    .B2(_13807_),
    .C1(_13808_),
    .C2(_12301_),
    .ZN(_13809_));
 BUF_X2 _36651_ (.A(_13809_),
    .Z(_13810_));
 MUX2_X1 _36652_ (.A(\core.keymem.key_mem[10][88] ),
    .B(_13810_),
    .S(_13742_),
    .Z(_01079_));
 OAI21_X1 _36653_ (.A(_13592_),
    .B1(_12142_),
    .B2(_12146_),
    .ZN(_13811_));
 NAND3_X1 _36654_ (.A1(_13223_),
    .A2(_13590_),
    .A3(_13591_),
    .ZN(_13812_));
 AOI21_X2 _36655_ (.A(_11989_),
    .B1(_13811_),
    .B2(_13812_),
    .ZN(_13813_));
 AND2_X1 _36656_ (.A1(_00108_),
    .A2(_11820_),
    .ZN(_13814_));
 OR2_X1 _36657_ (.A1(_11846_),
    .A2(_13814_),
    .ZN(_13815_));
 XNOR2_X1 _36658_ (.A(_13213_),
    .B(_12155_),
    .ZN(_13816_));
 OAI221_X2 _36659_ (.A(_13331_),
    .B1(_13813_),
    .B2(_13815_),
    .C1(_13816_),
    .C2(_12951_),
    .ZN(_13817_));
 BUF_X2 _36660_ (.A(_13817_),
    .Z(_13818_));
 MUX2_X1 _36661_ (.A(\core.keymem.key_mem[10][89] ),
    .B(_13818_),
    .S(_13742_),
    .Z(_01080_));
 AOI21_X1 _36662_ (.A(_11987_),
    .B1(_12101_),
    .B2(\core.key[8] ),
    .ZN(_13819_));
 INV_X1 _36663_ (.A(_13451_),
    .ZN(_13820_));
 MUX2_X2 _36664_ (.A(_07222_),
    .B(_10613_),
    .S(_11832_),
    .Z(_13821_));
 BUF_X2 _36665_ (.A(\core.keymem.prev_key0_reg[8] ),
    .Z(_13822_));
 INV_X1 _36666_ (.A(_13822_),
    .ZN(_13823_));
 NAND2_X1 _36667_ (.A1(_12666_),
    .A2(_12667_),
    .ZN(_13824_));
 NOR3_X1 _36668_ (.A1(_13823_),
    .A2(_11988_),
    .A3(_13824_),
    .ZN(_13825_));
 NAND3_X1 _36669_ (.A1(_13820_),
    .A2(_13821_),
    .A3(_13825_),
    .ZN(_13826_));
 OR3_X1 _36670_ (.A1(_13822_),
    .A2(_12667_),
    .A3(_13452_),
    .ZN(_13827_));
 NAND2_X1 _36671_ (.A1(_13822_),
    .A2(_13820_),
    .ZN(_13828_));
 OR3_X1 _36672_ (.A1(_12666_),
    .A2(_12667_),
    .A3(_13828_),
    .ZN(_13829_));
 AOI21_X1 _36673_ (.A(_12670_),
    .B1(_13827_),
    .B2(_13829_),
    .ZN(_13830_));
 NAND2_X1 _36674_ (.A1(_13822_),
    .A2(_13451_),
    .ZN(_13831_));
 NOR3_X1 _36675_ (.A1(_13821_),
    .A2(_13824_),
    .A3(_13831_),
    .ZN(_13832_));
 OAI21_X1 _36676_ (.A(_12099_),
    .B1(_13830_),
    .B2(_13832_),
    .ZN(_13833_));
 AND3_X1 _36677_ (.A1(_13819_),
    .A2(_13826_),
    .A3(_13833_),
    .ZN(_13834_));
 OR2_X1 _36678_ (.A1(_13822_),
    .A2(_13820_),
    .ZN(_13835_));
 INV_X1 _36679_ (.A(_12667_),
    .ZN(_13836_));
 NAND2_X1 _36680_ (.A1(_12666_),
    .A2(_13836_),
    .ZN(_13837_));
 OR2_X1 _36681_ (.A1(_12666_),
    .A2(_13836_),
    .ZN(_13838_));
 AOI221_X2 _36682_ (.A(_13821_),
    .B1(_13828_),
    .B2(_13835_),
    .C1(_13837_),
    .C2(_13838_),
    .ZN(_13839_));
 AOI21_X1 _36683_ (.A(_13831_),
    .B1(_13837_),
    .B2(_13838_),
    .ZN(_13840_));
 NOR3_X1 _36684_ (.A1(_13822_),
    .A2(_13451_),
    .A3(_13824_),
    .ZN(_13841_));
 MUX2_X1 _36685_ (.A(_13840_),
    .B(_13841_),
    .S(_12670_),
    .Z(_13842_));
 OR2_X1 _36686_ (.A1(_13839_),
    .A2(_13842_),
    .ZN(_13843_));
 NOR4_X1 _36687_ (.A1(_13822_),
    .A2(_13451_),
    .A3(_12666_),
    .A4(_12667_),
    .ZN(_13844_));
 NOR3_X1 _36688_ (.A1(_12666_),
    .A2(_12667_),
    .A3(_13831_),
    .ZN(_13845_));
 OAI21_X1 _36689_ (.A(_12670_),
    .B1(_13844_),
    .B2(_13845_),
    .ZN(_13846_));
 NOR3_X1 _36690_ (.A1(_13822_),
    .A2(_13451_),
    .A3(_13838_),
    .ZN(_13847_));
 NOR2_X1 _36691_ (.A1(_13824_),
    .A2(_13835_),
    .ZN(_13848_));
 OAI21_X1 _36692_ (.A(_13821_),
    .B1(_13847_),
    .B2(_13848_),
    .ZN(_13849_));
 NAND2_X1 _36693_ (.A1(_13846_),
    .A2(_13849_),
    .ZN(_13850_));
 OAI21_X2 _36694_ (.A(_12170_),
    .B1(_13843_),
    .B2(_13850_),
    .ZN(_13851_));
 XNOR2_X2 _36695_ (.A(_07261_),
    .B(_13455_),
    .ZN(_13852_));
 AOI22_X4 _36696_ (.A1(_13834_),
    .A2(_13851_),
    .B1(_13852_),
    .B2(_12028_),
    .ZN(_13853_));
 CLKBUF_X2 _36697_ (.A(_13853_),
    .Z(_13854_));
 MUX2_X1 _36698_ (.A(\core.keymem.key_mem[10][8] ),
    .B(_13854_),
    .S(_13742_),
    .Z(_01081_));
 XNOR2_X1 _36699_ (.A(_12279_),
    .B(_12901_),
    .ZN(_13855_));
 AOI21_X2 _36700_ (.A(_12779_),
    .B1(_13855_),
    .B2(_12808_),
    .ZN(_13856_));
 NAND2_X1 _36701_ (.A1(_00110_),
    .A2(_12629_),
    .ZN(_13857_));
 OAI21_X2 _36702_ (.A(_13857_),
    .B1(_13608_),
    .B2(_12345_),
    .ZN(_13858_));
 OAI21_X4 _36703_ (.A(_13856_),
    .B1(_13858_),
    .B2(_12292_),
    .ZN(_13859_));
 BUF_X2 _36704_ (.A(_13859_),
    .Z(_13860_));
 MUX2_X1 _36705_ (.A(\core.keymem.key_mem[10][90] ),
    .B(_13860_),
    .S(_12806_),
    .Z(_01082_));
 NAND2_X1 _36706_ (.A1(\core.keymem.key_mem[10][91] ),
    .A2(_12823_),
    .ZN(_13861_));
 INV_X1 _36707_ (.A(_13277_),
    .ZN(_13862_));
 XNOR2_X1 _36708_ (.A(_13862_),
    .B(_12168_),
    .ZN(_13863_));
 NAND2_X2 _36709_ (.A1(_12028_),
    .A2(_13863_),
    .ZN(_13864_));
 NAND2_X1 _36710_ (.A1(_00112_),
    .A2(_12345_),
    .ZN(_13865_));
 NOR2_X1 _36711_ (.A1(_12786_),
    .A2(_13865_),
    .ZN(_13866_));
 NOR2_X2 _36712_ (.A1(_12241_),
    .A2(_13267_),
    .ZN(_13867_));
 NOR2_X4 _36713_ (.A1(_13866_),
    .A2(_13867_),
    .ZN(_13868_));
 NAND2_X2 _36714_ (.A1(_13864_),
    .A2(_13868_),
    .ZN(_13869_));
 CLKBUF_X3 _36715_ (.A(_13869_),
    .Z(_13870_));
 OAI21_X1 _36716_ (.A(_13861_),
    .B1(_13870_),
    .B2(_12816_),
    .ZN(_01083_));
 NAND2_X1 _36717_ (.A1(\core.keymem.key_mem[10][92] ),
    .A2(_12823_),
    .ZN(_13871_));
 OAI21_X2 _36718_ (.A(_11901_),
    .B1(_13302_),
    .B2(_13311_),
    .ZN(_13872_));
 NAND2_X1 _36719_ (.A1(_00114_),
    .A2(_12345_),
    .ZN(_13873_));
 AND3_X2 _36720_ (.A1(_12301_),
    .A2(_13872_),
    .A3(_13873_),
    .ZN(_13874_));
 BUF_X4 _36721_ (.A(_12184_),
    .Z(_13875_));
 INV_X2 _36722_ (.A(_13317_),
    .ZN(_13876_));
 XNOR2_X1 _36723_ (.A(_13876_),
    .B(_12912_),
    .ZN(_13877_));
 OAI21_X2 _36724_ (.A(_13875_),
    .B1(_13877_),
    .B2(_06678_),
    .ZN(_13878_));
 NOR2_X2 _36725_ (.A1(_13874_),
    .A2(_13878_),
    .ZN(_13879_));
 CLKBUF_X3 _36726_ (.A(_13879_),
    .Z(_13880_));
 OAI21_X1 _36727_ (.A(_13871_),
    .B1(_13880_),
    .B2(_12816_),
    .ZN(_01084_));
 XNOR2_X2 _36728_ (.A(_12294_),
    .B(_12930_),
    .ZN(_13881_));
 AOI21_X2 _36729_ (.A(_12193_),
    .B1(_13881_),
    .B2(_12808_),
    .ZN(_13882_));
 NAND2_X1 _36730_ (.A1(_00116_),
    .A2(_12172_),
    .ZN(_13883_));
 NAND2_X1 _36731_ (.A1(_06678_),
    .A2(_13883_),
    .ZN(_13884_));
 NOR2_X1 _36732_ (.A1(_12307_),
    .A2(_12092_),
    .ZN(_13885_));
 AND2_X1 _36733_ (.A1(_12307_),
    .A2(_11945_),
    .ZN(_13886_));
 MUX2_X2 _36734_ (.A(_13885_),
    .B(_13886_),
    .S(_12306_),
    .Z(_13887_));
 OAI21_X4 _36735_ (.A(_13882_),
    .B1(_13884_),
    .B2(_13887_),
    .ZN(_13888_));
 BUF_X2 _36736_ (.A(_13888_),
    .Z(_13889_));
 MUX2_X1 _36737_ (.A(\core.keymem.key_mem[10][93] ),
    .B(_13889_),
    .S(_12806_),
    .Z(_01085_));
 NOR2_X1 _36738_ (.A1(_12629_),
    .A2(_13368_),
    .ZN(_13890_));
 NAND2_X1 _36739_ (.A1(_00118_),
    .A2(_12101_),
    .ZN(_13891_));
 NAND2_X1 _36740_ (.A1(_06677_),
    .A2(_13891_),
    .ZN(_13892_));
 INV_X1 _36741_ (.A(_13336_),
    .ZN(_13893_));
 XNOR2_X1 _36742_ (.A(_13893_),
    .B(_12196_),
    .ZN(_13894_));
 OAI221_X2 _36743_ (.A(_12834_),
    .B1(_13890_),
    .B2(_13892_),
    .C1(_13894_),
    .C2(_12301_),
    .ZN(_13895_));
 BUF_X2 _36744_ (.A(_13895_),
    .Z(_13896_));
 MUX2_X1 _36745_ (.A(\core.keymem.key_mem[10][94] ),
    .B(_13896_),
    .S(_12806_),
    .Z(_01086_));
 AND2_X1 _36746_ (.A1(_12099_),
    .A2(_13656_),
    .ZN(_13897_));
 NAND2_X1 _36747_ (.A1(_00120_),
    .A2(_12101_),
    .ZN(_13898_));
 NAND2_X1 _36748_ (.A1(_06677_),
    .A2(_13898_),
    .ZN(_13899_));
 INV_X1 _36749_ (.A(_13387_),
    .ZN(_13900_));
 XNOR2_X1 _36750_ (.A(_13900_),
    .B(_12943_),
    .ZN(_13901_));
 OAI221_X2 _36751_ (.A(_12834_),
    .B1(_13897_),
    .B2(_13899_),
    .C1(_13901_),
    .C2(_12301_),
    .ZN(_13902_));
 BUF_X2 _36752_ (.A(_13902_),
    .Z(_13903_));
 MUX2_X1 _36753_ (.A(\core.keymem.key_mem[10][95] ),
    .B(_13903_),
    .S(_12806_),
    .Z(_01087_));
 MUX2_X1 _36754_ (.A(\core.key[96] ),
    .B(_11835_),
    .S(_11860_),
    .Z(_13904_));
 MUX2_X1 _36755_ (.A(_12351_),
    .B(_13904_),
    .S(_12148_),
    .Z(_13905_));
 OR2_X1 _36756_ (.A1(_12860_),
    .A2(_13905_),
    .ZN(_13906_));
 CLKBUF_X2 _36757_ (.A(_13906_),
    .Z(_13907_));
 MUX2_X1 _36758_ (.A(\core.keymem.key_mem[10][96] ),
    .B(_13907_),
    .S(_12806_),
    .Z(_01088_));
 NAND2_X1 _36759_ (.A1(\core.keymem.key_mem[10][97] ),
    .A2(_12823_),
    .ZN(_13908_));
 OAI21_X1 _36760_ (.A(_13908_),
    .B1(_12824_),
    .B2(_12777_),
    .ZN(_01089_));
 NAND2_X1 _36761_ (.A1(\core.keymem.key_mem[10][98] ),
    .A2(_12823_),
    .ZN(_13909_));
 CLKBUF_X3 _36762_ (.A(_12787_),
    .Z(_13910_));
 OAI21_X1 _36763_ (.A(_13909_),
    .B1(_12824_),
    .B2(_13910_),
    .ZN(_01090_));
 MUX2_X1 _36764_ (.A(\core.keymem.key_mem[10][99] ),
    .B(_12800_),
    .S(_12806_),
    .Z(_01091_));
 NOR2_X1 _36765_ (.A1(\core.key[9] ),
    .A2(_11827_),
    .ZN(_13911_));
 NAND2_X1 _36766_ (.A1(_11908_),
    .A2(_13911_),
    .ZN(_13912_));
 NAND2_X1 _36767_ (.A1(_11960_),
    .A2(_13912_),
    .ZN(_13913_));
 XNOR2_X1 _36768_ (.A(\core.keymem.prev_key0_reg[9] ),
    .B(_13463_),
    .ZN(_13914_));
 XNOR2_X1 _36769_ (.A(_12678_),
    .B(_13914_),
    .ZN(_13915_));
 NOR2_X1 _36770_ (.A1(_12959_),
    .A2(_13915_),
    .ZN(_13916_));
 XNOR2_X1 _36771_ (.A(\core.keymem.prev_key1_reg[9] ),
    .B(_13460_),
    .ZN(_13917_));
 AOI211_X2 _36772_ (.A(_13913_),
    .B(_13916_),
    .C1(_12971_),
    .C2(_13917_),
    .ZN(_13918_));
 BUF_X2 _36773_ (.A(_13918_),
    .Z(_13919_));
 MUX2_X1 _36774_ (.A(\core.keymem.key_mem[10][9] ),
    .B(_13919_),
    .S(_12806_),
    .Z(_01092_));
 BUF_X2 _36775_ (.A(_22112_),
    .Z(_13920_));
 NAND2_X4 _36776_ (.A1(_16222_),
    .A2(_13920_),
    .ZN(_13921_));
 NOR2_X4 _36777_ (.A1(_12803_),
    .A2(_13921_),
    .ZN(_13922_));
 BUF_X4 _36778_ (.A(_13922_),
    .Z(_13923_));
 BUF_X4 _36779_ (.A(_13923_),
    .Z(_13924_));
 MUX2_X1 _36780_ (.A(\core.keymem.key_mem[11][0] ),
    .B(_11844_),
    .S(_13924_),
    .Z(_01093_));
 MUX2_X1 _36781_ (.A(\core.keymem.key_mem[11][100] ),
    .B(_11873_),
    .S(_13924_),
    .Z(_01094_));
 MUX2_X1 _36782_ (.A(\core.keymem.key_mem[11][101] ),
    .B(_12813_),
    .S(_13924_),
    .Z(_01095_));
 MUX2_X1 _36783_ (.A(\core.keymem.key_mem[11][102] ),
    .B(_11906_),
    .S(_13924_),
    .Z(_01096_));
 MUX2_X1 _36784_ (.A(\core.keymem.key_mem[11][103] ),
    .B(_11929_),
    .S(_13924_),
    .Z(_01097_));
 OR2_X1 _36785_ (.A1(_12803_),
    .A2(_13921_),
    .ZN(_13925_));
 CLKBUF_X3 _36786_ (.A(_13925_),
    .Z(_13926_));
 BUF_X4 _36787_ (.A(_13926_),
    .Z(_13927_));
 NAND2_X1 _36788_ (.A1(\core.keymem.key_mem[11][104] ),
    .A2(_13927_),
    .ZN(_13928_));
 BUF_X4 _36789_ (.A(_13926_),
    .Z(_13929_));
 BUF_X4 _36790_ (.A(_13929_),
    .Z(_13930_));
 OAI21_X1 _36791_ (.A(_13928_),
    .B1(_13930_),
    .B2(_12822_),
    .ZN(_01098_));
 MUX2_X1 _36792_ (.A(\core.keymem.key_mem[11][105] ),
    .B(_12830_),
    .S(_13924_),
    .Z(_01099_));
 BUF_X4 _36793_ (.A(_13923_),
    .Z(_13931_));
 MUX2_X1 _36794_ (.A(\core.keymem.key_mem[11][106] ),
    .B(_12832_),
    .S(_13931_),
    .Z(_01100_));
 MUX2_X1 _36795_ (.A(\core.keymem.key_mem[11][107] ),
    .B(_11967_),
    .S(_13931_),
    .Z(_01101_));
 MUX2_X1 _36796_ (.A(\core.keymem.key_mem[11][108] ),
    .B(_11981_),
    .S(_13931_),
    .Z(_01102_));
 MUX2_X1 _36797_ (.A(\core.keymem.key_mem[11][109] ),
    .B(_12842_),
    .S(_13931_),
    .Z(_01103_));
 NAND2_X1 _36798_ (.A1(\core.keymem.key_mem[11][10] ),
    .A2(_13927_),
    .ZN(_13932_));
 OAI21_X1 _36799_ (.A(_13932_),
    .B1(_13930_),
    .B2(_12858_),
    .ZN(_01104_));
 MUX2_X1 _36800_ (.A(\core.keymem.key_mem[11][110] ),
    .B(_12859_),
    .S(_13931_),
    .Z(_01105_));
 MUX2_X1 _36801_ (.A(\core.keymem.key_mem[11][111] ),
    .B(_12017_),
    .S(_13931_),
    .Z(_01106_));
 MUX2_X1 _36802_ (.A(\core.keymem.key_mem[11][112] ),
    .B(_12031_),
    .S(_13931_),
    .Z(_01107_));
 MUX2_X1 _36803_ (.A(\core.keymem.key_mem[11][113] ),
    .B(_12868_),
    .S(_13931_),
    .Z(_01108_));
 MUX2_X1 _36804_ (.A(\core.keymem.key_mem[11][114] ),
    .B(_12869_),
    .S(_13931_),
    .Z(_01109_));
 MUX2_X1 _36805_ (.A(\core.keymem.key_mem[11][115] ),
    .B(_12059_),
    .S(_13931_),
    .Z(_01110_));
 BUF_X4 _36806_ (.A(_13923_),
    .Z(_13933_));
 MUX2_X1 _36807_ (.A(\core.keymem.key_mem[11][116] ),
    .B(_12077_),
    .S(_13933_),
    .Z(_01111_));
 MUX2_X1 _36808_ (.A(\core.keymem.key_mem[11][117] ),
    .B(_12877_),
    .S(_13933_),
    .Z(_01112_));
 MUX2_X1 _36809_ (.A(\core.keymem.key_mem[11][118] ),
    .B(_12882_),
    .S(_13933_),
    .Z(_01113_));
 MUX2_X1 _36810_ (.A(\core.keymem.key_mem[11][119] ),
    .B(_12096_),
    .S(_13933_),
    .Z(_01114_));
 NAND2_X1 _36811_ (.A1(\core.keymem.key_mem[11][11] ),
    .A2(_13927_),
    .ZN(_13934_));
 OAI21_X1 _36812_ (.A(_13934_),
    .B1(_13930_),
    .B2(_12895_),
    .ZN(_01115_));
 MUX2_X1 _36813_ (.A(\core.keymem.key_mem[11][120] ),
    .B(_12124_),
    .S(_13933_),
    .Z(_01116_));
 MUX2_X1 _36814_ (.A(\core.keymem.key_mem[11][121] ),
    .B(_12160_),
    .S(_13933_),
    .Z(_01117_));
 MUX2_X1 _36815_ (.A(\core.keymem.key_mem[11][122] ),
    .B(_12903_),
    .S(_13933_),
    .Z(_01118_));
 NAND2_X1 _36816_ (.A1(\core.keymem.key_mem[11][123] ),
    .A2(_13927_),
    .ZN(_13935_));
 OAI21_X1 _36817_ (.A(_13935_),
    .B1(_13930_),
    .B2(_12182_),
    .ZN(_01119_));
 NAND2_X1 _36818_ (.A1(\core.keymem.key_mem[11][124] ),
    .A2(_13927_),
    .ZN(_13936_));
 OAI21_X1 _36819_ (.A(_13936_),
    .B1(_13930_),
    .B2(_12926_),
    .ZN(_01120_));
 MUX2_X1 _36820_ (.A(\core.keymem.key_mem[11][125] ),
    .B(_12932_),
    .S(_13933_),
    .Z(_01121_));
 NAND2_X1 _36821_ (.A1(\core.keymem.key_mem[11][126] ),
    .A2(_13927_),
    .ZN(_13937_));
 OAI21_X1 _36822_ (.A(_13937_),
    .B1(_13930_),
    .B2(_12207_),
    .ZN(_01122_));
 MUX2_X1 _36823_ (.A(\core.keymem.key_mem[11][127] ),
    .B(_12945_),
    .S(_13933_),
    .Z(_01123_));
 MUX2_X1 _36824_ (.A(\core.keymem.key_mem[11][12] ),
    .B(_12958_),
    .S(_13933_),
    .Z(_01124_));
 BUF_X8 _36825_ (.A(_13922_),
    .Z(_13938_));
 MUX2_X1 _36826_ (.A(\core.keymem.key_mem[11][13] ),
    .B(_12974_),
    .S(_13938_),
    .Z(_01125_));
 NOR2_X1 _36827_ (.A1(\core.keymem.key_mem[11][14] ),
    .A2(_13924_),
    .ZN(_13939_));
 AOI21_X1 _36828_ (.A(_13939_),
    .B1(_13924_),
    .B2(_13007_),
    .ZN(_01126_));
 MUX2_X1 _36829_ (.A(\core.keymem.key_mem[11][15] ),
    .B(_13017_),
    .S(_13938_),
    .Z(_01127_));
 MUX2_X1 _36830_ (.A(\core.keymem.key_mem[11][16] ),
    .B(_13029_),
    .S(_13938_),
    .Z(_01128_));
 NAND2_X1 _36831_ (.A1(\core.keymem.key_mem[11][17] ),
    .A2(_13927_),
    .ZN(_13940_));
 OAI21_X1 _36832_ (.A(_13940_),
    .B1(_13930_),
    .B2(_13042_),
    .ZN(_01129_));
 MUX2_X1 _36833_ (.A(\core.keymem.key_mem[11][18] ),
    .B(_13094_),
    .S(_13938_),
    .Z(_01130_));
 BUF_X4 _36834_ (.A(_13926_),
    .Z(_13941_));
 NAND2_X1 _36835_ (.A1(\core.keymem.key_mem[11][19] ),
    .A2(_13941_),
    .ZN(_13942_));
 OAI21_X1 _36836_ (.A(_13942_),
    .B1(_13930_),
    .B2(_13109_),
    .ZN(_01131_));
 MUX2_X1 _36837_ (.A(\core.keymem.key_mem[11][1] ),
    .B(_13134_),
    .S(_13938_),
    .Z(_01132_));
 MUX2_X1 _36838_ (.A(\core.keymem.key_mem[11][20] ),
    .B(_13146_),
    .S(_13938_),
    .Z(_01133_));
 MUX2_X1 _36839_ (.A(\core.keymem.key_mem[11][21] ),
    .B(_13155_),
    .S(_13938_),
    .Z(_01134_));
 NOR2_X1 _36840_ (.A1(\core.keymem.key_mem[11][22] ),
    .A2(_13924_),
    .ZN(_13943_));
 AOI21_X1 _36841_ (.A(_13943_),
    .B1(_13924_),
    .B2(_13191_),
    .ZN(_01135_));
 MUX2_X1 _36842_ (.A(\core.keymem.key_mem[11][23] ),
    .B(_13196_),
    .S(_13938_),
    .Z(_01136_));
 NAND2_X1 _36843_ (.A1(\core.keymem.key_mem[11][24] ),
    .A2(_13941_),
    .ZN(_13944_));
 OAI21_X1 _36844_ (.A(_13944_),
    .B1(_13930_),
    .B2(_13212_),
    .ZN(_01137_));
 MUX2_X1 _36845_ (.A(\core.keymem.key_mem[11][25] ),
    .B(_13233_),
    .S(_13938_),
    .Z(_01138_));
 MUX2_X1 _36846_ (.A(\core.keymem.key_mem[11][26] ),
    .B(_13241_),
    .S(_13938_),
    .Z(_01139_));
 BUF_X4 _36847_ (.A(_13922_),
    .Z(_13945_));
 MUX2_X1 _36848_ (.A(\core.keymem.key_mem[11][27] ),
    .B(_13284_),
    .S(_13945_),
    .Z(_01140_));
 MUX2_X1 _36849_ (.A(\core.keymem.key_mem[11][28] ),
    .B(_13325_),
    .S(_13945_),
    .Z(_01141_));
 MUX2_X1 _36850_ (.A(\core.keymem.key_mem[11][29] ),
    .B(_13329_),
    .S(_13945_),
    .Z(_01142_));
 NAND2_X1 _36851_ (.A1(\core.keymem.key_mem[11][2] ),
    .A2(_13941_),
    .ZN(_13946_));
 OAI21_X1 _36852_ (.A(_13946_),
    .B1(_13930_),
    .B2(_13335_),
    .ZN(_01143_));
 MUX2_X1 _36853_ (.A(\core.keymem.key_mem[11][30] ),
    .B(_13379_),
    .S(_13945_),
    .Z(_01144_));
 MUX2_X1 _36854_ (.A(\core.keymem.key_mem[11][31] ),
    .B(_13395_),
    .S(_13945_),
    .Z(_01145_));
 MUX2_X1 _36855_ (.A(\core.keymem.key_mem[11][32] ),
    .B(_13396_),
    .S(_13945_),
    .Z(_01146_));
 MUX2_X1 _36856_ (.A(\core.keymem.key_mem[11][33] ),
    .B(_13402_),
    .S(_13945_),
    .Z(_01147_));
 MUX2_X1 _36857_ (.A(\core.keymem.key_mem[11][34] ),
    .B(_13403_),
    .S(_13945_),
    .Z(_01148_));
 MUX2_X1 _36858_ (.A(\core.keymem.key_mem[11][35] ),
    .B(_13405_),
    .S(_13945_),
    .Z(_01149_));
 NAND2_X1 _36859_ (.A1(\core.keymem.key_mem[11][36] ),
    .A2(_13941_),
    .ZN(_13947_));
 BUF_X4 _36860_ (.A(_13929_),
    .Z(_13948_));
 OAI21_X1 _36861_ (.A(_13947_),
    .B1(_13948_),
    .B2(_13407_),
    .ZN(_01150_));
 NAND2_X1 _36862_ (.A1(\core.keymem.key_mem[11][37] ),
    .A2(_13941_),
    .ZN(_13949_));
 OAI21_X1 _36863_ (.A(_13949_),
    .B1(_13948_),
    .B2(_12439_),
    .ZN(_01151_));
 MUX2_X1 _36864_ (.A(\core.keymem.key_mem[11][38] ),
    .B(_13410_),
    .S(_13945_),
    .Z(_01152_));
 NAND2_X1 _36865_ (.A1(\core.keymem.key_mem[11][39] ),
    .A2(_13941_),
    .ZN(_13950_));
 OAI21_X1 _36866_ (.A(_13950_),
    .B1(_13948_),
    .B2(_13435_),
    .ZN(_01153_));
 NAND2_X1 _36867_ (.A1(\core.keymem.key_mem[11][3] ),
    .A2(_13941_),
    .ZN(_13951_));
 OAI21_X1 _36868_ (.A(_13951_),
    .B1(_13948_),
    .B2(_13448_),
    .ZN(_01154_));
 NAND2_X1 _36869_ (.A1(\core.keymem.key_mem[11][40] ),
    .A2(_13941_),
    .ZN(_13952_));
 OAI21_X1 _36870_ (.A(_13952_),
    .B1(_13948_),
    .B2(_13457_),
    .ZN(_01155_));
 BUF_X4 _36871_ (.A(_13922_),
    .Z(_13953_));
 MUX2_X1 _36872_ (.A(\core.keymem.key_mem[11][41] ),
    .B(_13467_),
    .S(_13953_),
    .Z(_01156_));
 MUX2_X1 _36873_ (.A(\core.keymem.key_mem[11][42] ),
    .B(_13490_),
    .S(_13953_),
    .Z(_01157_));
 NAND2_X1 _36874_ (.A1(\core.keymem.key_mem[11][43] ),
    .A2(_13941_),
    .ZN(_13954_));
 OAI21_X1 _36875_ (.A(_13954_),
    .B1(_13948_),
    .B2(_13496_),
    .ZN(_01158_));
 MUX2_X1 _36876_ (.A(\core.keymem.key_mem[11][44] ),
    .B(_13497_),
    .S(_13953_),
    .Z(_01159_));
 NAND2_X1 _36877_ (.A1(\core.keymem.key_mem[11][45] ),
    .A2(_13941_),
    .ZN(_13955_));
 OAI21_X1 _36878_ (.A(_13955_),
    .B1(_13948_),
    .B2(_13510_),
    .ZN(_01160_));
 BUF_X4 _36879_ (.A(_13926_),
    .Z(_13956_));
 NAND2_X1 _36880_ (.A1(\core.keymem.key_mem[11][46] ),
    .A2(_13956_),
    .ZN(_13957_));
 OAI21_X1 _36881_ (.A(_13957_),
    .B1(_13948_),
    .B2(_13517_),
    .ZN(_01161_));
 NAND2_X1 _36882_ (.A1(\core.keymem.key_mem[11][47] ),
    .A2(_13956_),
    .ZN(_13958_));
 OAI21_X1 _36883_ (.A(_13958_),
    .B1(_13948_),
    .B2(_12520_),
    .ZN(_01162_));
 NAND2_X1 _36884_ (.A1(\core.keymem.key_mem[11][48] ),
    .A2(_13956_),
    .ZN(_13959_));
 OAI21_X1 _36885_ (.A(_13959_),
    .B1(_13948_),
    .B2(_12532_),
    .ZN(_01163_));
 NAND2_X1 _36886_ (.A1(\core.keymem.key_mem[11][49] ),
    .A2(_13956_),
    .ZN(_13960_));
 BUF_X4 _36887_ (.A(_13929_),
    .Z(_13961_));
 OAI21_X1 _36888_ (.A(_13960_),
    .B1(_13961_),
    .B2(_13529_),
    .ZN(_01164_));
 MUX2_X1 _36889_ (.A(\core.keymem.key_mem[11][4] ),
    .B(_13538_),
    .S(_13953_),
    .Z(_01165_));
 MUX2_X1 _36890_ (.A(\core.keymem.key_mem[11][50] ),
    .B(_13557_),
    .S(_13953_),
    .Z(_01166_));
 MUX2_X1 _36891_ (.A(\core.keymem.key_mem[11][51] ),
    .B(_13564_),
    .S(_13953_),
    .Z(_01167_));
 NAND2_X1 _36892_ (.A1(\core.keymem.key_mem[11][52] ),
    .A2(_13956_),
    .ZN(_13962_));
 OAI21_X1 _36893_ (.A(_13962_),
    .B1(_13961_),
    .B2(_12568_),
    .ZN(_01168_));
 NAND2_X1 _36894_ (.A1(\core.keymem.key_mem[11][53] ),
    .A2(_13956_),
    .ZN(_13963_));
 OAI21_X1 _36895_ (.A(_13963_),
    .B1(_13961_),
    .B2(_12584_),
    .ZN(_01169_));
 NAND2_X1 _36896_ (.A1(\core.keymem.key_mem[11][54] ),
    .A2(_13956_),
    .ZN(_13964_));
 OAI21_X1 _36897_ (.A(_13964_),
    .B1(_13961_),
    .B2(_13575_),
    .ZN(_01170_));
 MUX2_X1 _36898_ (.A(\core.keymem.key_mem[11][55] ),
    .B(_13581_),
    .S(_13953_),
    .Z(_01171_));
 MUX2_X1 _36899_ (.A(\core.keymem.key_mem[11][56] ),
    .B(_13589_),
    .S(_13953_),
    .Z(_01172_));
 MUX2_X1 _36900_ (.A(\core.keymem.key_mem[11][57] ),
    .B(_13604_),
    .S(_13953_),
    .Z(_01173_));
 MUX2_X1 _36901_ (.A(\core.keymem.key_mem[11][58] ),
    .B(_13611_),
    .S(_13953_),
    .Z(_01174_));
 BUF_X4 _36902_ (.A(_13922_),
    .Z(_13965_));
 MUX2_X1 _36903_ (.A(\core.keymem.key_mem[11][59] ),
    .B(_13616_),
    .S(_13965_),
    .Z(_01175_));
 MUX2_X1 _36904_ (.A(\core.keymem.key_mem[11][5] ),
    .B(_12606_),
    .S(_13965_),
    .Z(_01176_));
 MUX2_X1 _36905_ (.A(\core.keymem.key_mem[11][60] ),
    .B(_13622_),
    .S(_13965_),
    .Z(_01177_));
 MUX2_X1 _36906_ (.A(\core.keymem.key_mem[11][61] ),
    .B(_13632_),
    .S(_13965_),
    .Z(_01178_));
 MUX2_X1 _36907_ (.A(\core.keymem.key_mem[11][62] ),
    .B(_13637_),
    .S(_13965_),
    .Z(_01179_));
 MUX2_X1 _36908_ (.A(\core.keymem.key_mem[11][63] ),
    .B(_13659_),
    .S(_13965_),
    .Z(_01180_));
 MUX2_X1 _36909_ (.A(\core.keymem.key_mem[11][64] ),
    .B(_12622_),
    .S(_13965_),
    .Z(_01181_));
 NAND2_X1 _36910_ (.A1(\core.keymem.key_mem[11][65] ),
    .A2(_13956_),
    .ZN(_13966_));
 OAI21_X1 _36911_ (.A(_13966_),
    .B1(_13961_),
    .B2(_13673_),
    .ZN(_01182_));
 MUX2_X1 _36912_ (.A(\core.keymem.key_mem[11][66] ),
    .B(_13681_),
    .S(_13965_),
    .Z(_01183_));
 NAND2_X1 _36913_ (.A1(\core.keymem.key_mem[11][67] ),
    .A2(_13956_),
    .ZN(_13967_));
 OAI21_X1 _36914_ (.A(_13967_),
    .B1(_13961_),
    .B2(_13690_),
    .ZN(_01184_));
 NAND2_X1 _36915_ (.A1(\core.keymem.key_mem[11][68] ),
    .A2(_13956_),
    .ZN(_13968_));
 OAI21_X1 _36916_ (.A(_13968_),
    .B1(_13961_),
    .B2(_12635_),
    .ZN(_01185_));
 BUF_X4 _36917_ (.A(_13926_),
    .Z(_13969_));
 NAND2_X1 _36918_ (.A1(\core.keymem.key_mem[11][69] ),
    .A2(_13969_),
    .ZN(_13970_));
 OAI21_X1 _36919_ (.A(_13970_),
    .B1(_13961_),
    .B2(_13700_),
    .ZN(_01186_));
 MUX2_X1 _36920_ (.A(\core.keymem.key_mem[11][6] ),
    .B(_13711_),
    .S(_13965_),
    .Z(_01187_));
 MUX2_X1 _36921_ (.A(\core.keymem.key_mem[11][70] ),
    .B(_13713_),
    .S(_13965_),
    .Z(_01188_));
 NAND2_X1 _36922_ (.A1(\core.keymem.key_mem[11][71] ),
    .A2(_13969_),
    .ZN(_13971_));
 OAI21_X1 _36923_ (.A(_13971_),
    .B1(_13961_),
    .B2(_12659_),
    .ZN(_01189_));
 NAND2_X1 _36924_ (.A1(\core.keymem.key_mem[11][72] ),
    .A2(_13969_),
    .ZN(_13972_));
 OAI21_X1 _36925_ (.A(_13972_),
    .B1(_13961_),
    .B2(_13716_),
    .ZN(_01190_));
 NAND2_X1 _36926_ (.A1(\core.keymem.key_mem[11][73] ),
    .A2(_13969_),
    .ZN(_13973_));
 BUF_X4 _36927_ (.A(_13929_),
    .Z(_13974_));
 OAI21_X1 _36928_ (.A(_13973_),
    .B1(_13974_),
    .B2(_12688_),
    .ZN(_01191_));
 NAND2_X1 _36929_ (.A1(\core.keymem.key_mem[11][74] ),
    .A2(_13969_),
    .ZN(_13975_));
 OAI21_X1 _36930_ (.A(_13975_),
    .B1(_13974_),
    .B2(_13726_),
    .ZN(_01192_));
 NAND2_X1 _36931_ (.A1(\core.keymem.key_mem[11][75] ),
    .A2(_13969_),
    .ZN(_13976_));
 OAI21_X1 _36932_ (.A(_13976_),
    .B1(_13974_),
    .B2(_13733_),
    .ZN(_01193_));
 BUF_X4 _36933_ (.A(_13922_),
    .Z(_13977_));
 MUX2_X1 _36934_ (.A(\core.keymem.key_mem[11][76] ),
    .B(_13741_),
    .S(_13977_),
    .Z(_01194_));
 MUX2_X1 _36935_ (.A(\core.keymem.key_mem[11][77] ),
    .B(_13751_),
    .S(_13977_),
    .Z(_01195_));
 NAND2_X1 _36936_ (.A1(\core.keymem.key_mem[11][78] ),
    .A2(_13969_),
    .ZN(_13978_));
 OAI21_X1 _36937_ (.A(_13978_),
    .B1(_13974_),
    .B2(_12708_),
    .ZN(_01196_));
 MUX2_X1 _36938_ (.A(\core.keymem.key_mem[11][79] ),
    .B(_13758_),
    .S(_13977_),
    .Z(_01197_));
 NAND2_X1 _36939_ (.A1(\core.keymem.key_mem[11][7] ),
    .A2(_13969_),
    .ZN(_13979_));
 OAI21_X1 _36940_ (.A(_13979_),
    .B1(_13974_),
    .B2(_13767_),
    .ZN(_01198_));
 MUX2_X1 _36941_ (.A(\core.keymem.key_mem[11][80] ),
    .B(_13769_),
    .S(_13977_),
    .Z(_01199_));
 NAND2_X1 _36942_ (.A1(\core.keymem.key_mem[11][81] ),
    .A2(_13969_),
    .ZN(_13980_));
 OAI21_X1 _36943_ (.A(_13980_),
    .B1(_13974_),
    .B2(_13775_),
    .ZN(_01200_));
 NAND2_X1 _36944_ (.A1(\core.keymem.key_mem[11][82] ),
    .A2(_13969_),
    .ZN(_13981_));
 OAI21_X1 _36945_ (.A(_13981_),
    .B1(_13974_),
    .B2(_13783_),
    .ZN(_01201_));
 NAND2_X1 _36946_ (.A1(\core.keymem.key_mem[11][83] ),
    .A2(_13929_),
    .ZN(_13982_));
 OAI21_X1 _36947_ (.A(_13982_),
    .B1(_13974_),
    .B2(_13791_),
    .ZN(_01202_));
 NAND2_X1 _36948_ (.A1(\core.keymem.key_mem[11][84] ),
    .A2(_13929_),
    .ZN(_13983_));
 OAI21_X1 _36949_ (.A(_13983_),
    .B1(_13974_),
    .B2(_12725_),
    .ZN(_01203_));
 MUX2_X1 _36950_ (.A(\core.keymem.key_mem[11][85] ),
    .B(_13798_),
    .S(_13977_),
    .Z(_01204_));
 MUX2_X1 _36951_ (.A(\core.keymem.key_mem[11][86] ),
    .B(_12741_),
    .S(_13977_),
    .Z(_01205_));
 MUX2_X1 _36952_ (.A(\core.keymem.key_mem[11][87] ),
    .B(_13804_),
    .S(_13977_),
    .Z(_01206_));
 MUX2_X1 _36953_ (.A(\core.keymem.key_mem[11][88] ),
    .B(_13810_),
    .S(_13977_),
    .Z(_01207_));
 MUX2_X1 _36954_ (.A(\core.keymem.key_mem[11][89] ),
    .B(_13818_),
    .S(_13977_),
    .Z(_01208_));
 MUX2_X1 _36955_ (.A(\core.keymem.key_mem[11][8] ),
    .B(_13854_),
    .S(_13977_),
    .Z(_01209_));
 MUX2_X1 _36956_ (.A(\core.keymem.key_mem[11][90] ),
    .B(_13860_),
    .S(_13923_),
    .Z(_01210_));
 NAND2_X1 _36957_ (.A1(\core.keymem.key_mem[11][91] ),
    .A2(_13929_),
    .ZN(_13984_));
 OAI21_X1 _36958_ (.A(_13984_),
    .B1(_13974_),
    .B2(_13870_),
    .ZN(_01211_));
 NAND2_X1 _36959_ (.A1(\core.keymem.key_mem[11][92] ),
    .A2(_13929_),
    .ZN(_13985_));
 OAI21_X1 _36960_ (.A(_13985_),
    .B1(_13927_),
    .B2(_13880_),
    .ZN(_01212_));
 MUX2_X1 _36961_ (.A(\core.keymem.key_mem[11][93] ),
    .B(_13889_),
    .S(_13923_),
    .Z(_01213_));
 MUX2_X1 _36962_ (.A(\core.keymem.key_mem[11][94] ),
    .B(_13896_),
    .S(_13923_),
    .Z(_01214_));
 MUX2_X1 _36963_ (.A(\core.keymem.key_mem[11][95] ),
    .B(_13903_),
    .S(_13923_),
    .Z(_01215_));
 MUX2_X1 _36964_ (.A(\core.keymem.key_mem[11][96] ),
    .B(_13907_),
    .S(_13923_),
    .Z(_01216_));
 NAND2_X1 _36965_ (.A1(\core.keymem.key_mem[11][97] ),
    .A2(_13929_),
    .ZN(_13986_));
 OAI21_X1 _36966_ (.A(_13986_),
    .B1(_13927_),
    .B2(_12777_),
    .ZN(_01217_));
 NAND2_X1 _36967_ (.A1(\core.keymem.key_mem[11][98] ),
    .A2(_13929_),
    .ZN(_13987_));
 OAI21_X1 _36968_ (.A(_13987_),
    .B1(_13927_),
    .B2(_13910_),
    .ZN(_01218_));
 MUX2_X1 _36969_ (.A(\core.keymem.key_mem[11][99] ),
    .B(_12800_),
    .S(_13923_),
    .Z(_01219_));
 MUX2_X1 _36970_ (.A(\core.keymem.key_mem[11][9] ),
    .B(_13919_),
    .S(_13923_),
    .Z(_01220_));
 NAND2_X4 _36971_ (.A1(_11794_),
    .A2(_16218_),
    .ZN(_13988_));
 NAND2_X4 _36972_ (.A1(_16222_),
    .A2(_11793_),
    .ZN(_13989_));
 NOR2_X4 _36973_ (.A1(_13988_),
    .A2(_13989_),
    .ZN(_13990_));
 BUF_X4 _36974_ (.A(_13990_),
    .Z(_13991_));
 BUF_X4 _36975_ (.A(_13991_),
    .Z(_13992_));
 MUX2_X1 _36976_ (.A(\core.keymem.key_mem[12][0] ),
    .B(_11844_),
    .S(_13992_),
    .Z(_01221_));
 MUX2_X1 _36977_ (.A(\core.keymem.key_mem[12][100] ),
    .B(_11873_),
    .S(_13992_),
    .Z(_01222_));
 MUX2_X1 _36978_ (.A(\core.keymem.key_mem[12][101] ),
    .B(_12813_),
    .S(_13992_),
    .Z(_01223_));
 MUX2_X1 _36979_ (.A(\core.keymem.key_mem[12][102] ),
    .B(_11906_),
    .S(_13992_),
    .Z(_01224_));
 MUX2_X1 _36980_ (.A(\core.keymem.key_mem[12][103] ),
    .B(_11929_),
    .S(_13992_),
    .Z(_01225_));
 OR2_X1 _36981_ (.A1(_13988_),
    .A2(_13989_),
    .ZN(_13993_));
 CLKBUF_X3 _36982_ (.A(_13993_),
    .Z(_13994_));
 BUF_X4 _36983_ (.A(_13994_),
    .Z(_13995_));
 NAND2_X1 _36984_ (.A1(\core.keymem.key_mem[12][104] ),
    .A2(_13995_),
    .ZN(_13996_));
 BUF_X4 _36985_ (.A(_13994_),
    .Z(_13997_));
 BUF_X4 _36986_ (.A(_13997_),
    .Z(_13998_));
 OAI21_X1 _36987_ (.A(_13996_),
    .B1(_13998_),
    .B2(_12822_),
    .ZN(_01226_));
 MUX2_X1 _36988_ (.A(\core.keymem.key_mem[12][105] ),
    .B(_12830_),
    .S(_13992_),
    .Z(_01227_));
 BUF_X4 _36989_ (.A(_13991_),
    .Z(_13999_));
 MUX2_X1 _36990_ (.A(\core.keymem.key_mem[12][106] ),
    .B(_12832_),
    .S(_13999_),
    .Z(_01228_));
 MUX2_X1 _36991_ (.A(\core.keymem.key_mem[12][107] ),
    .B(_11967_),
    .S(_13999_),
    .Z(_01229_));
 MUX2_X1 _36992_ (.A(\core.keymem.key_mem[12][108] ),
    .B(_11981_),
    .S(_13999_),
    .Z(_01230_));
 MUX2_X1 _36993_ (.A(\core.keymem.key_mem[12][109] ),
    .B(_12842_),
    .S(_13999_),
    .Z(_01231_));
 NAND2_X1 _36994_ (.A1(\core.keymem.key_mem[12][10] ),
    .A2(_13995_),
    .ZN(_14000_));
 OAI21_X1 _36995_ (.A(_14000_),
    .B1(_13998_),
    .B2(_12858_),
    .ZN(_01232_));
 MUX2_X1 _36996_ (.A(\core.keymem.key_mem[12][110] ),
    .B(_12859_),
    .S(_13999_),
    .Z(_01233_));
 MUX2_X1 _36997_ (.A(\core.keymem.key_mem[12][111] ),
    .B(_12017_),
    .S(_13999_),
    .Z(_01234_));
 MUX2_X1 _36998_ (.A(\core.keymem.key_mem[12][112] ),
    .B(_12031_),
    .S(_13999_),
    .Z(_01235_));
 MUX2_X1 _36999_ (.A(\core.keymem.key_mem[12][113] ),
    .B(_12868_),
    .S(_13999_),
    .Z(_01236_));
 MUX2_X1 _37000_ (.A(\core.keymem.key_mem[12][114] ),
    .B(_12869_),
    .S(_13999_),
    .Z(_01237_));
 MUX2_X1 _37001_ (.A(\core.keymem.key_mem[12][115] ),
    .B(_12059_),
    .S(_13999_),
    .Z(_01238_));
 BUF_X4 _37002_ (.A(_13991_),
    .Z(_14001_));
 MUX2_X1 _37003_ (.A(\core.keymem.key_mem[12][116] ),
    .B(_12077_),
    .S(_14001_),
    .Z(_01239_));
 MUX2_X1 _37004_ (.A(\core.keymem.key_mem[12][117] ),
    .B(_12877_),
    .S(_14001_),
    .Z(_01240_));
 MUX2_X1 _37005_ (.A(\core.keymem.key_mem[12][118] ),
    .B(_12882_),
    .S(_14001_),
    .Z(_01241_));
 MUX2_X1 _37006_ (.A(\core.keymem.key_mem[12][119] ),
    .B(_12096_),
    .S(_14001_),
    .Z(_01242_));
 NAND2_X1 _37007_ (.A1(\core.keymem.key_mem[12][11] ),
    .A2(_13995_),
    .ZN(_14002_));
 OAI21_X1 _37008_ (.A(_14002_),
    .B1(_13998_),
    .B2(_12895_),
    .ZN(_01243_));
 MUX2_X1 _37009_ (.A(\core.keymem.key_mem[12][120] ),
    .B(_12124_),
    .S(_14001_),
    .Z(_01244_));
 MUX2_X1 _37010_ (.A(\core.keymem.key_mem[12][121] ),
    .B(_12160_),
    .S(_14001_),
    .Z(_01245_));
 MUX2_X1 _37011_ (.A(\core.keymem.key_mem[12][122] ),
    .B(_12903_),
    .S(_14001_),
    .Z(_01246_));
 NAND2_X1 _37012_ (.A1(\core.keymem.key_mem[12][123] ),
    .A2(_13995_),
    .ZN(_14003_));
 OAI21_X1 _37013_ (.A(_14003_),
    .B1(_13998_),
    .B2(_12182_),
    .ZN(_01247_));
 NAND2_X1 _37014_ (.A1(\core.keymem.key_mem[12][124] ),
    .A2(_13995_),
    .ZN(_14004_));
 OAI21_X1 _37015_ (.A(_14004_),
    .B1(_13998_),
    .B2(_12926_),
    .ZN(_01248_));
 MUX2_X1 _37016_ (.A(\core.keymem.key_mem[12][125] ),
    .B(_12932_),
    .S(_14001_),
    .Z(_01249_));
 NAND2_X1 _37017_ (.A1(\core.keymem.key_mem[12][126] ),
    .A2(_13995_),
    .ZN(_14005_));
 OAI21_X1 _37018_ (.A(_14005_),
    .B1(_13998_),
    .B2(_12207_),
    .ZN(_01250_));
 MUX2_X1 _37019_ (.A(\core.keymem.key_mem[12][127] ),
    .B(_12945_),
    .S(_14001_),
    .Z(_01251_));
 MUX2_X1 _37020_ (.A(\core.keymem.key_mem[12][12] ),
    .B(_12958_),
    .S(_14001_),
    .Z(_01252_));
 BUF_X4 _37021_ (.A(_13990_),
    .Z(_14006_));
 MUX2_X1 _37022_ (.A(\core.keymem.key_mem[12][13] ),
    .B(_12974_),
    .S(_14006_),
    .Z(_01253_));
 NOR2_X1 _37023_ (.A1(\core.keymem.key_mem[12][14] ),
    .A2(_13992_),
    .ZN(_14007_));
 AOI21_X1 _37024_ (.A(_14007_),
    .B1(_13992_),
    .B2(_13007_),
    .ZN(_01254_));
 MUX2_X1 _37025_ (.A(\core.keymem.key_mem[12][15] ),
    .B(_13017_),
    .S(_14006_),
    .Z(_01255_));
 MUX2_X1 _37026_ (.A(\core.keymem.key_mem[12][16] ),
    .B(_13029_),
    .S(_14006_),
    .Z(_01256_));
 NAND2_X1 _37027_ (.A1(\core.keymem.key_mem[12][17] ),
    .A2(_13995_),
    .ZN(_14008_));
 OAI21_X1 _37028_ (.A(_14008_),
    .B1(_13998_),
    .B2(_13042_),
    .ZN(_01257_));
 MUX2_X1 _37029_ (.A(\core.keymem.key_mem[12][18] ),
    .B(_13094_),
    .S(_14006_),
    .Z(_01258_));
 BUF_X4 _37030_ (.A(_13994_),
    .Z(_14009_));
 NAND2_X1 _37031_ (.A1(\core.keymem.key_mem[12][19] ),
    .A2(_14009_),
    .ZN(_14010_));
 OAI21_X1 _37032_ (.A(_14010_),
    .B1(_13998_),
    .B2(_13109_),
    .ZN(_01259_));
 MUX2_X1 _37033_ (.A(\core.keymem.key_mem[12][1] ),
    .B(_13134_),
    .S(_14006_),
    .Z(_01260_));
 MUX2_X1 _37034_ (.A(\core.keymem.key_mem[12][20] ),
    .B(_13146_),
    .S(_14006_),
    .Z(_01261_));
 MUX2_X1 _37035_ (.A(\core.keymem.key_mem[12][21] ),
    .B(_13155_),
    .S(_14006_),
    .Z(_01262_));
 NOR2_X1 _37036_ (.A1(\core.keymem.key_mem[12][22] ),
    .A2(_13992_),
    .ZN(_14011_));
 AOI21_X1 _37037_ (.A(_14011_),
    .B1(_13992_),
    .B2(_13191_),
    .ZN(_01263_));
 MUX2_X1 _37038_ (.A(\core.keymem.key_mem[12][23] ),
    .B(_13196_),
    .S(_14006_),
    .Z(_01264_));
 NAND2_X1 _37039_ (.A1(\core.keymem.key_mem[12][24] ),
    .A2(_14009_),
    .ZN(_14012_));
 OAI21_X1 _37040_ (.A(_14012_),
    .B1(_13998_),
    .B2(_13212_),
    .ZN(_01265_));
 MUX2_X1 _37041_ (.A(\core.keymem.key_mem[12][25] ),
    .B(_13233_),
    .S(_14006_),
    .Z(_01266_));
 MUX2_X1 _37042_ (.A(\core.keymem.key_mem[12][26] ),
    .B(_13241_),
    .S(_14006_),
    .Z(_01267_));
 BUF_X4 _37043_ (.A(_13990_),
    .Z(_14013_));
 MUX2_X1 _37044_ (.A(\core.keymem.key_mem[12][27] ),
    .B(_13284_),
    .S(_14013_),
    .Z(_01268_));
 MUX2_X1 _37045_ (.A(\core.keymem.key_mem[12][28] ),
    .B(_13325_),
    .S(_14013_),
    .Z(_01269_));
 MUX2_X1 _37046_ (.A(\core.keymem.key_mem[12][29] ),
    .B(_13329_),
    .S(_14013_),
    .Z(_01270_));
 NAND2_X1 _37047_ (.A1(\core.keymem.key_mem[12][2] ),
    .A2(_14009_),
    .ZN(_14014_));
 OAI21_X1 _37048_ (.A(_14014_),
    .B1(_13998_),
    .B2(_13335_),
    .ZN(_01271_));
 MUX2_X1 _37049_ (.A(\core.keymem.key_mem[12][30] ),
    .B(_13379_),
    .S(_14013_),
    .Z(_01272_));
 MUX2_X1 _37050_ (.A(\core.keymem.key_mem[12][31] ),
    .B(_13395_),
    .S(_14013_),
    .Z(_01273_));
 MUX2_X1 _37051_ (.A(\core.keymem.key_mem[12][32] ),
    .B(_13396_),
    .S(_14013_),
    .Z(_01274_));
 MUX2_X1 _37052_ (.A(\core.keymem.key_mem[12][33] ),
    .B(_13402_),
    .S(_14013_),
    .Z(_01275_));
 MUX2_X1 _37053_ (.A(\core.keymem.key_mem[12][34] ),
    .B(_13403_),
    .S(_14013_),
    .Z(_01276_));
 MUX2_X1 _37054_ (.A(\core.keymem.key_mem[12][35] ),
    .B(_13405_),
    .S(_14013_),
    .Z(_01277_));
 NAND2_X1 _37055_ (.A1(\core.keymem.key_mem[12][36] ),
    .A2(_14009_),
    .ZN(_14015_));
 BUF_X4 _37056_ (.A(_13997_),
    .Z(_14016_));
 OAI21_X1 _37057_ (.A(_14015_),
    .B1(_14016_),
    .B2(_13407_),
    .ZN(_01278_));
 NAND2_X1 _37058_ (.A1(\core.keymem.key_mem[12][37] ),
    .A2(_14009_),
    .ZN(_14017_));
 OAI21_X1 _37059_ (.A(_14017_),
    .B1(_14016_),
    .B2(_12439_),
    .ZN(_01279_));
 MUX2_X1 _37060_ (.A(\core.keymem.key_mem[12][38] ),
    .B(_13410_),
    .S(_14013_),
    .Z(_01280_));
 NAND2_X1 _37061_ (.A1(\core.keymem.key_mem[12][39] ),
    .A2(_14009_),
    .ZN(_14018_));
 OAI21_X1 _37062_ (.A(_14018_),
    .B1(_14016_),
    .B2(_13435_),
    .ZN(_01281_));
 NAND2_X1 _37063_ (.A1(\core.keymem.key_mem[12][3] ),
    .A2(_14009_),
    .ZN(_14019_));
 OAI21_X1 _37064_ (.A(_14019_),
    .B1(_14016_),
    .B2(_13448_),
    .ZN(_01282_));
 NAND2_X1 _37065_ (.A1(\core.keymem.key_mem[12][40] ),
    .A2(_14009_),
    .ZN(_14020_));
 OAI21_X1 _37066_ (.A(_14020_),
    .B1(_14016_),
    .B2(_13457_),
    .ZN(_01283_));
 BUF_X4 _37067_ (.A(_13990_),
    .Z(_14021_));
 MUX2_X1 _37068_ (.A(\core.keymem.key_mem[12][41] ),
    .B(_13467_),
    .S(_14021_),
    .Z(_01284_));
 MUX2_X1 _37069_ (.A(\core.keymem.key_mem[12][42] ),
    .B(_13490_),
    .S(_14021_),
    .Z(_01285_));
 NAND2_X1 _37070_ (.A1(\core.keymem.key_mem[12][43] ),
    .A2(_14009_),
    .ZN(_14022_));
 OAI21_X1 _37071_ (.A(_14022_),
    .B1(_14016_),
    .B2(_13496_),
    .ZN(_01286_));
 MUX2_X1 _37072_ (.A(\core.keymem.key_mem[12][44] ),
    .B(_13497_),
    .S(_14021_),
    .Z(_01287_));
 NAND2_X1 _37073_ (.A1(\core.keymem.key_mem[12][45] ),
    .A2(_14009_),
    .ZN(_14023_));
 OAI21_X1 _37074_ (.A(_14023_),
    .B1(_14016_),
    .B2(_13510_),
    .ZN(_01288_));
 BUF_X4 _37075_ (.A(_13994_),
    .Z(_14024_));
 NAND2_X1 _37076_ (.A1(\core.keymem.key_mem[12][46] ),
    .A2(_14024_),
    .ZN(_14025_));
 OAI21_X1 _37077_ (.A(_14025_),
    .B1(_14016_),
    .B2(_13517_),
    .ZN(_01289_));
 NAND2_X1 _37078_ (.A1(\core.keymem.key_mem[12][47] ),
    .A2(_14024_),
    .ZN(_14026_));
 OAI21_X1 _37079_ (.A(_14026_),
    .B1(_14016_),
    .B2(_12520_),
    .ZN(_01290_));
 NAND2_X1 _37080_ (.A1(\core.keymem.key_mem[12][48] ),
    .A2(_14024_),
    .ZN(_14027_));
 OAI21_X1 _37081_ (.A(_14027_),
    .B1(_14016_),
    .B2(_12532_),
    .ZN(_01291_));
 NAND2_X1 _37082_ (.A1(\core.keymem.key_mem[12][49] ),
    .A2(_14024_),
    .ZN(_14028_));
 BUF_X4 _37083_ (.A(_13997_),
    .Z(_14029_));
 OAI21_X1 _37084_ (.A(_14028_),
    .B1(_14029_),
    .B2(_13529_),
    .ZN(_01292_));
 MUX2_X1 _37085_ (.A(\core.keymem.key_mem[12][4] ),
    .B(_13538_),
    .S(_14021_),
    .Z(_01293_));
 MUX2_X1 _37086_ (.A(\core.keymem.key_mem[12][50] ),
    .B(_13557_),
    .S(_14021_),
    .Z(_01294_));
 MUX2_X1 _37087_ (.A(\core.keymem.key_mem[12][51] ),
    .B(_13564_),
    .S(_14021_),
    .Z(_01295_));
 NAND2_X1 _37088_ (.A1(\core.keymem.key_mem[12][52] ),
    .A2(_14024_),
    .ZN(_14030_));
 OAI21_X1 _37089_ (.A(_14030_),
    .B1(_14029_),
    .B2(_12568_),
    .ZN(_01296_));
 NAND2_X1 _37090_ (.A1(\core.keymem.key_mem[12][53] ),
    .A2(_14024_),
    .ZN(_14031_));
 OAI21_X1 _37091_ (.A(_14031_),
    .B1(_14029_),
    .B2(_12584_),
    .ZN(_01297_));
 NAND2_X1 _37092_ (.A1(\core.keymem.key_mem[12][54] ),
    .A2(_14024_),
    .ZN(_14032_));
 OAI21_X1 _37093_ (.A(_14032_),
    .B1(_14029_),
    .B2(_13575_),
    .ZN(_01298_));
 MUX2_X1 _37094_ (.A(\core.keymem.key_mem[12][55] ),
    .B(_13581_),
    .S(_14021_),
    .Z(_01299_));
 MUX2_X1 _37095_ (.A(\core.keymem.key_mem[12][56] ),
    .B(_13589_),
    .S(_14021_),
    .Z(_01300_));
 MUX2_X1 _37096_ (.A(\core.keymem.key_mem[12][57] ),
    .B(_13604_),
    .S(_14021_),
    .Z(_01301_));
 MUX2_X1 _37097_ (.A(\core.keymem.key_mem[12][58] ),
    .B(_13611_),
    .S(_14021_),
    .Z(_01302_));
 BUF_X4 _37098_ (.A(_13990_),
    .Z(_14033_));
 MUX2_X1 _37099_ (.A(\core.keymem.key_mem[12][59] ),
    .B(_13616_),
    .S(_14033_),
    .Z(_01303_));
 MUX2_X1 _37100_ (.A(\core.keymem.key_mem[12][5] ),
    .B(_12606_),
    .S(_14033_),
    .Z(_01304_));
 MUX2_X1 _37101_ (.A(\core.keymem.key_mem[12][60] ),
    .B(_13622_),
    .S(_14033_),
    .Z(_01305_));
 MUX2_X1 _37102_ (.A(\core.keymem.key_mem[12][61] ),
    .B(_13632_),
    .S(_14033_),
    .Z(_01306_));
 MUX2_X1 _37103_ (.A(\core.keymem.key_mem[12][62] ),
    .B(_13637_),
    .S(_14033_),
    .Z(_01307_));
 MUX2_X1 _37104_ (.A(\core.keymem.key_mem[12][63] ),
    .B(_13659_),
    .S(_14033_),
    .Z(_01308_));
 MUX2_X1 _37105_ (.A(\core.keymem.key_mem[12][64] ),
    .B(_12622_),
    .S(_14033_),
    .Z(_01309_));
 NAND2_X1 _37106_ (.A1(\core.keymem.key_mem[12][65] ),
    .A2(_14024_),
    .ZN(_14034_));
 OAI21_X1 _37107_ (.A(_14034_),
    .B1(_14029_),
    .B2(_13673_),
    .ZN(_01310_));
 MUX2_X1 _37108_ (.A(\core.keymem.key_mem[12][66] ),
    .B(_13681_),
    .S(_14033_),
    .Z(_01311_));
 NAND2_X1 _37109_ (.A1(\core.keymem.key_mem[12][67] ),
    .A2(_14024_),
    .ZN(_14035_));
 OAI21_X1 _37110_ (.A(_14035_),
    .B1(_14029_),
    .B2(_13690_),
    .ZN(_01312_));
 NAND2_X1 _37111_ (.A1(\core.keymem.key_mem[12][68] ),
    .A2(_14024_),
    .ZN(_14036_));
 OAI21_X1 _37112_ (.A(_14036_),
    .B1(_14029_),
    .B2(_12635_),
    .ZN(_01313_));
 BUF_X4 _37113_ (.A(_13994_),
    .Z(_14037_));
 NAND2_X1 _37114_ (.A1(\core.keymem.key_mem[12][69] ),
    .A2(_14037_),
    .ZN(_14038_));
 OAI21_X1 _37115_ (.A(_14038_),
    .B1(_14029_),
    .B2(_13700_),
    .ZN(_01314_));
 MUX2_X1 _37116_ (.A(\core.keymem.key_mem[12][6] ),
    .B(_13711_),
    .S(_14033_),
    .Z(_01315_));
 MUX2_X1 _37117_ (.A(\core.keymem.key_mem[12][70] ),
    .B(_13713_),
    .S(_14033_),
    .Z(_01316_));
 NAND2_X1 _37118_ (.A1(\core.keymem.key_mem[12][71] ),
    .A2(_14037_),
    .ZN(_14039_));
 OAI21_X1 _37119_ (.A(_14039_),
    .B1(_14029_),
    .B2(_12659_),
    .ZN(_01317_));
 NAND2_X1 _37120_ (.A1(\core.keymem.key_mem[12][72] ),
    .A2(_14037_),
    .ZN(_14040_));
 OAI21_X1 _37121_ (.A(_14040_),
    .B1(_14029_),
    .B2(_13716_),
    .ZN(_01318_));
 NAND2_X1 _37122_ (.A1(\core.keymem.key_mem[12][73] ),
    .A2(_14037_),
    .ZN(_14041_));
 BUF_X4 _37123_ (.A(_13997_),
    .Z(_14042_));
 OAI21_X1 _37124_ (.A(_14041_),
    .B1(_14042_),
    .B2(_12688_),
    .ZN(_01319_));
 NAND2_X1 _37125_ (.A1(\core.keymem.key_mem[12][74] ),
    .A2(_14037_),
    .ZN(_14043_));
 OAI21_X1 _37126_ (.A(_14043_),
    .B1(_14042_),
    .B2(_13726_),
    .ZN(_01320_));
 NAND2_X1 _37127_ (.A1(\core.keymem.key_mem[12][75] ),
    .A2(_14037_),
    .ZN(_14044_));
 OAI21_X1 _37128_ (.A(_14044_),
    .B1(_14042_),
    .B2(_13733_),
    .ZN(_01321_));
 BUF_X4 _37129_ (.A(_13990_),
    .Z(_14045_));
 MUX2_X1 _37130_ (.A(\core.keymem.key_mem[12][76] ),
    .B(_13741_),
    .S(_14045_),
    .Z(_01322_));
 MUX2_X1 _37131_ (.A(\core.keymem.key_mem[12][77] ),
    .B(_13751_),
    .S(_14045_),
    .Z(_01323_));
 NAND2_X1 _37132_ (.A1(\core.keymem.key_mem[12][78] ),
    .A2(_14037_),
    .ZN(_14046_));
 OAI21_X1 _37133_ (.A(_14046_),
    .B1(_14042_),
    .B2(_12708_),
    .ZN(_01324_));
 MUX2_X1 _37134_ (.A(\core.keymem.key_mem[12][79] ),
    .B(_13758_),
    .S(_14045_),
    .Z(_01325_));
 NAND2_X1 _37135_ (.A1(\core.keymem.key_mem[12][7] ),
    .A2(_14037_),
    .ZN(_14047_));
 OAI21_X1 _37136_ (.A(_14047_),
    .B1(_14042_),
    .B2(_13767_),
    .ZN(_01326_));
 MUX2_X1 _37137_ (.A(\core.keymem.key_mem[12][80] ),
    .B(_13769_),
    .S(_14045_),
    .Z(_01327_));
 NAND2_X1 _37138_ (.A1(\core.keymem.key_mem[12][81] ),
    .A2(_14037_),
    .ZN(_14048_));
 OAI21_X1 _37139_ (.A(_14048_),
    .B1(_14042_),
    .B2(_13775_),
    .ZN(_01328_));
 NAND2_X1 _37140_ (.A1(\core.keymem.key_mem[12][82] ),
    .A2(_14037_),
    .ZN(_14049_));
 OAI21_X1 _37141_ (.A(_14049_),
    .B1(_14042_),
    .B2(_13783_),
    .ZN(_01329_));
 NAND2_X1 _37142_ (.A1(\core.keymem.key_mem[12][83] ),
    .A2(_13997_),
    .ZN(_14050_));
 OAI21_X1 _37143_ (.A(_14050_),
    .B1(_14042_),
    .B2(_13791_),
    .ZN(_01330_));
 NAND2_X1 _37144_ (.A1(\core.keymem.key_mem[12][84] ),
    .A2(_13997_),
    .ZN(_14051_));
 OAI21_X1 _37145_ (.A(_14051_),
    .B1(_14042_),
    .B2(_12725_),
    .ZN(_01331_));
 MUX2_X1 _37146_ (.A(\core.keymem.key_mem[12][85] ),
    .B(_13798_),
    .S(_14045_),
    .Z(_01332_));
 MUX2_X1 _37147_ (.A(\core.keymem.key_mem[12][86] ),
    .B(_12741_),
    .S(_14045_),
    .Z(_01333_));
 MUX2_X1 _37148_ (.A(\core.keymem.key_mem[12][87] ),
    .B(_13804_),
    .S(_14045_),
    .Z(_01334_));
 MUX2_X1 _37149_ (.A(\core.keymem.key_mem[12][88] ),
    .B(_13810_),
    .S(_14045_),
    .Z(_01335_));
 MUX2_X1 _37150_ (.A(\core.keymem.key_mem[12][89] ),
    .B(_13818_),
    .S(_14045_),
    .Z(_01336_));
 MUX2_X1 _37151_ (.A(\core.keymem.key_mem[12][8] ),
    .B(_13854_),
    .S(_14045_),
    .Z(_01337_));
 MUX2_X1 _37152_ (.A(\core.keymem.key_mem[12][90] ),
    .B(_13860_),
    .S(_13991_),
    .Z(_01338_));
 NAND2_X1 _37153_ (.A1(\core.keymem.key_mem[12][91] ),
    .A2(_13997_),
    .ZN(_14052_));
 OAI21_X1 _37154_ (.A(_14052_),
    .B1(_14042_),
    .B2(_13870_),
    .ZN(_01339_));
 NAND2_X1 _37155_ (.A1(\core.keymem.key_mem[12][92] ),
    .A2(_13997_),
    .ZN(_14053_));
 OAI21_X1 _37156_ (.A(_14053_),
    .B1(_13995_),
    .B2(_13880_),
    .ZN(_01340_));
 MUX2_X1 _37157_ (.A(\core.keymem.key_mem[12][93] ),
    .B(_13889_),
    .S(_13991_),
    .Z(_01341_));
 MUX2_X1 _37158_ (.A(\core.keymem.key_mem[12][94] ),
    .B(_13896_),
    .S(_13991_),
    .Z(_01342_));
 MUX2_X1 _37159_ (.A(\core.keymem.key_mem[12][95] ),
    .B(_13903_),
    .S(_13991_),
    .Z(_01343_));
 MUX2_X1 _37160_ (.A(\core.keymem.key_mem[12][96] ),
    .B(_13907_),
    .S(_13991_),
    .Z(_01344_));
 NAND2_X1 _37161_ (.A1(\core.keymem.key_mem[12][97] ),
    .A2(_13997_),
    .ZN(_14054_));
 OAI21_X1 _37162_ (.A(_14054_),
    .B1(_13995_),
    .B2(_12777_),
    .ZN(_01345_));
 NAND2_X1 _37163_ (.A1(\core.keymem.key_mem[12][98] ),
    .A2(_13997_),
    .ZN(_14055_));
 OAI21_X1 _37164_ (.A(_14055_),
    .B1(_13995_),
    .B2(_13910_),
    .ZN(_01346_));
 MUX2_X1 _37165_ (.A(\core.keymem.key_mem[12][99] ),
    .B(_12800_),
    .S(_13991_),
    .Z(_01347_));
 MUX2_X1 _37166_ (.A(\core.keymem.key_mem[12][9] ),
    .B(_13919_),
    .S(_13991_),
    .Z(_01348_));
 NAND2_X4 _37167_ (.A1(_16222_),
    .A2(_11816_),
    .ZN(_14056_));
 NOR2_X4 _37168_ (.A1(_13988_),
    .A2(_14056_),
    .ZN(_14057_));
 BUF_X4 _37169_ (.A(_14057_),
    .Z(_14058_));
 BUF_X4 _37170_ (.A(_14058_),
    .Z(_14059_));
 MUX2_X1 _37171_ (.A(\core.keymem.key_mem[13][0] ),
    .B(_11844_),
    .S(_14059_),
    .Z(_01349_));
 MUX2_X1 _37172_ (.A(\core.keymem.key_mem[13][100] ),
    .B(_11873_),
    .S(_14059_),
    .Z(_01350_));
 MUX2_X1 _37173_ (.A(\core.keymem.key_mem[13][101] ),
    .B(_12813_),
    .S(_14059_),
    .Z(_01351_));
 MUX2_X1 _37174_ (.A(\core.keymem.key_mem[13][102] ),
    .B(_11906_),
    .S(_14059_),
    .Z(_01352_));
 MUX2_X1 _37175_ (.A(\core.keymem.key_mem[13][103] ),
    .B(_11929_),
    .S(_14059_),
    .Z(_01353_));
 OR2_X1 _37176_ (.A1(_13988_),
    .A2(_14056_),
    .ZN(_14060_));
 CLKBUF_X3 _37177_ (.A(_14060_),
    .Z(_14061_));
 BUF_X4 _37178_ (.A(_14061_),
    .Z(_14062_));
 NAND2_X1 _37179_ (.A1(\core.keymem.key_mem[13][104] ),
    .A2(_14062_),
    .ZN(_14063_));
 BUF_X4 _37180_ (.A(_14061_),
    .Z(_14064_));
 BUF_X4 _37181_ (.A(_14064_),
    .Z(_14065_));
 OAI21_X1 _37182_ (.A(_14063_),
    .B1(_14065_),
    .B2(_12822_),
    .ZN(_01354_));
 MUX2_X1 _37183_ (.A(\core.keymem.key_mem[13][105] ),
    .B(_12830_),
    .S(_14059_),
    .Z(_01355_));
 BUF_X4 _37184_ (.A(_14058_),
    .Z(_14066_));
 MUX2_X1 _37185_ (.A(\core.keymem.key_mem[13][106] ),
    .B(_12832_),
    .S(_14066_),
    .Z(_01356_));
 MUX2_X1 _37186_ (.A(\core.keymem.key_mem[13][107] ),
    .B(_11967_),
    .S(_14066_),
    .Z(_01357_));
 MUX2_X1 _37187_ (.A(\core.keymem.key_mem[13][108] ),
    .B(_11981_),
    .S(_14066_),
    .Z(_01358_));
 MUX2_X1 _37188_ (.A(\core.keymem.key_mem[13][109] ),
    .B(_12842_),
    .S(_14066_),
    .Z(_01359_));
 NAND2_X1 _37189_ (.A1(\core.keymem.key_mem[13][10] ),
    .A2(_14062_),
    .ZN(_14067_));
 OAI21_X1 _37190_ (.A(_14067_),
    .B1(_14065_),
    .B2(_12858_),
    .ZN(_01360_));
 MUX2_X1 _37191_ (.A(\core.keymem.key_mem[13][110] ),
    .B(_12859_),
    .S(_14066_),
    .Z(_01361_));
 MUX2_X1 _37192_ (.A(\core.keymem.key_mem[13][111] ),
    .B(_12017_),
    .S(_14066_),
    .Z(_01362_));
 MUX2_X1 _37193_ (.A(\core.keymem.key_mem[13][112] ),
    .B(_12031_),
    .S(_14066_),
    .Z(_01363_));
 MUX2_X1 _37194_ (.A(\core.keymem.key_mem[13][113] ),
    .B(_12868_),
    .S(_14066_),
    .Z(_01364_));
 MUX2_X1 _37195_ (.A(\core.keymem.key_mem[13][114] ),
    .B(_12869_),
    .S(_14066_),
    .Z(_01365_));
 MUX2_X1 _37196_ (.A(\core.keymem.key_mem[13][115] ),
    .B(_12059_),
    .S(_14066_),
    .Z(_01366_));
 BUF_X4 _37197_ (.A(_14058_),
    .Z(_14068_));
 MUX2_X1 _37198_ (.A(\core.keymem.key_mem[13][116] ),
    .B(_12077_),
    .S(_14068_),
    .Z(_01367_));
 MUX2_X1 _37199_ (.A(\core.keymem.key_mem[13][117] ),
    .B(_12877_),
    .S(_14068_),
    .Z(_01368_));
 MUX2_X1 _37200_ (.A(\core.keymem.key_mem[13][118] ),
    .B(_12882_),
    .S(_14068_),
    .Z(_01369_));
 MUX2_X1 _37201_ (.A(\core.keymem.key_mem[13][119] ),
    .B(_12096_),
    .S(_14068_),
    .Z(_01370_));
 NAND2_X1 _37202_ (.A1(\core.keymem.key_mem[13][11] ),
    .A2(_14062_),
    .ZN(_14069_));
 OAI21_X1 _37203_ (.A(_14069_),
    .B1(_14065_),
    .B2(_12895_),
    .ZN(_01371_));
 MUX2_X1 _37204_ (.A(\core.keymem.key_mem[13][120] ),
    .B(_12124_),
    .S(_14068_),
    .Z(_01372_));
 MUX2_X1 _37205_ (.A(\core.keymem.key_mem[13][121] ),
    .B(_12160_),
    .S(_14068_),
    .Z(_01373_));
 MUX2_X1 _37206_ (.A(\core.keymem.key_mem[13][122] ),
    .B(_12903_),
    .S(_14068_),
    .Z(_01374_));
 NAND2_X1 _37207_ (.A1(\core.keymem.key_mem[13][123] ),
    .A2(_14062_),
    .ZN(_14070_));
 OAI21_X1 _37208_ (.A(_14070_),
    .B1(_14065_),
    .B2(_12182_),
    .ZN(_01375_));
 NAND2_X1 _37209_ (.A1(\core.keymem.key_mem[13][124] ),
    .A2(_14062_),
    .ZN(_14071_));
 OAI21_X1 _37210_ (.A(_14071_),
    .B1(_14065_),
    .B2(_12926_),
    .ZN(_01376_));
 MUX2_X1 _37211_ (.A(\core.keymem.key_mem[13][125] ),
    .B(_12932_),
    .S(_14068_),
    .Z(_01377_));
 NAND2_X1 _37212_ (.A1(\core.keymem.key_mem[13][126] ),
    .A2(_14062_),
    .ZN(_14072_));
 OAI21_X1 _37213_ (.A(_14072_),
    .B1(_14065_),
    .B2(_12207_),
    .ZN(_01378_));
 MUX2_X1 _37214_ (.A(\core.keymem.key_mem[13][127] ),
    .B(_12945_),
    .S(_14068_),
    .Z(_01379_));
 MUX2_X1 _37215_ (.A(\core.keymem.key_mem[13][12] ),
    .B(_12958_),
    .S(_14068_),
    .Z(_01380_));
 BUF_X4 _37216_ (.A(_14057_),
    .Z(_14073_));
 MUX2_X1 _37217_ (.A(\core.keymem.key_mem[13][13] ),
    .B(_12974_),
    .S(_14073_),
    .Z(_01381_));
 NOR2_X1 _37218_ (.A1(\core.keymem.key_mem[13][14] ),
    .A2(_14059_),
    .ZN(_14074_));
 AOI21_X1 _37219_ (.A(_14074_),
    .B1(_14059_),
    .B2(_13007_),
    .ZN(_01382_));
 MUX2_X1 _37220_ (.A(\core.keymem.key_mem[13][15] ),
    .B(_13017_),
    .S(_14073_),
    .Z(_01383_));
 MUX2_X1 _37221_ (.A(\core.keymem.key_mem[13][16] ),
    .B(_13029_),
    .S(_14073_),
    .Z(_01384_));
 NAND2_X1 _37222_ (.A1(\core.keymem.key_mem[13][17] ),
    .A2(_14062_),
    .ZN(_14075_));
 OAI21_X1 _37223_ (.A(_14075_),
    .B1(_14065_),
    .B2(_13042_),
    .ZN(_01385_));
 MUX2_X1 _37224_ (.A(\core.keymem.key_mem[13][18] ),
    .B(_13094_),
    .S(_14073_),
    .Z(_01386_));
 BUF_X4 _37225_ (.A(_14061_),
    .Z(_14076_));
 NAND2_X1 _37226_ (.A1(\core.keymem.key_mem[13][19] ),
    .A2(_14076_),
    .ZN(_14077_));
 OAI21_X1 _37227_ (.A(_14077_),
    .B1(_14065_),
    .B2(_13109_),
    .ZN(_01387_));
 MUX2_X1 _37228_ (.A(\core.keymem.key_mem[13][1] ),
    .B(_13134_),
    .S(_14073_),
    .Z(_01388_));
 MUX2_X1 _37229_ (.A(\core.keymem.key_mem[13][20] ),
    .B(_13146_),
    .S(_14073_),
    .Z(_01389_));
 MUX2_X1 _37230_ (.A(\core.keymem.key_mem[13][21] ),
    .B(_13155_),
    .S(_14073_),
    .Z(_01390_));
 NOR2_X1 _37231_ (.A1(\core.keymem.key_mem[13][22] ),
    .A2(_14059_),
    .ZN(_14078_));
 AOI21_X1 _37232_ (.A(_14078_),
    .B1(_14059_),
    .B2(_13191_),
    .ZN(_01391_));
 MUX2_X1 _37233_ (.A(\core.keymem.key_mem[13][23] ),
    .B(_13196_),
    .S(_14073_),
    .Z(_01392_));
 NAND2_X1 _37234_ (.A1(\core.keymem.key_mem[13][24] ),
    .A2(_14076_),
    .ZN(_14079_));
 OAI21_X1 _37235_ (.A(_14079_),
    .B1(_14065_),
    .B2(_13212_),
    .ZN(_01393_));
 MUX2_X1 _37236_ (.A(\core.keymem.key_mem[13][25] ),
    .B(_13233_),
    .S(_14073_),
    .Z(_01394_));
 MUX2_X1 _37237_ (.A(\core.keymem.key_mem[13][26] ),
    .B(_13241_),
    .S(_14073_),
    .Z(_01395_));
 BUF_X4 _37238_ (.A(_14057_),
    .Z(_14080_));
 MUX2_X1 _37239_ (.A(\core.keymem.key_mem[13][27] ),
    .B(_13284_),
    .S(_14080_),
    .Z(_01396_));
 MUX2_X1 _37240_ (.A(\core.keymem.key_mem[13][28] ),
    .B(_13325_),
    .S(_14080_),
    .Z(_01397_));
 MUX2_X1 _37241_ (.A(\core.keymem.key_mem[13][29] ),
    .B(_13329_),
    .S(_14080_),
    .Z(_01398_));
 NAND2_X1 _37242_ (.A1(\core.keymem.key_mem[13][2] ),
    .A2(_14076_),
    .ZN(_14081_));
 OAI21_X1 _37243_ (.A(_14081_),
    .B1(_14065_),
    .B2(_13335_),
    .ZN(_01399_));
 MUX2_X1 _37244_ (.A(\core.keymem.key_mem[13][30] ),
    .B(_13379_),
    .S(_14080_),
    .Z(_01400_));
 MUX2_X1 _37245_ (.A(\core.keymem.key_mem[13][31] ),
    .B(_13395_),
    .S(_14080_),
    .Z(_01401_));
 MUX2_X1 _37246_ (.A(\core.keymem.key_mem[13][32] ),
    .B(_13396_),
    .S(_14080_),
    .Z(_01402_));
 MUX2_X1 _37247_ (.A(\core.keymem.key_mem[13][33] ),
    .B(_13402_),
    .S(_14080_),
    .Z(_01403_));
 MUX2_X1 _37248_ (.A(\core.keymem.key_mem[13][34] ),
    .B(_13403_),
    .S(_14080_),
    .Z(_01404_));
 MUX2_X1 _37249_ (.A(\core.keymem.key_mem[13][35] ),
    .B(_13405_),
    .S(_14080_),
    .Z(_01405_));
 NAND2_X1 _37250_ (.A1(\core.keymem.key_mem[13][36] ),
    .A2(_14076_),
    .ZN(_14082_));
 BUF_X4 _37251_ (.A(_14064_),
    .Z(_14083_));
 OAI21_X1 _37252_ (.A(_14082_),
    .B1(_14083_),
    .B2(_13407_),
    .ZN(_01406_));
 NAND2_X1 _37253_ (.A1(\core.keymem.key_mem[13][37] ),
    .A2(_14076_),
    .ZN(_14084_));
 OAI21_X1 _37254_ (.A(_14084_),
    .B1(_14083_),
    .B2(_12439_),
    .ZN(_01407_));
 MUX2_X1 _37255_ (.A(\core.keymem.key_mem[13][38] ),
    .B(_13410_),
    .S(_14080_),
    .Z(_01408_));
 NAND2_X1 _37256_ (.A1(\core.keymem.key_mem[13][39] ),
    .A2(_14076_),
    .ZN(_14085_));
 OAI21_X1 _37257_ (.A(_14085_),
    .B1(_14083_),
    .B2(_13435_),
    .ZN(_01409_));
 NAND2_X1 _37258_ (.A1(\core.keymem.key_mem[13][3] ),
    .A2(_14076_),
    .ZN(_14086_));
 OAI21_X1 _37259_ (.A(_14086_),
    .B1(_14083_),
    .B2(_13448_),
    .ZN(_01410_));
 NAND2_X1 _37260_ (.A1(\core.keymem.key_mem[13][40] ),
    .A2(_14076_),
    .ZN(_14087_));
 OAI21_X1 _37261_ (.A(_14087_),
    .B1(_14083_),
    .B2(_13457_),
    .ZN(_01411_));
 BUF_X4 _37262_ (.A(_14057_),
    .Z(_14088_));
 MUX2_X1 _37263_ (.A(\core.keymem.key_mem[13][41] ),
    .B(_13467_),
    .S(_14088_),
    .Z(_01412_));
 MUX2_X1 _37264_ (.A(\core.keymem.key_mem[13][42] ),
    .B(_13490_),
    .S(_14088_),
    .Z(_01413_));
 NAND2_X1 _37265_ (.A1(\core.keymem.key_mem[13][43] ),
    .A2(_14076_),
    .ZN(_14089_));
 OAI21_X1 _37266_ (.A(_14089_),
    .B1(_14083_),
    .B2(_13496_),
    .ZN(_01414_));
 MUX2_X1 _37267_ (.A(\core.keymem.key_mem[13][44] ),
    .B(_13497_),
    .S(_14088_),
    .Z(_01415_));
 NAND2_X1 _37268_ (.A1(\core.keymem.key_mem[13][45] ),
    .A2(_14076_),
    .ZN(_14090_));
 OAI21_X1 _37269_ (.A(_14090_),
    .B1(_14083_),
    .B2(_13510_),
    .ZN(_01416_));
 BUF_X4 _37270_ (.A(_14061_),
    .Z(_14091_));
 NAND2_X1 _37271_ (.A1(\core.keymem.key_mem[13][46] ),
    .A2(_14091_),
    .ZN(_14092_));
 OAI21_X1 _37272_ (.A(_14092_),
    .B1(_14083_),
    .B2(_13517_),
    .ZN(_01417_));
 NAND2_X1 _37273_ (.A1(\core.keymem.key_mem[13][47] ),
    .A2(_14091_),
    .ZN(_14093_));
 OAI21_X1 _37274_ (.A(_14093_),
    .B1(_14083_),
    .B2(_12520_),
    .ZN(_01418_));
 NAND2_X1 _37275_ (.A1(\core.keymem.key_mem[13][48] ),
    .A2(_14091_),
    .ZN(_14094_));
 OAI21_X1 _37276_ (.A(_14094_),
    .B1(_14083_),
    .B2(_12532_),
    .ZN(_01419_));
 NAND2_X1 _37277_ (.A1(\core.keymem.key_mem[13][49] ),
    .A2(_14091_),
    .ZN(_14095_));
 BUF_X4 _37278_ (.A(_14064_),
    .Z(_14096_));
 OAI21_X1 _37279_ (.A(_14095_),
    .B1(_14096_),
    .B2(_13529_),
    .ZN(_01420_));
 MUX2_X1 _37280_ (.A(\core.keymem.key_mem[13][4] ),
    .B(_13538_),
    .S(_14088_),
    .Z(_01421_));
 MUX2_X1 _37281_ (.A(\core.keymem.key_mem[13][50] ),
    .B(_13557_),
    .S(_14088_),
    .Z(_01422_));
 MUX2_X1 _37282_ (.A(\core.keymem.key_mem[13][51] ),
    .B(_13564_),
    .S(_14088_),
    .Z(_01423_));
 NAND2_X1 _37283_ (.A1(\core.keymem.key_mem[13][52] ),
    .A2(_14091_),
    .ZN(_14097_));
 OAI21_X1 _37284_ (.A(_14097_),
    .B1(_14096_),
    .B2(_12568_),
    .ZN(_01424_));
 NAND2_X1 _37285_ (.A1(\core.keymem.key_mem[13][53] ),
    .A2(_14091_),
    .ZN(_14098_));
 OAI21_X1 _37286_ (.A(_14098_),
    .B1(_14096_),
    .B2(_12584_),
    .ZN(_01425_));
 NAND2_X1 _37287_ (.A1(\core.keymem.key_mem[13][54] ),
    .A2(_14091_),
    .ZN(_14099_));
 OAI21_X1 _37288_ (.A(_14099_),
    .B1(_14096_),
    .B2(_13575_),
    .ZN(_01426_));
 MUX2_X1 _37289_ (.A(\core.keymem.key_mem[13][55] ),
    .B(_13581_),
    .S(_14088_),
    .Z(_01427_));
 MUX2_X1 _37290_ (.A(\core.keymem.key_mem[13][56] ),
    .B(_13589_),
    .S(_14088_),
    .Z(_01428_));
 MUX2_X1 _37291_ (.A(\core.keymem.key_mem[13][57] ),
    .B(_13604_),
    .S(_14088_),
    .Z(_01429_));
 MUX2_X1 _37292_ (.A(\core.keymem.key_mem[13][58] ),
    .B(_13611_),
    .S(_14088_),
    .Z(_01430_));
 BUF_X4 _37293_ (.A(_14057_),
    .Z(_14100_));
 MUX2_X1 _37294_ (.A(\core.keymem.key_mem[13][59] ),
    .B(_13616_),
    .S(_14100_),
    .Z(_01431_));
 MUX2_X1 _37295_ (.A(\core.keymem.key_mem[13][5] ),
    .B(_12606_),
    .S(_14100_),
    .Z(_01432_));
 MUX2_X1 _37296_ (.A(\core.keymem.key_mem[13][60] ),
    .B(_13622_),
    .S(_14100_),
    .Z(_01433_));
 MUX2_X1 _37297_ (.A(\core.keymem.key_mem[13][61] ),
    .B(_13632_),
    .S(_14100_),
    .Z(_01434_));
 MUX2_X1 _37298_ (.A(\core.keymem.key_mem[13][62] ),
    .B(_13637_),
    .S(_14100_),
    .Z(_01435_));
 MUX2_X1 _37299_ (.A(\core.keymem.key_mem[13][63] ),
    .B(_13659_),
    .S(_14100_),
    .Z(_01436_));
 MUX2_X1 _37300_ (.A(\core.keymem.key_mem[13][64] ),
    .B(_12622_),
    .S(_14100_),
    .Z(_01437_));
 NAND2_X1 _37301_ (.A1(\core.keymem.key_mem[13][65] ),
    .A2(_14091_),
    .ZN(_14101_));
 OAI21_X1 _37302_ (.A(_14101_),
    .B1(_14096_),
    .B2(_13673_),
    .ZN(_01438_));
 MUX2_X1 _37303_ (.A(\core.keymem.key_mem[13][66] ),
    .B(_13681_),
    .S(_14100_),
    .Z(_01439_));
 NAND2_X1 _37304_ (.A1(\core.keymem.key_mem[13][67] ),
    .A2(_14091_),
    .ZN(_14102_));
 OAI21_X1 _37305_ (.A(_14102_),
    .B1(_14096_),
    .B2(_13690_),
    .ZN(_01440_));
 NAND2_X1 _37306_ (.A1(\core.keymem.key_mem[13][68] ),
    .A2(_14091_),
    .ZN(_14103_));
 OAI21_X1 _37307_ (.A(_14103_),
    .B1(_14096_),
    .B2(_12635_),
    .ZN(_01441_));
 BUF_X4 _37308_ (.A(_14061_),
    .Z(_14104_));
 NAND2_X1 _37309_ (.A1(\core.keymem.key_mem[13][69] ),
    .A2(_14104_),
    .ZN(_14105_));
 OAI21_X1 _37310_ (.A(_14105_),
    .B1(_14096_),
    .B2(_13700_),
    .ZN(_01442_));
 MUX2_X1 _37311_ (.A(\core.keymem.key_mem[13][6] ),
    .B(_13711_),
    .S(_14100_),
    .Z(_01443_));
 MUX2_X1 _37312_ (.A(\core.keymem.key_mem[13][70] ),
    .B(_13713_),
    .S(_14100_),
    .Z(_01444_));
 NAND2_X1 _37313_ (.A1(\core.keymem.key_mem[13][71] ),
    .A2(_14104_),
    .ZN(_14106_));
 OAI21_X1 _37314_ (.A(_14106_),
    .B1(_14096_),
    .B2(_12659_),
    .ZN(_01445_));
 NAND2_X1 _37315_ (.A1(\core.keymem.key_mem[13][72] ),
    .A2(_14104_),
    .ZN(_14107_));
 OAI21_X1 _37316_ (.A(_14107_),
    .B1(_14096_),
    .B2(_13716_),
    .ZN(_01446_));
 NAND2_X1 _37317_ (.A1(\core.keymem.key_mem[13][73] ),
    .A2(_14104_),
    .ZN(_14108_));
 BUF_X4 _37318_ (.A(_14064_),
    .Z(_14109_));
 OAI21_X1 _37319_ (.A(_14108_),
    .B1(_14109_),
    .B2(_12688_),
    .ZN(_01447_));
 NAND2_X1 _37320_ (.A1(\core.keymem.key_mem[13][74] ),
    .A2(_14104_),
    .ZN(_14110_));
 OAI21_X1 _37321_ (.A(_14110_),
    .B1(_14109_),
    .B2(_13726_),
    .ZN(_01448_));
 NAND2_X1 _37322_ (.A1(\core.keymem.key_mem[13][75] ),
    .A2(_14104_),
    .ZN(_14111_));
 OAI21_X1 _37323_ (.A(_14111_),
    .B1(_14109_),
    .B2(_13733_),
    .ZN(_01449_));
 BUF_X4 _37324_ (.A(_14057_),
    .Z(_14112_));
 MUX2_X1 _37325_ (.A(\core.keymem.key_mem[13][76] ),
    .B(_13741_),
    .S(_14112_),
    .Z(_01450_));
 MUX2_X1 _37326_ (.A(\core.keymem.key_mem[13][77] ),
    .B(_13751_),
    .S(_14112_),
    .Z(_01451_));
 NAND2_X1 _37327_ (.A1(\core.keymem.key_mem[13][78] ),
    .A2(_14104_),
    .ZN(_14113_));
 OAI21_X1 _37328_ (.A(_14113_),
    .B1(_14109_),
    .B2(_12708_),
    .ZN(_01452_));
 MUX2_X1 _37329_ (.A(\core.keymem.key_mem[13][79] ),
    .B(_13758_),
    .S(_14112_),
    .Z(_01453_));
 NAND2_X1 _37330_ (.A1(\core.keymem.key_mem[13][7] ),
    .A2(_14104_),
    .ZN(_14114_));
 OAI21_X1 _37331_ (.A(_14114_),
    .B1(_14109_),
    .B2(_13767_),
    .ZN(_01454_));
 MUX2_X1 _37332_ (.A(\core.keymem.key_mem[13][80] ),
    .B(_13769_),
    .S(_14112_),
    .Z(_01455_));
 NAND2_X1 _37333_ (.A1(\core.keymem.key_mem[13][81] ),
    .A2(_14104_),
    .ZN(_14115_));
 OAI21_X1 _37334_ (.A(_14115_),
    .B1(_14109_),
    .B2(_13775_),
    .ZN(_01456_));
 NAND2_X1 _37335_ (.A1(\core.keymem.key_mem[13][82] ),
    .A2(_14104_),
    .ZN(_14116_));
 OAI21_X1 _37336_ (.A(_14116_),
    .B1(_14109_),
    .B2(_13783_),
    .ZN(_01457_));
 NAND2_X1 _37337_ (.A1(\core.keymem.key_mem[13][83] ),
    .A2(_14064_),
    .ZN(_14117_));
 OAI21_X1 _37338_ (.A(_14117_),
    .B1(_14109_),
    .B2(_13791_),
    .ZN(_01458_));
 NAND2_X1 _37339_ (.A1(\core.keymem.key_mem[13][84] ),
    .A2(_14064_),
    .ZN(_14118_));
 OAI21_X1 _37340_ (.A(_14118_),
    .B1(_14109_),
    .B2(_12725_),
    .ZN(_01459_));
 MUX2_X1 _37341_ (.A(\core.keymem.key_mem[13][85] ),
    .B(_13798_),
    .S(_14112_),
    .Z(_01460_));
 MUX2_X1 _37342_ (.A(\core.keymem.key_mem[13][86] ),
    .B(_12741_),
    .S(_14112_),
    .Z(_01461_));
 MUX2_X1 _37343_ (.A(\core.keymem.key_mem[13][87] ),
    .B(_13804_),
    .S(_14112_),
    .Z(_01462_));
 MUX2_X1 _37344_ (.A(\core.keymem.key_mem[13][88] ),
    .B(_13810_),
    .S(_14112_),
    .Z(_01463_));
 MUX2_X1 _37345_ (.A(\core.keymem.key_mem[13][89] ),
    .B(_13818_),
    .S(_14112_),
    .Z(_01464_));
 MUX2_X1 _37346_ (.A(\core.keymem.key_mem[13][8] ),
    .B(_13854_),
    .S(_14112_),
    .Z(_01465_));
 MUX2_X1 _37347_ (.A(\core.keymem.key_mem[13][90] ),
    .B(_13860_),
    .S(_14058_),
    .Z(_01466_));
 NAND2_X1 _37348_ (.A1(\core.keymem.key_mem[13][91] ),
    .A2(_14064_),
    .ZN(_14119_));
 OAI21_X1 _37349_ (.A(_14119_),
    .B1(_14109_),
    .B2(_13870_),
    .ZN(_01467_));
 NAND2_X1 _37350_ (.A1(\core.keymem.key_mem[13][92] ),
    .A2(_14064_),
    .ZN(_14120_));
 OAI21_X1 _37351_ (.A(_14120_),
    .B1(_14062_),
    .B2(_13880_),
    .ZN(_01468_));
 MUX2_X1 _37352_ (.A(\core.keymem.key_mem[13][93] ),
    .B(_13889_),
    .S(_14058_),
    .Z(_01469_));
 MUX2_X1 _37353_ (.A(\core.keymem.key_mem[13][94] ),
    .B(_13896_),
    .S(_14058_),
    .Z(_01470_));
 MUX2_X1 _37354_ (.A(\core.keymem.key_mem[13][95] ),
    .B(_13903_),
    .S(_14058_),
    .Z(_01471_));
 MUX2_X1 _37355_ (.A(\core.keymem.key_mem[13][96] ),
    .B(_13907_),
    .S(_14058_),
    .Z(_01472_));
 NAND2_X1 _37356_ (.A1(\core.keymem.key_mem[13][97] ),
    .A2(_14064_),
    .ZN(_14121_));
 OAI21_X1 _37357_ (.A(_14121_),
    .B1(_14062_),
    .B2(_12777_),
    .ZN(_01473_));
 NAND2_X1 _37358_ (.A1(\core.keymem.key_mem[13][98] ),
    .A2(_14064_),
    .ZN(_14122_));
 OAI21_X1 _37359_ (.A(_14122_),
    .B1(_14062_),
    .B2(_13910_),
    .ZN(_01474_));
 MUX2_X1 _37360_ (.A(\core.keymem.key_mem[13][99] ),
    .B(_12800_),
    .S(_14058_),
    .Z(_01475_));
 MUX2_X1 _37361_ (.A(\core.keymem.key_mem[13][9] ),
    .B(_13919_),
    .S(_14058_),
    .Z(_01476_));
 NOR2_X4 _37362_ (.A1(_12804_),
    .A2(_13988_),
    .ZN(_14123_));
 BUF_X4 _37363_ (.A(_14123_),
    .Z(_14124_));
 BUF_X4 _37364_ (.A(_14124_),
    .Z(_14125_));
 MUX2_X1 _37365_ (.A(\core.keymem.key_mem[14][0] ),
    .B(_11844_),
    .S(_14125_),
    .Z(_01477_));
 MUX2_X1 _37366_ (.A(\core.keymem.key_mem[14][100] ),
    .B(_11873_),
    .S(_14125_),
    .Z(_01478_));
 MUX2_X1 _37367_ (.A(\core.keymem.key_mem[14][101] ),
    .B(_12813_),
    .S(_14125_),
    .Z(_01479_));
 MUX2_X1 _37368_ (.A(\core.keymem.key_mem[14][102] ),
    .B(_11906_),
    .S(_14125_),
    .Z(_01480_));
 MUX2_X1 _37369_ (.A(\core.keymem.key_mem[14][103] ),
    .B(_11929_),
    .S(_14125_),
    .Z(_01481_));
 OR2_X1 _37370_ (.A1(_12804_),
    .A2(_13988_),
    .ZN(_14126_));
 CLKBUF_X3 _37371_ (.A(_14126_),
    .Z(_14127_));
 BUF_X4 _37372_ (.A(_14127_),
    .Z(_14128_));
 NAND2_X1 _37373_ (.A1(\core.keymem.key_mem[14][104] ),
    .A2(_14128_),
    .ZN(_14129_));
 BUF_X4 _37374_ (.A(_14127_),
    .Z(_14130_));
 BUF_X4 _37375_ (.A(_14130_),
    .Z(_14131_));
 OAI21_X1 _37376_ (.A(_14129_),
    .B1(_14131_),
    .B2(_12822_),
    .ZN(_01482_));
 MUX2_X1 _37377_ (.A(\core.keymem.key_mem[14][105] ),
    .B(_12830_),
    .S(_14125_),
    .Z(_01483_));
 BUF_X4 _37378_ (.A(_14124_),
    .Z(_14132_));
 MUX2_X1 _37379_ (.A(\core.keymem.key_mem[14][106] ),
    .B(_12832_),
    .S(_14132_),
    .Z(_01484_));
 MUX2_X1 _37380_ (.A(\core.keymem.key_mem[14][107] ),
    .B(_11967_),
    .S(_14132_),
    .Z(_01485_));
 MUX2_X1 _37381_ (.A(\core.keymem.key_mem[14][108] ),
    .B(_11981_),
    .S(_14132_),
    .Z(_01486_));
 MUX2_X1 _37382_ (.A(\core.keymem.key_mem[14][109] ),
    .B(_12842_),
    .S(_14132_),
    .Z(_01487_));
 NAND2_X1 _37383_ (.A1(\core.keymem.key_mem[14][10] ),
    .A2(_14128_),
    .ZN(_14133_));
 OAI21_X1 _37384_ (.A(_14133_),
    .B1(_14131_),
    .B2(_12858_),
    .ZN(_01488_));
 MUX2_X1 _37385_ (.A(\core.keymem.key_mem[14][110] ),
    .B(_12859_),
    .S(_14132_),
    .Z(_01489_));
 MUX2_X1 _37386_ (.A(\core.keymem.key_mem[14][111] ),
    .B(_12017_),
    .S(_14132_),
    .Z(_01490_));
 MUX2_X1 _37387_ (.A(\core.keymem.key_mem[14][112] ),
    .B(_12031_),
    .S(_14132_),
    .Z(_01491_));
 MUX2_X1 _37388_ (.A(\core.keymem.key_mem[14][113] ),
    .B(_12868_),
    .S(_14132_),
    .Z(_01492_));
 MUX2_X1 _37389_ (.A(\core.keymem.key_mem[14][114] ),
    .B(_12869_),
    .S(_14132_),
    .Z(_01493_));
 MUX2_X1 _37390_ (.A(\core.keymem.key_mem[14][115] ),
    .B(_12059_),
    .S(_14132_),
    .Z(_01494_));
 BUF_X4 _37391_ (.A(_14124_),
    .Z(_14134_));
 MUX2_X1 _37392_ (.A(\core.keymem.key_mem[14][116] ),
    .B(_12077_),
    .S(_14134_),
    .Z(_01495_));
 MUX2_X1 _37393_ (.A(\core.keymem.key_mem[14][117] ),
    .B(_12877_),
    .S(_14134_),
    .Z(_01496_));
 MUX2_X1 _37394_ (.A(\core.keymem.key_mem[14][118] ),
    .B(_12882_),
    .S(_14134_),
    .Z(_01497_));
 MUX2_X1 _37395_ (.A(\core.keymem.key_mem[14][119] ),
    .B(_12096_),
    .S(_14134_),
    .Z(_01498_));
 NAND2_X1 _37396_ (.A1(\core.keymem.key_mem[14][11] ),
    .A2(_14128_),
    .ZN(_14135_));
 OAI21_X1 _37397_ (.A(_14135_),
    .B1(_14131_),
    .B2(_12895_),
    .ZN(_01499_));
 MUX2_X1 _37398_ (.A(\core.keymem.key_mem[14][120] ),
    .B(_12124_),
    .S(_14134_),
    .Z(_01500_));
 MUX2_X1 _37399_ (.A(\core.keymem.key_mem[14][121] ),
    .B(_12160_),
    .S(_14134_),
    .Z(_01501_));
 MUX2_X1 _37400_ (.A(\core.keymem.key_mem[14][122] ),
    .B(_12903_),
    .S(_14134_),
    .Z(_01502_));
 NAND2_X1 _37401_ (.A1(\core.keymem.key_mem[14][123] ),
    .A2(_14128_),
    .ZN(_14136_));
 OAI21_X1 _37402_ (.A(_14136_),
    .B1(_14131_),
    .B2(_12182_),
    .ZN(_01503_));
 NAND2_X1 _37403_ (.A1(\core.keymem.key_mem[14][124] ),
    .A2(_14128_),
    .ZN(_14137_));
 OAI21_X1 _37404_ (.A(_14137_),
    .B1(_14131_),
    .B2(_12926_),
    .ZN(_01504_));
 MUX2_X1 _37405_ (.A(\core.keymem.key_mem[14][125] ),
    .B(_12932_),
    .S(_14134_),
    .Z(_01505_));
 NAND2_X1 _37406_ (.A1(\core.keymem.key_mem[14][126] ),
    .A2(_14128_),
    .ZN(_14138_));
 OAI21_X1 _37407_ (.A(_14138_),
    .B1(_14131_),
    .B2(_12207_),
    .ZN(_01506_));
 MUX2_X1 _37408_ (.A(\core.keymem.key_mem[14][127] ),
    .B(_12945_),
    .S(_14134_),
    .Z(_01507_));
 MUX2_X1 _37409_ (.A(\core.keymem.key_mem[14][12] ),
    .B(_12958_),
    .S(_14134_),
    .Z(_01508_));
 BUF_X4 _37410_ (.A(_14123_),
    .Z(_14139_));
 MUX2_X1 _37411_ (.A(\core.keymem.key_mem[14][13] ),
    .B(_12974_),
    .S(_14139_),
    .Z(_01509_));
 NOR2_X1 _37412_ (.A1(\core.keymem.key_mem[14][14] ),
    .A2(_14125_),
    .ZN(_14140_));
 AOI21_X1 _37413_ (.A(_14140_),
    .B1(_14125_),
    .B2(_13007_),
    .ZN(_01510_));
 MUX2_X1 _37414_ (.A(\core.keymem.key_mem[14][15] ),
    .B(_13017_),
    .S(_14139_),
    .Z(_01511_));
 MUX2_X1 _37415_ (.A(\core.keymem.key_mem[14][16] ),
    .B(_13029_),
    .S(_14139_),
    .Z(_01512_));
 NAND2_X1 _37416_ (.A1(\core.keymem.key_mem[14][17] ),
    .A2(_14128_),
    .ZN(_14141_));
 OAI21_X1 _37417_ (.A(_14141_),
    .B1(_14131_),
    .B2(_13042_),
    .ZN(_01513_));
 MUX2_X1 _37418_ (.A(\core.keymem.key_mem[14][18] ),
    .B(_13094_),
    .S(_14139_),
    .Z(_01514_));
 BUF_X4 _37419_ (.A(_14127_),
    .Z(_14142_));
 NAND2_X1 _37420_ (.A1(\core.keymem.key_mem[14][19] ),
    .A2(_14142_),
    .ZN(_14143_));
 OAI21_X1 _37421_ (.A(_14143_),
    .B1(_14131_),
    .B2(_13109_),
    .ZN(_01515_));
 MUX2_X1 _37422_ (.A(\core.keymem.key_mem[14][1] ),
    .B(_13134_),
    .S(_14139_),
    .Z(_01516_));
 MUX2_X1 _37423_ (.A(\core.keymem.key_mem[14][20] ),
    .B(_13146_),
    .S(_14139_),
    .Z(_01517_));
 MUX2_X1 _37424_ (.A(\core.keymem.key_mem[14][21] ),
    .B(_13155_),
    .S(_14139_),
    .Z(_01518_));
 NOR2_X1 _37425_ (.A1(\core.keymem.key_mem[14][22] ),
    .A2(_14125_),
    .ZN(_14144_));
 AOI21_X1 _37426_ (.A(_14144_),
    .B1(_14125_),
    .B2(_13191_),
    .ZN(_01519_));
 MUX2_X1 _37427_ (.A(\core.keymem.key_mem[14][23] ),
    .B(_13196_),
    .S(_14139_),
    .Z(_01520_));
 NAND2_X1 _37428_ (.A1(\core.keymem.key_mem[14][24] ),
    .A2(_14142_),
    .ZN(_14145_));
 OAI21_X1 _37429_ (.A(_14145_),
    .B1(_14131_),
    .B2(_13212_),
    .ZN(_01521_));
 MUX2_X1 _37430_ (.A(\core.keymem.key_mem[14][25] ),
    .B(_13233_),
    .S(_14139_),
    .Z(_01522_));
 MUX2_X1 _37431_ (.A(\core.keymem.key_mem[14][26] ),
    .B(_13241_),
    .S(_14139_),
    .Z(_01523_));
 BUF_X4 _37432_ (.A(_14123_),
    .Z(_14146_));
 MUX2_X1 _37433_ (.A(\core.keymem.key_mem[14][27] ),
    .B(_13284_),
    .S(_14146_),
    .Z(_01524_));
 MUX2_X1 _37434_ (.A(\core.keymem.key_mem[14][28] ),
    .B(_13325_),
    .S(_14146_),
    .Z(_01525_));
 MUX2_X1 _37435_ (.A(\core.keymem.key_mem[14][29] ),
    .B(_13329_),
    .S(_14146_),
    .Z(_01526_));
 NAND2_X1 _37436_ (.A1(\core.keymem.key_mem[14][2] ),
    .A2(_14142_),
    .ZN(_14147_));
 OAI21_X1 _37437_ (.A(_14147_),
    .B1(_14131_),
    .B2(_13335_),
    .ZN(_01527_));
 MUX2_X1 _37438_ (.A(\core.keymem.key_mem[14][30] ),
    .B(_13379_),
    .S(_14146_),
    .Z(_01528_));
 MUX2_X1 _37439_ (.A(\core.keymem.key_mem[14][31] ),
    .B(_13395_),
    .S(_14146_),
    .Z(_01529_));
 MUX2_X1 _37440_ (.A(\core.keymem.key_mem[14][32] ),
    .B(_13396_),
    .S(_14146_),
    .Z(_01530_));
 MUX2_X1 _37441_ (.A(\core.keymem.key_mem[14][33] ),
    .B(_13402_),
    .S(_14146_),
    .Z(_01531_));
 MUX2_X1 _37442_ (.A(\core.keymem.key_mem[14][34] ),
    .B(_13403_),
    .S(_14146_),
    .Z(_01532_));
 MUX2_X1 _37443_ (.A(\core.keymem.key_mem[14][35] ),
    .B(_13405_),
    .S(_14146_),
    .Z(_01533_));
 NAND2_X1 _37444_ (.A1(\core.keymem.key_mem[14][36] ),
    .A2(_14142_),
    .ZN(_14148_));
 BUF_X4 _37445_ (.A(_14130_),
    .Z(_14149_));
 OAI21_X1 _37446_ (.A(_14148_),
    .B1(_14149_),
    .B2(_13407_),
    .ZN(_01534_));
 NAND2_X1 _37447_ (.A1(\core.keymem.key_mem[14][37] ),
    .A2(_14142_),
    .ZN(_14150_));
 OAI21_X1 _37448_ (.A(_14150_),
    .B1(_14149_),
    .B2(_12439_),
    .ZN(_01535_));
 MUX2_X1 _37449_ (.A(\core.keymem.key_mem[14][38] ),
    .B(_13410_),
    .S(_14146_),
    .Z(_01536_));
 NAND2_X1 _37450_ (.A1(\core.keymem.key_mem[14][39] ),
    .A2(_14142_),
    .ZN(_14151_));
 OAI21_X1 _37451_ (.A(_14151_),
    .B1(_14149_),
    .B2(_13435_),
    .ZN(_01537_));
 NAND2_X1 _37452_ (.A1(\core.keymem.key_mem[14][3] ),
    .A2(_14142_),
    .ZN(_14152_));
 OAI21_X1 _37453_ (.A(_14152_),
    .B1(_14149_),
    .B2(_13448_),
    .ZN(_01538_));
 NAND2_X1 _37454_ (.A1(\core.keymem.key_mem[14][40] ),
    .A2(_14142_),
    .ZN(_14153_));
 OAI21_X1 _37455_ (.A(_14153_),
    .B1(_14149_),
    .B2(_13457_),
    .ZN(_01539_));
 BUF_X4 _37456_ (.A(_14123_),
    .Z(_14154_));
 MUX2_X1 _37457_ (.A(\core.keymem.key_mem[14][41] ),
    .B(_13467_),
    .S(_14154_),
    .Z(_01540_));
 MUX2_X1 _37458_ (.A(\core.keymem.key_mem[14][42] ),
    .B(_13490_),
    .S(_14154_),
    .Z(_01541_));
 NAND2_X1 _37459_ (.A1(\core.keymem.key_mem[14][43] ),
    .A2(_14142_),
    .ZN(_14155_));
 OAI21_X1 _37460_ (.A(_14155_),
    .B1(_14149_),
    .B2(_13496_),
    .ZN(_01542_));
 MUX2_X1 _37461_ (.A(\core.keymem.key_mem[14][44] ),
    .B(_13497_),
    .S(_14154_),
    .Z(_01543_));
 NAND2_X1 _37462_ (.A1(\core.keymem.key_mem[14][45] ),
    .A2(_14142_),
    .ZN(_14156_));
 OAI21_X1 _37463_ (.A(_14156_),
    .B1(_14149_),
    .B2(_13510_),
    .ZN(_01544_));
 BUF_X4 _37464_ (.A(_14127_),
    .Z(_14157_));
 NAND2_X1 _37465_ (.A1(\core.keymem.key_mem[14][46] ),
    .A2(_14157_),
    .ZN(_14158_));
 OAI21_X1 _37466_ (.A(_14158_),
    .B1(_14149_),
    .B2(_13517_),
    .ZN(_01545_));
 NAND2_X1 _37467_ (.A1(\core.keymem.key_mem[14][47] ),
    .A2(_14157_),
    .ZN(_14159_));
 OAI21_X1 _37468_ (.A(_14159_),
    .B1(_14149_),
    .B2(_12520_),
    .ZN(_01546_));
 NAND2_X1 _37469_ (.A1(\core.keymem.key_mem[14][48] ),
    .A2(_14157_),
    .ZN(_14160_));
 OAI21_X1 _37470_ (.A(_14160_),
    .B1(_14149_),
    .B2(_12532_),
    .ZN(_01547_));
 NAND2_X1 _37471_ (.A1(\core.keymem.key_mem[14][49] ),
    .A2(_14157_),
    .ZN(_14161_));
 BUF_X4 _37472_ (.A(_14130_),
    .Z(_14162_));
 OAI21_X1 _37473_ (.A(_14161_),
    .B1(_14162_),
    .B2(_13529_),
    .ZN(_01548_));
 MUX2_X1 _37474_ (.A(\core.keymem.key_mem[14][4] ),
    .B(_13538_),
    .S(_14154_),
    .Z(_01549_));
 MUX2_X1 _37475_ (.A(\core.keymem.key_mem[14][50] ),
    .B(_13557_),
    .S(_14154_),
    .Z(_01550_));
 MUX2_X1 _37476_ (.A(\core.keymem.key_mem[14][51] ),
    .B(_13564_),
    .S(_14154_),
    .Z(_01551_));
 NAND2_X1 _37477_ (.A1(\core.keymem.key_mem[14][52] ),
    .A2(_14157_),
    .ZN(_14163_));
 OAI21_X1 _37478_ (.A(_14163_),
    .B1(_14162_),
    .B2(_12568_),
    .ZN(_01552_));
 NAND2_X1 _37479_ (.A1(\core.keymem.key_mem[14][53] ),
    .A2(_14157_),
    .ZN(_14164_));
 OAI21_X1 _37480_ (.A(_14164_),
    .B1(_14162_),
    .B2(_12584_),
    .ZN(_01553_));
 NAND2_X1 _37481_ (.A1(\core.keymem.key_mem[14][54] ),
    .A2(_14157_),
    .ZN(_14165_));
 OAI21_X1 _37482_ (.A(_14165_),
    .B1(_14162_),
    .B2(_13575_),
    .ZN(_01554_));
 MUX2_X1 _37483_ (.A(\core.keymem.key_mem[14][55] ),
    .B(_13581_),
    .S(_14154_),
    .Z(_01555_));
 MUX2_X1 _37484_ (.A(\core.keymem.key_mem[14][56] ),
    .B(_13589_),
    .S(_14154_),
    .Z(_01556_));
 MUX2_X1 _37485_ (.A(\core.keymem.key_mem[14][57] ),
    .B(_13604_),
    .S(_14154_),
    .Z(_01557_));
 MUX2_X1 _37486_ (.A(\core.keymem.key_mem[14][58] ),
    .B(_13611_),
    .S(_14154_),
    .Z(_01558_));
 BUF_X4 _37487_ (.A(_14123_),
    .Z(_14166_));
 MUX2_X1 _37488_ (.A(\core.keymem.key_mem[14][59] ),
    .B(_13616_),
    .S(_14166_),
    .Z(_01559_));
 MUX2_X1 _37489_ (.A(\core.keymem.key_mem[14][5] ),
    .B(_12606_),
    .S(_14166_),
    .Z(_01560_));
 MUX2_X1 _37490_ (.A(\core.keymem.key_mem[14][60] ),
    .B(_13622_),
    .S(_14166_),
    .Z(_01561_));
 MUX2_X1 _37491_ (.A(\core.keymem.key_mem[14][61] ),
    .B(_13632_),
    .S(_14166_),
    .Z(_01562_));
 MUX2_X1 _37492_ (.A(\core.keymem.key_mem[14][62] ),
    .B(_13637_),
    .S(_14166_),
    .Z(_01563_));
 MUX2_X1 _37493_ (.A(\core.keymem.key_mem[14][63] ),
    .B(_13659_),
    .S(_14166_),
    .Z(_01564_));
 MUX2_X1 _37494_ (.A(\core.keymem.key_mem[14][64] ),
    .B(_12622_),
    .S(_14166_),
    .Z(_01565_));
 NAND2_X1 _37495_ (.A1(\core.keymem.key_mem[14][65] ),
    .A2(_14157_),
    .ZN(_14167_));
 OAI21_X1 _37496_ (.A(_14167_),
    .B1(_14162_),
    .B2(_13673_),
    .ZN(_01566_));
 MUX2_X1 _37497_ (.A(\core.keymem.key_mem[14][66] ),
    .B(_13681_),
    .S(_14166_),
    .Z(_01567_));
 NAND2_X1 _37498_ (.A1(\core.keymem.key_mem[14][67] ),
    .A2(_14157_),
    .ZN(_14168_));
 OAI21_X1 _37499_ (.A(_14168_),
    .B1(_14162_),
    .B2(_13690_),
    .ZN(_01568_));
 NAND2_X1 _37500_ (.A1(\core.keymem.key_mem[14][68] ),
    .A2(_14157_),
    .ZN(_14169_));
 OAI21_X1 _37501_ (.A(_14169_),
    .B1(_14162_),
    .B2(_12635_),
    .ZN(_01569_));
 BUF_X4 _37502_ (.A(_14127_),
    .Z(_14170_));
 NAND2_X1 _37503_ (.A1(\core.keymem.key_mem[14][69] ),
    .A2(_14170_),
    .ZN(_14171_));
 OAI21_X1 _37504_ (.A(_14171_),
    .B1(_14162_),
    .B2(_13700_),
    .ZN(_01570_));
 MUX2_X1 _37505_ (.A(\core.keymem.key_mem[14][6] ),
    .B(_13711_),
    .S(_14166_),
    .Z(_01571_));
 MUX2_X1 _37506_ (.A(\core.keymem.key_mem[14][70] ),
    .B(_13713_),
    .S(_14166_),
    .Z(_01572_));
 NAND2_X1 _37507_ (.A1(\core.keymem.key_mem[14][71] ),
    .A2(_14170_),
    .ZN(_14172_));
 OAI21_X1 _37508_ (.A(_14172_),
    .B1(_14162_),
    .B2(_12659_),
    .ZN(_01573_));
 NAND2_X1 _37509_ (.A1(\core.keymem.key_mem[14][72] ),
    .A2(_14170_),
    .ZN(_14173_));
 OAI21_X1 _37510_ (.A(_14173_),
    .B1(_14162_),
    .B2(_13716_),
    .ZN(_01574_));
 NAND2_X1 _37511_ (.A1(\core.keymem.key_mem[14][73] ),
    .A2(_14170_),
    .ZN(_14174_));
 BUF_X4 _37512_ (.A(_14130_),
    .Z(_14175_));
 OAI21_X1 _37513_ (.A(_14174_),
    .B1(_14175_),
    .B2(_12688_),
    .ZN(_01575_));
 NAND2_X1 _37514_ (.A1(\core.keymem.key_mem[14][74] ),
    .A2(_14170_),
    .ZN(_14176_));
 OAI21_X1 _37515_ (.A(_14176_),
    .B1(_14175_),
    .B2(_13726_),
    .ZN(_01576_));
 NAND2_X1 _37516_ (.A1(\core.keymem.key_mem[14][75] ),
    .A2(_14170_),
    .ZN(_14177_));
 OAI21_X1 _37517_ (.A(_14177_),
    .B1(_14175_),
    .B2(_13733_),
    .ZN(_01577_));
 BUF_X4 _37518_ (.A(_14123_),
    .Z(_14178_));
 MUX2_X1 _37519_ (.A(\core.keymem.key_mem[14][76] ),
    .B(_13741_),
    .S(_14178_),
    .Z(_01578_));
 MUX2_X1 _37520_ (.A(\core.keymem.key_mem[14][77] ),
    .B(_13751_),
    .S(_14178_),
    .Z(_01579_));
 NAND2_X1 _37521_ (.A1(\core.keymem.key_mem[14][78] ),
    .A2(_14170_),
    .ZN(_14179_));
 OAI21_X1 _37522_ (.A(_14179_),
    .B1(_14175_),
    .B2(_12708_),
    .ZN(_01580_));
 MUX2_X1 _37523_ (.A(\core.keymem.key_mem[14][79] ),
    .B(_13758_),
    .S(_14178_),
    .Z(_01581_));
 NAND2_X1 _37524_ (.A1(\core.keymem.key_mem[14][7] ),
    .A2(_14170_),
    .ZN(_14180_));
 OAI21_X1 _37525_ (.A(_14180_),
    .B1(_14175_),
    .B2(_13767_),
    .ZN(_01582_));
 MUX2_X1 _37526_ (.A(\core.keymem.key_mem[14][80] ),
    .B(_13769_),
    .S(_14178_),
    .Z(_01583_));
 NAND2_X1 _37527_ (.A1(\core.keymem.key_mem[14][81] ),
    .A2(_14170_),
    .ZN(_14181_));
 OAI21_X1 _37528_ (.A(_14181_),
    .B1(_14175_),
    .B2(_13775_),
    .ZN(_01584_));
 NAND2_X1 _37529_ (.A1(\core.keymem.key_mem[14][82] ),
    .A2(_14170_),
    .ZN(_14182_));
 OAI21_X1 _37530_ (.A(_14182_),
    .B1(_14175_),
    .B2(_13783_),
    .ZN(_01585_));
 NAND2_X1 _37531_ (.A1(\core.keymem.key_mem[14][83] ),
    .A2(_14130_),
    .ZN(_14183_));
 OAI21_X1 _37532_ (.A(_14183_),
    .B1(_14175_),
    .B2(_13791_),
    .ZN(_01586_));
 NAND2_X1 _37533_ (.A1(\core.keymem.key_mem[14][84] ),
    .A2(_14130_),
    .ZN(_14184_));
 OAI21_X1 _37534_ (.A(_14184_),
    .B1(_14175_),
    .B2(_12725_),
    .ZN(_01587_));
 MUX2_X1 _37535_ (.A(\core.keymem.key_mem[14][85] ),
    .B(_13798_),
    .S(_14178_),
    .Z(_01588_));
 MUX2_X1 _37536_ (.A(\core.keymem.key_mem[14][86] ),
    .B(_12741_),
    .S(_14178_),
    .Z(_01589_));
 MUX2_X1 _37537_ (.A(\core.keymem.key_mem[14][87] ),
    .B(_13804_),
    .S(_14178_),
    .Z(_01590_));
 MUX2_X1 _37538_ (.A(\core.keymem.key_mem[14][88] ),
    .B(_13810_),
    .S(_14178_),
    .Z(_01591_));
 MUX2_X1 _37539_ (.A(\core.keymem.key_mem[14][89] ),
    .B(_13818_),
    .S(_14178_),
    .Z(_01592_));
 MUX2_X1 _37540_ (.A(\core.keymem.key_mem[14][8] ),
    .B(_13854_),
    .S(_14178_),
    .Z(_01593_));
 MUX2_X1 _37541_ (.A(\core.keymem.key_mem[14][90] ),
    .B(_13860_),
    .S(_14124_),
    .Z(_01594_));
 NAND2_X1 _37542_ (.A1(\core.keymem.key_mem[14][91] ),
    .A2(_14130_),
    .ZN(_14185_));
 OAI21_X1 _37543_ (.A(_14185_),
    .B1(_14175_),
    .B2(_13870_),
    .ZN(_01595_));
 NAND2_X1 _37544_ (.A1(\core.keymem.key_mem[14][92] ),
    .A2(_14130_),
    .ZN(_14186_));
 OAI21_X1 _37545_ (.A(_14186_),
    .B1(_14128_),
    .B2(_13880_),
    .ZN(_01596_));
 MUX2_X1 _37546_ (.A(\core.keymem.key_mem[14][93] ),
    .B(_13889_),
    .S(_14124_),
    .Z(_01597_));
 MUX2_X1 _37547_ (.A(\core.keymem.key_mem[14][94] ),
    .B(_13896_),
    .S(_14124_),
    .Z(_01598_));
 MUX2_X1 _37548_ (.A(\core.keymem.key_mem[14][95] ),
    .B(_13903_),
    .S(_14124_),
    .Z(_01599_));
 MUX2_X1 _37549_ (.A(\core.keymem.key_mem[14][96] ),
    .B(_13907_),
    .S(_14124_),
    .Z(_01600_));
 NAND2_X1 _37550_ (.A1(\core.keymem.key_mem[14][97] ),
    .A2(_14130_),
    .ZN(_14187_));
 OAI21_X1 _37551_ (.A(_14187_),
    .B1(_14128_),
    .B2(_12777_),
    .ZN(_01601_));
 NAND2_X1 _37552_ (.A1(\core.keymem.key_mem[14][98] ),
    .A2(_14130_),
    .ZN(_14188_));
 OAI21_X1 _37553_ (.A(_14188_),
    .B1(_14128_),
    .B2(_13910_),
    .ZN(_01602_));
 MUX2_X1 _37554_ (.A(\core.keymem.key_mem[14][99] ),
    .B(_12800_),
    .S(_14124_),
    .Z(_01603_));
 MUX2_X1 _37555_ (.A(\core.keymem.key_mem[14][9] ),
    .B(_13919_),
    .S(_14124_),
    .Z(_01604_));
 NAND2_X4 _37556_ (.A1(_11792_),
    .A2(_11997_),
    .ZN(_14189_));
 BUF_X8 _37557_ (.A(_14189_),
    .Z(_14190_));
 BUF_X4 _37558_ (.A(_14190_),
    .Z(_14191_));
 NOR2_X4 _37559_ (.A1(_11804_),
    .A2(_14189_),
    .ZN(_14192_));
 BUF_X4 _37560_ (.A(_14192_),
    .Z(_14193_));
 AOI22_X1 _37561_ (.A1(\core.keymem.key_mem[1][0] ),
    .A2(_14191_),
    .B1(_14193_),
    .B2(_11844_),
    .ZN(_14194_));
 INV_X1 _37562_ (.A(_14194_),
    .ZN(_01605_));
 NOR2_X4 _37563_ (.A1(_16224_),
    .A2(_12365_),
    .ZN(_14195_));
 BUF_X4 _37564_ (.A(_14195_),
    .Z(_14196_));
 MUX2_X1 _37565_ (.A(\core.keymem.key_mem[1][100] ),
    .B(_11873_),
    .S(_14196_),
    .Z(_01606_));
 INV_X1 _37566_ (.A(\core.keymem.key_mem[1][101] ),
    .ZN(_14197_));
 BUF_X4 _37567_ (.A(_14195_),
    .Z(_14198_));
 BUF_X4 _37568_ (.A(_14198_),
    .Z(_14199_));
 NAND2_X4 _37569_ (.A1(_16229_),
    .A2(_14195_),
    .ZN(_14200_));
 BUF_X8 _37570_ (.A(_12871_),
    .Z(_14201_));
 OAI21_X4 _37571_ (.A(_12812_),
    .B1(_14201_),
    .B2(_11879_),
    .ZN(_14202_));
 OAI22_X1 _37572_ (.A1(_14197_),
    .A2(_14199_),
    .B1(_14200_),
    .B2(_14202_),
    .ZN(_01607_));
 AOI22_X1 _37573_ (.A1(\core.keymem.key_mem[1][102] ),
    .A2(_14191_),
    .B1(_14193_),
    .B2(_11906_),
    .ZN(_14203_));
 INV_X1 _37574_ (.A(_14203_),
    .ZN(_01608_));
 MUX2_X1 _37575_ (.A(\core.keymem.key_mem[1][103] ),
    .B(_11929_),
    .S(_14196_),
    .Z(_01609_));
 INV_X1 _37576_ (.A(\core.keymem.key_mem[1][104] ),
    .ZN(_14204_));
 BUF_X8 _37577_ (.A(_12779_),
    .Z(_14205_));
 BUF_X4 _37578_ (.A(_14205_),
    .Z(_14206_));
 NAND2_X1 _37579_ (.A1(_00133_),
    .A2(_14206_),
    .ZN(_14207_));
 NAND3_X1 _37580_ (.A1(_16285_),
    .A2(_14196_),
    .A3(_14207_),
    .ZN(_14208_));
 OAI22_X1 _37581_ (.A1(_14204_),
    .A2(_14199_),
    .B1(_14208_),
    .B2(_12821_),
    .ZN(_01610_));
 BUF_X4 _37582_ (.A(_14190_),
    .Z(_14209_));
 NAND2_X1 _37583_ (.A1(\core.keymem.key_mem[1][105] ),
    .A2(_14209_),
    .ZN(_14210_));
 BUF_X8 _37584_ (.A(_11952_),
    .Z(_14211_));
 BUF_X8 _37585_ (.A(_12193_),
    .Z(_14212_));
 NAND2_X1 _37586_ (.A1(_00134_),
    .A2(_14212_),
    .ZN(_14213_));
 NAND3_X1 _37587_ (.A1(_14211_),
    .A2(_12830_),
    .A3(_14213_),
    .ZN(_14214_));
 OAI21_X1 _37588_ (.A(_14210_),
    .B1(_14214_),
    .B2(_14209_),
    .ZN(_01611_));
 NAND2_X1 _37589_ (.A1(\core.keymem.key_mem[1][106] ),
    .A2(_14209_),
    .ZN(_14215_));
 BUF_X4 _37590_ (.A(_14200_),
    .Z(_14216_));
 OAI21_X1 _37591_ (.A(_14215_),
    .B1(_14216_),
    .B2(_11951_),
    .ZN(_01612_));
 MUX2_X1 _37592_ (.A(\core.keymem.key_mem[1][107] ),
    .B(_11967_),
    .S(_14196_),
    .Z(_01613_));
 MUX2_X1 _37593_ (.A(\core.keymem.key_mem[1][108] ),
    .B(_11981_),
    .S(_14196_),
    .Z(_01614_));
 BUF_X4 _37594_ (.A(_14192_),
    .Z(_14217_));
 NAND2_X1 _37595_ (.A1(_00141_),
    .A2(_14212_),
    .ZN(_14218_));
 NAND3_X1 _37596_ (.A1(_12842_),
    .A2(_14217_),
    .A3(_14218_),
    .ZN(_14219_));
 BUF_X4 _37597_ (.A(_14198_),
    .Z(_14220_));
 INV_X1 _37598_ (.A(\core.keymem.key_mem[1][109] ),
    .ZN(_14221_));
 OAI21_X1 _37599_ (.A(_14219_),
    .B1(_14220_),
    .B2(_14221_),
    .ZN(_01615_));
 BUF_X4 _37600_ (.A(_13720_),
    .Z(_14222_));
 NOR4_X1 _37601_ (.A1(_11805_),
    .A2(_11983_),
    .A3(_14222_),
    .A4(_14189_),
    .ZN(_14223_));
 BUF_X8 _37602_ (.A(_14190_),
    .Z(_14224_));
 AOI21_X1 _37603_ (.A(_14223_),
    .B1(_14224_),
    .B2(\core.keymem.key_mem[1][10] ),
    .ZN(_14225_));
 BUF_X4 _37604_ (.A(_12186_),
    .Z(_14226_));
 BUF_X8 _37605_ (.A(_14198_),
    .Z(_14227_));
 NAND3_X1 _37606_ (.A1(_16285_),
    .A2(_14226_),
    .A3(_14227_),
    .ZN(_14228_));
 NAND2_X1 _37607_ (.A1(_06678_),
    .A2(_12851_),
    .ZN(_14229_));
 OAI22_X2 _37608_ (.A1(_06680_),
    .A2(_12856_),
    .B1(_14229_),
    .B2(_12850_),
    .ZN(_14230_));
 OAI21_X1 _37609_ (.A(_14225_),
    .B1(_14228_),
    .B2(_14230_),
    .ZN(_01616_));
 NAND2_X1 _37610_ (.A1(\core.keymem.key_mem[1][110] ),
    .A2(_14209_),
    .ZN(_14231_));
 BUF_X4 _37611_ (.A(_14190_),
    .Z(_14232_));
 OAI21_X1 _37612_ (.A(_14231_),
    .B1(_14232_),
    .B2(_12004_),
    .ZN(_01617_));
 MUX2_X1 _37613_ (.A(\core.keymem.key_mem[1][111] ),
    .B(_12017_),
    .S(_14196_),
    .Z(_01618_));
 AOI22_X1 _37614_ (.A1(\core.keymem.key_mem[1][112] ),
    .A2(_14224_),
    .B1(_14193_),
    .B2(_12031_),
    .ZN(_14233_));
 INV_X1 _37615_ (.A(_14233_),
    .ZN(_01619_));
 NAND2_X1 _37616_ (.A1(\core.keymem.key_mem[1][113] ),
    .A2(_14209_),
    .ZN(_14234_));
 BUF_X4 _37617_ (.A(_14198_),
    .Z(_14235_));
 NAND2_X1 _37618_ (.A1(_00146_),
    .A2(_14206_),
    .ZN(_14236_));
 NAND3_X1 _37619_ (.A1(_14211_),
    .A2(_14235_),
    .A3(_14236_),
    .ZN(_14237_));
 BUF_X8 _37620_ (.A(_14212_),
    .Z(_14238_));
 NOR2_X1 _37621_ (.A1(_14238_),
    .A2(_12866_),
    .ZN(_14239_));
 OAI21_X1 _37622_ (.A(_14234_),
    .B1(_14237_),
    .B2(_14239_),
    .ZN(_01620_));
 NAND2_X1 _37623_ (.A1(\core.keymem.key_mem[1][114] ),
    .A2(_14209_),
    .ZN(_14240_));
 OAI21_X1 _37624_ (.A(_14240_),
    .B1(_14232_),
    .B2(_12049_),
    .ZN(_01621_));
 MUX2_X1 _37625_ (.A(\core.keymem.key_mem[1][115] ),
    .B(_12059_),
    .S(_14196_),
    .Z(_01622_));
 MUX2_X1 _37626_ (.A(\core.keymem.key_mem[1][116] ),
    .B(_12077_),
    .S(_14196_),
    .Z(_01623_));
 INV_X1 _37627_ (.A(\core.keymem.key_mem[1][117] ),
    .ZN(_14241_));
 BUF_X4 _37628_ (.A(_12860_),
    .Z(_14242_));
 NAND2_X2 _37629_ (.A1(_00153_),
    .A2(_14242_),
    .ZN(_14243_));
 NAND3_X1 _37630_ (.A1(_16285_),
    .A2(_14196_),
    .A3(_14243_),
    .ZN(_14244_));
 BUF_X4 _37631_ (.A(_13875_),
    .Z(_14245_));
 AND3_X2 _37632_ (.A1(_14245_),
    .A2(_12874_),
    .A3(_12875_),
    .ZN(_14246_));
 OAI22_X1 _37633_ (.A1(_14241_),
    .A2(_14199_),
    .B1(_14244_),
    .B2(_14246_),
    .ZN(_01624_));
 NAND2_X1 _37634_ (.A1(\core.keymem.key_mem[1][118] ),
    .A2(_14209_),
    .ZN(_14247_));
 BUF_X8 _37635_ (.A(_14222_),
    .Z(_14248_));
 OAI21_X4 _37636_ (.A(_12881_),
    .B1(_14248_),
    .B2(_12079_),
    .ZN(_14249_));
 BUF_X4 _37637_ (.A(_14200_),
    .Z(_14250_));
 OAI21_X1 _37638_ (.A(_14247_),
    .B1(_14249_),
    .B2(_14250_),
    .ZN(_01625_));
 MUX2_X1 _37639_ (.A(\core.keymem.key_mem[1][119] ),
    .B(_12096_),
    .S(_14196_),
    .Z(_01626_));
 BUF_X4 _37640_ (.A(_14190_),
    .Z(_14251_));
 NAND2_X1 _37641_ (.A1(\core.keymem.key_mem[1][11] ),
    .A2(_14251_),
    .ZN(_14252_));
 NOR2_X2 _37642_ (.A1(_00406_),
    .A2(_14222_),
    .ZN(_14253_));
 MUX2_X1 _37643_ (.A(_12888_),
    .B(_12893_),
    .S(_13132_),
    .Z(_14254_));
 AOI21_X4 _37644_ (.A(_14253_),
    .B1(_14254_),
    .B2(_14248_),
    .ZN(_14255_));
 OAI21_X1 _37645_ (.A(_14252_),
    .B1(_14255_),
    .B2(_14250_),
    .ZN(_01627_));
 AOI22_X1 _37646_ (.A1(\core.keymem.key_mem[1][120] ),
    .A2(_14224_),
    .B1(_14193_),
    .B2(_12124_),
    .ZN(_14256_));
 INV_X1 _37647_ (.A(_14256_),
    .ZN(_01628_));
 NAND2_X1 _37648_ (.A1(_12160_),
    .A2(_14217_),
    .ZN(_14257_));
 INV_X1 _37649_ (.A(\core.keymem.key_mem[1][121] ),
    .ZN(_14258_));
 OAI21_X1 _37650_ (.A(_14257_),
    .B1(_14220_),
    .B2(_14258_),
    .ZN(_01629_));
 AOI22_X1 _37651_ (.A1(\core.keymem.key_mem[1][122] ),
    .A2(_14224_),
    .B1(_14193_),
    .B2(_12903_),
    .ZN(_14259_));
 INV_X1 _37652_ (.A(_14259_),
    .ZN(_01630_));
 NAND2_X1 _37653_ (.A1(\core.keymem.key_mem[1][123] ),
    .A2(_14251_),
    .ZN(_14260_));
 OAI21_X1 _37654_ (.A(_14260_),
    .B1(_14216_),
    .B2(_12182_),
    .ZN(_01631_));
 NOR2_X1 _37655_ (.A1(_11930_),
    .A2(_12925_),
    .ZN(_14261_));
 BUF_X8 _37656_ (.A(_14195_),
    .Z(_14262_));
 MUX2_X1 _37657_ (.A(\core.keymem.key_mem[1][124] ),
    .B(_14261_),
    .S(_14262_),
    .Z(_01632_));
 NAND2_X1 _37658_ (.A1(\core.keymem.key_mem[1][125] ),
    .A2(_14251_),
    .ZN(_14263_));
 BUF_X8 _37659_ (.A(_14205_),
    .Z(_14264_));
 BUF_X4 _37660_ (.A(_12028_),
    .Z(_14265_));
 AOI22_X2 _37661_ (.A1(_12189_),
    .A2(_14264_),
    .B1(_14265_),
    .B2(_12930_),
    .ZN(_14266_));
 BUF_X4 _37662_ (.A(_12844_),
    .Z(_14267_));
 AND2_X1 _37663_ (.A1(_14267_),
    .A2(_12306_),
    .ZN(_14268_));
 OAI21_X2 _37664_ (.A(_14266_),
    .B1(_12928_),
    .B2(_14268_),
    .ZN(_14269_));
 OAI21_X1 _37665_ (.A(_14263_),
    .B1(_14216_),
    .B2(_14269_),
    .ZN(_01633_));
 NAND2_X1 _37666_ (.A1(\core.keymem.key_mem[1][126] ),
    .A2(_14251_),
    .ZN(_14270_));
 OAI21_X1 _37667_ (.A(_14270_),
    .B1(_14216_),
    .B2(_12207_),
    .ZN(_01634_));
 AOI22_X1 _37668_ (.A1(\core.keymem.key_mem[1][127] ),
    .A2(_14224_),
    .B1(_14193_),
    .B2(_12945_),
    .ZN(_14271_));
 INV_X1 _37669_ (.A(_14271_),
    .ZN(_01635_));
 NAND2_X1 _37670_ (.A1(\core.keymem.key_mem[1][12] ),
    .A2(_14251_),
    .ZN(_14272_));
 OR2_X1 _37671_ (.A1(_12947_),
    .A2(_12948_),
    .ZN(_14273_));
 BUF_X4 _37672_ (.A(_12156_),
    .Z(_14274_));
 NOR2_X1 _37673_ (.A1(_14274_),
    .A2(_12950_),
    .ZN(_14275_));
 NOR2_X1 _37674_ (.A1(_14242_),
    .A2(_14275_),
    .ZN(_14276_));
 BUF_X4 _37675_ (.A(_12345_),
    .Z(_14277_));
 BUF_X4 _37676_ (.A(_14277_),
    .Z(_14278_));
 XOR2_X2 _37677_ (.A(_11974_),
    .B(_12954_),
    .Z(_14279_));
 OAI21_X2 _37678_ (.A(_06679_),
    .B1(_14278_),
    .B2(_14279_),
    .ZN(_14280_));
 AOI21_X4 _37679_ (.A(_14273_),
    .B1(_14276_),
    .B2(_14280_),
    .ZN(_14281_));
 OAI21_X1 _37680_ (.A(_14272_),
    .B1(_14281_),
    .B2(_14250_),
    .ZN(_01636_));
 BUF_X4 _37681_ (.A(_11842_),
    .Z(_14282_));
 NAND2_X2 _37682_ (.A1(_12213_),
    .A2(_14282_),
    .ZN(_14283_));
 NOR3_X1 _37683_ (.A1(_12183_),
    .A2(_14189_),
    .A3(_14283_),
    .ZN(_14284_));
 AOI21_X1 _37684_ (.A(_14284_),
    .B1(_14224_),
    .B2(\core.keymem.key_mem[1][13] ),
    .ZN(_14285_));
 INV_X1 _37685_ (.A(_12967_),
    .ZN(_14286_));
 INV_X1 _37686_ (.A(\core.keymem.prev_key1_reg[13] ),
    .ZN(_14287_));
 XNOR2_X1 _37687_ (.A(_14287_),
    .B(_12969_),
    .ZN(_14288_));
 BUF_X4 _37688_ (.A(_14274_),
    .Z(_14289_));
 OAI21_X2 _37689_ (.A(_14286_),
    .B1(_14288_),
    .B2(_14289_),
    .ZN(_14290_));
 OAI21_X1 _37690_ (.A(_14285_),
    .B1(_14228_),
    .B2(_14290_),
    .ZN(_01637_));
 NAND2_X1 _37691_ (.A1(\core.keymem.key_mem[1][14] ),
    .A2(_14251_),
    .ZN(_14291_));
 NOR2_X1 _37692_ (.A1(_06680_),
    .A2(_13004_),
    .ZN(_14292_));
 BUF_X4 _37693_ (.A(_12972_),
    .Z(_14293_));
 INV_X1 _37694_ (.A(_12978_),
    .ZN(_14294_));
 NAND2_X1 _37695_ (.A1(_14294_),
    .A2(_11992_),
    .ZN(_14295_));
 NAND2_X1 _37696_ (.A1(_12979_),
    .A2(_12698_),
    .ZN(_14296_));
 OAI22_X1 _37697_ (.A1(_11992_),
    .A2(_12981_),
    .B1(_14295_),
    .B2(_14296_),
    .ZN(_14297_));
 NAND3_X1 _37698_ (.A1(_12149_),
    .A2(net11),
    .A3(_14297_),
    .ZN(_14298_));
 NOR2_X1 _37699_ (.A1(_11841_),
    .A2(_12977_),
    .ZN(_14299_));
 AOI21_X1 _37700_ (.A(_14293_),
    .B1(_14298_),
    .B2(_14299_),
    .ZN(_14300_));
 NOR2_X2 _37701_ (.A1(_14292_),
    .A2(_14300_),
    .ZN(_14301_));
 NAND2_X2 _37702_ (.A1(_00409_),
    .A2(_14282_),
    .ZN(_14302_));
 NAND3_X1 _37703_ (.A1(_11986_),
    .A2(_14227_),
    .A3(_14302_),
    .ZN(_14303_));
 OAI21_X1 _37704_ (.A(_14291_),
    .B1(_14301_),
    .B2(_14303_),
    .ZN(_01638_));
 BUF_X4 _37705_ (.A(_11800_),
    .Z(_14304_));
 NAND2_X2 _37706_ (.A1(_12217_),
    .A2(_14304_),
    .ZN(_14305_));
 AOI21_X4 _37707_ (.A(_13015_),
    .B1(_14305_),
    .B2(_13012_),
    .ZN(_14306_));
 MUX2_X1 _37708_ (.A(\core.keymem.key_mem[1][15] ),
    .B(_14306_),
    .S(_14262_),
    .Z(_01639_));
 NAND2_X2 _37709_ (.A1(_00411_),
    .A2(_14212_),
    .ZN(_14307_));
 NAND4_X1 _37710_ (.A1(_12751_),
    .A2(_13029_),
    .A3(_14227_),
    .A4(_14307_),
    .ZN(_14308_));
 INV_X1 _37711_ (.A(\core.keymem.key_mem[1][16] ),
    .ZN(_14309_));
 OAI21_X1 _37712_ (.A(_14308_),
    .B1(_14220_),
    .B2(_14309_),
    .ZN(_01640_));
 NAND2_X1 _37713_ (.A1(\core.keymem.key_mem[1][17] ),
    .A2(_14251_),
    .ZN(_14310_));
 NAND2_X1 _37714_ (.A1(_12301_),
    .A2(_13036_),
    .ZN(_14311_));
 OAI22_X1 _37715_ (.A1(_14274_),
    .A2(_13040_),
    .B1(_14311_),
    .B2(_13035_),
    .ZN(_14312_));
 BUF_X4 _37716_ (.A(_12834_),
    .Z(_14313_));
 MUX2_X2 _37717_ (.A(_00434_),
    .B(_14312_),
    .S(_14313_),
    .Z(_14314_));
 BUF_X4 _37718_ (.A(_14200_),
    .Z(_14315_));
 OAI21_X1 _37719_ (.A(_14310_),
    .B1(_14314_),
    .B2(_14315_),
    .ZN(_01641_));
 NAND2_X2 _37720_ (.A1(_00435_),
    .A2(_11800_),
    .ZN(_14316_));
 NAND4_X1 _37721_ (.A1(_14211_),
    .A2(_13094_),
    .A3(_14227_),
    .A4(_14316_),
    .ZN(_14317_));
 INV_X1 _37722_ (.A(\core.keymem.key_mem[1][18] ),
    .ZN(_14318_));
 OAI21_X1 _37723_ (.A(_14317_),
    .B1(_14220_),
    .B2(_14318_),
    .ZN(_01642_));
 NAND2_X1 _37724_ (.A1(\core.keymem.key_mem[1][19] ),
    .A2(_14251_),
    .ZN(_14319_));
 AOI21_X1 _37725_ (.A(_12292_),
    .B1(\core.key[19] ),
    .B2(_13415_),
    .ZN(_14320_));
 OAI21_X2 _37726_ (.A(_14320_),
    .B1(_13106_),
    .B2(_14277_),
    .ZN(_14321_));
 AOI22_X4 _37727_ (.A1(_12224_),
    .A2(_14238_),
    .B1(_13103_),
    .B2(_14321_),
    .ZN(_14322_));
 OAI21_X1 _37728_ (.A(_14319_),
    .B1(_14322_),
    .B2(_14315_),
    .ZN(_01643_));
 OAI22_X2 _37729_ (.A1(_12227_),
    .A2(_12347_),
    .B1(_12302_),
    .B2(\core.key[1] ),
    .ZN(_14323_));
 AOI221_X2 _37730_ (.A(_13115_),
    .B1(_14323_),
    .B2(_12951_),
    .C1(_12311_),
    .C2(_13121_),
    .ZN(_14324_));
 MUX2_X1 _37731_ (.A(\core.keymem.key_mem[1][1] ),
    .B(_14324_),
    .S(_14262_),
    .Z(_01644_));
 NAND2_X2 _37732_ (.A1(_12231_),
    .A2(_14304_),
    .ZN(_14325_));
 AOI21_X4 _37733_ (.A(_13144_),
    .B1(_14325_),
    .B2(_13141_),
    .ZN(_14326_));
 MUX2_X1 _37734_ (.A(\core.keymem.key_mem[1][20] ),
    .B(_14326_),
    .S(_14262_),
    .Z(_01645_));
 AOI21_X1 _37735_ (.A(_11846_),
    .B1(\core.key[21] ),
    .B2(_11892_),
    .ZN(_14327_));
 AOI221_X2 _37736_ (.A(_12680_),
    .B1(_13150_),
    .B2(_14327_),
    .C1(_13153_),
    .C2(_12971_),
    .ZN(_14328_));
 NOR2_X2 _37737_ (.A1(_00438_),
    .A2(_12185_),
    .ZN(_14329_));
 OAI21_X1 _37738_ (.A(_14217_),
    .B1(_14328_),
    .B2(_14329_),
    .ZN(_14330_));
 INV_X1 _37739_ (.A(\core.keymem.key_mem[1][21] ),
    .ZN(_14331_));
 OAI21_X1 _37740_ (.A(_14330_),
    .B1(_14220_),
    .B2(_14331_),
    .ZN(_01646_));
 NAND2_X4 _37741_ (.A1(_12235_),
    .A2(_14304_),
    .ZN(_14332_));
 AOI21_X1 _37742_ (.A(_12183_),
    .B1(_13190_),
    .B2(_14332_),
    .ZN(_14333_));
 MUX2_X1 _37743_ (.A(\core.keymem.key_mem[1][22] ),
    .B(_14333_),
    .S(_14262_),
    .Z(_01647_));
 NAND2_X1 _37744_ (.A1(\core.keymem.key_mem[1][23] ),
    .A2(_14251_),
    .ZN(_14334_));
 OAI21_X1 _37745_ (.A(_14334_),
    .B1(_14216_),
    .B2(_12272_),
    .ZN(_01648_));
 NOR2_X2 _37746_ (.A1(_11952_),
    .A2(_14189_),
    .ZN(_14335_));
 NOR4_X2 _37747_ (.A1(_13203_),
    .A2(_13209_),
    .A3(_13210_),
    .A4(_14189_),
    .ZN(_14336_));
 NOR2_X1 _37748_ (.A1(\core.keymem.key_mem[1][24] ),
    .A2(_14198_),
    .ZN(_14337_));
 NOR3_X1 _37749_ (.A1(_14335_),
    .A2(_14336_),
    .A3(_14337_),
    .ZN(_01649_));
 NAND2_X1 _37750_ (.A1(_00020_),
    .A2(_14212_),
    .ZN(_14338_));
 NAND3_X1 _37751_ (.A1(_13233_),
    .A2(_14217_),
    .A3(_14338_),
    .ZN(_14339_));
 INV_X1 _37752_ (.A(\core.keymem.key_mem[1][25] ),
    .ZN(_14340_));
 OAI21_X1 _37753_ (.A(_14339_),
    .B1(_14220_),
    .B2(_14340_),
    .ZN(_01650_));
 NAND3_X1 _37754_ (.A1(_12751_),
    .A2(_13241_),
    .A3(_14235_),
    .ZN(_14341_));
 INV_X1 _37755_ (.A(\core.keymem.key_mem[1][26] ),
    .ZN(_14342_));
 OAI21_X1 _37756_ (.A(_14341_),
    .B1(_14220_),
    .B2(_14342_),
    .ZN(_01651_));
 OAI21_X1 _37757_ (.A(_14217_),
    .B1(_13282_),
    .B2(_13276_),
    .ZN(_14343_));
 OAI21_X1 _37758_ (.A(_14343_),
    .B1(_14220_),
    .B2(_03322_),
    .ZN(_01652_));
 AOI21_X1 _37759_ (.A(_12183_),
    .B1(_13315_),
    .B2(_13323_),
    .ZN(_14344_));
 MUX2_X1 _37760_ (.A(\core.keymem.key_mem[1][28] ),
    .B(_14344_),
    .S(_14262_),
    .Z(_01653_));
 NAND2_X1 _37761_ (.A1(\core.keymem.key_mem[1][29] ),
    .A2(_14251_),
    .ZN(_14345_));
 OAI21_X1 _37762_ (.A(_14345_),
    .B1(_14216_),
    .B2(_12312_),
    .ZN(_01654_));
 INV_X1 _37763_ (.A(\core.keymem.key_mem[1][2] ),
    .ZN(_14346_));
 OAI22_X1 _37764_ (.A1(_14346_),
    .A2(_14199_),
    .B1(_14200_),
    .B2(_12337_),
    .ZN(_01655_));
 OAI21_X1 _37765_ (.A(_14217_),
    .B1(_13375_),
    .B2(_13341_),
    .ZN(_14347_));
 INV_X1 _37766_ (.A(\core.keymem.key_mem[1][30] ),
    .ZN(_14348_));
 OAI21_X1 _37767_ (.A(_14347_),
    .B1(_14220_),
    .B2(_14348_),
    .ZN(_01656_));
 BUF_X4 _37768_ (.A(_14190_),
    .Z(_14349_));
 NAND2_X1 _37769_ (.A1(\core.keymem.key_mem[1][31] ),
    .A2(_14349_),
    .ZN(_14350_));
 OAI21_X1 _37770_ (.A(_11986_),
    .B1(_13386_),
    .B2(_13393_),
    .ZN(_14351_));
 OAI21_X1 _37771_ (.A(_14350_),
    .B1(_14351_),
    .B2(_14209_),
    .ZN(_01657_));
 NAND2_X1 _37772_ (.A1(\core.keymem.key_mem[1][32] ),
    .A2(_14349_),
    .ZN(_14352_));
 OAI21_X1 _37773_ (.A(_14352_),
    .B1(_14232_),
    .B2(_12355_),
    .ZN(_01658_));
 NAND3_X1 _37774_ (.A1(_12751_),
    .A2(_13402_),
    .A3(_14235_),
    .ZN(_14353_));
 INV_X1 _37775_ (.A(\core.keymem.key_mem[1][33] ),
    .ZN(_14354_));
 OAI21_X1 _37776_ (.A(_14353_),
    .B1(_14220_),
    .B2(_14354_),
    .ZN(_01659_));
 NAND2_X1 _37777_ (.A1(\core.keymem.key_mem[1][34] ),
    .A2(_14349_),
    .ZN(_14355_));
 OAI21_X1 _37778_ (.A(_14355_),
    .B1(_14232_),
    .B2(_12376_),
    .ZN(_01660_));
 NAND2_X1 _37779_ (.A1(\core.keymem.key_mem[1][35] ),
    .A2(_14349_),
    .ZN(_14356_));
 OAI21_X1 _37780_ (.A(_14356_),
    .B1(_14216_),
    .B2(_12413_),
    .ZN(_01661_));
 MUX2_X1 _37781_ (.A(\core.keymem.key_mem[1][36] ),
    .B(_12423_),
    .S(_14262_),
    .Z(_01662_));
 NAND2_X1 _37782_ (.A1(\core.keymem.key_mem[1][37] ),
    .A2(_14349_),
    .ZN(_14357_));
 OAI21_X1 _37783_ (.A(_14357_),
    .B1(_14216_),
    .B2(_12439_),
    .ZN(_01663_));
 INV_X1 _37784_ (.A(\core.keymem.key_mem[1][38] ),
    .ZN(_14358_));
 OAI22_X1 _37785_ (.A1(_14358_),
    .A2(_14199_),
    .B1(_14200_),
    .B2(_12468_),
    .ZN(_01664_));
 NAND2_X1 _37786_ (.A1(\core.keymem.key_mem[1][39] ),
    .A2(_14349_),
    .ZN(_14359_));
 NAND2_X2 _37787_ (.A1(_00048_),
    .A2(_14264_),
    .ZN(_14360_));
 NAND3_X1 _37788_ (.A1(_14211_),
    .A2(_14235_),
    .A3(_14360_),
    .ZN(_14361_));
 OAI21_X1 _37789_ (.A(_14359_),
    .B1(_14361_),
    .B2(_13435_),
    .ZN(_01665_));
 BUF_X4 _37790_ (.A(_13132_),
    .Z(_14362_));
 OAI21_X2 _37791_ (.A(_13439_),
    .B1(_13440_),
    .B2(_12263_),
    .ZN(_14363_));
 NAND2_X1 _37792_ (.A1(\core.key[3] ),
    .A2(_12345_),
    .ZN(_14364_));
 NAND2_X1 _37793_ (.A1(_12158_),
    .A2(_14364_),
    .ZN(_14365_));
 XNOR2_X1 _37794_ (.A(_12796_),
    .B(_13444_),
    .ZN(_14366_));
 BUF_X4 _37795_ (.A(_12170_),
    .Z(_14367_));
 AOI21_X2 _37796_ (.A(_14365_),
    .B1(_14366_),
    .B2(_14367_),
    .ZN(_14368_));
 OAI221_X2 _37797_ (.A(_13439_),
    .B1(_13440_),
    .B2(_12263_),
    .C1(_12470_),
    .C2(_12185_),
    .ZN(_14369_));
 OAI22_X4 _37798_ (.A1(_14362_),
    .A2(_14363_),
    .B1(_14368_),
    .B2(_14369_),
    .ZN(_14370_));
 MUX2_X1 _37799_ (.A(\core.keymem.key_mem[1][3] ),
    .B(_14370_),
    .S(_14262_),
    .Z(_01666_));
 NAND2_X1 _37800_ (.A1(\core.keymem.key_mem[1][40] ),
    .A2(_14349_),
    .ZN(_14371_));
 NAND2_X1 _37801_ (.A1(_00049_),
    .A2(_14206_),
    .ZN(_14372_));
 NAND3_X1 _37802_ (.A1(_14211_),
    .A2(_14235_),
    .A3(_14372_),
    .ZN(_14373_));
 OAI21_X1 _37803_ (.A(_14371_),
    .B1(_14373_),
    .B2(_13457_),
    .ZN(_01667_));
 NAND3_X1 _37804_ (.A1(_12751_),
    .A2(_13467_),
    .A3(_14235_),
    .ZN(_14374_));
 BUF_X8 _37805_ (.A(_14198_),
    .Z(_14375_));
 INV_X1 _37806_ (.A(\core.keymem.key_mem[1][41] ),
    .ZN(_14376_));
 OAI21_X1 _37807_ (.A(_14374_),
    .B1(_14375_),
    .B2(_14376_),
    .ZN(_01668_));
 NAND2_X1 _37808_ (.A1(\core.keymem.key_mem[1][42] ),
    .A2(_14349_),
    .ZN(_14377_));
 OAI21_X4 _37809_ (.A(_13489_),
    .B1(_14248_),
    .B2(_12476_),
    .ZN(_14378_));
 OAI21_X1 _37810_ (.A(_14377_),
    .B1(_14378_),
    .B2(_14315_),
    .ZN(_01669_));
 NAND2_X1 _37811_ (.A1(\core.keymem.key_mem[1][43] ),
    .A2(_14349_),
    .ZN(_14379_));
 NAND2_X1 _37812_ (.A1(_00052_),
    .A2(_14238_),
    .ZN(_14380_));
 NAND3_X1 _37813_ (.A1(_14211_),
    .A2(_14235_),
    .A3(_14380_),
    .ZN(_14381_));
 OAI21_X1 _37814_ (.A(_14379_),
    .B1(_14381_),
    .B2(_13496_),
    .ZN(_01670_));
 NAND2_X1 _37815_ (.A1(\core.keymem.key_mem[1][44] ),
    .A2(_14349_),
    .ZN(_14382_));
 OAI21_X1 _37816_ (.A(_14382_),
    .B1(_14232_),
    .B2(_12506_),
    .ZN(_01671_));
 AND2_X1 _37817_ (.A1(_00054_),
    .A2(_14205_),
    .ZN(_14383_));
 NOR3_X1 _37818_ (.A1(_12183_),
    .A2(_14383_),
    .A3(_13509_),
    .ZN(_14384_));
 MUX2_X1 _37819_ (.A(\core.keymem.key_mem[1][45] ),
    .B(_14384_),
    .S(_14262_),
    .Z(_01672_));
 BUF_X4 _37820_ (.A(_14190_),
    .Z(_14385_));
 NAND2_X1 _37821_ (.A1(\core.keymem.key_mem[1][46] ),
    .A2(_14385_),
    .ZN(_14386_));
 NAND2_X1 _37822_ (.A1(_00055_),
    .A2(_14238_),
    .ZN(_14387_));
 NAND3_X1 _37823_ (.A1(_11986_),
    .A2(_14235_),
    .A3(_14387_),
    .ZN(_14388_));
 OAI21_X1 _37824_ (.A(_14386_),
    .B1(_14388_),
    .B2(_13517_),
    .ZN(_01673_));
 NAND2_X1 _37825_ (.A1(\core.keymem.key_mem[1][47] ),
    .A2(_14385_),
    .ZN(_14389_));
 OAI21_X1 _37826_ (.A(_14389_),
    .B1(_14232_),
    .B2(_12520_),
    .ZN(_01674_));
 NAND2_X1 _37827_ (.A1(\core.keymem.key_mem[1][48] ),
    .A2(_14385_),
    .ZN(_14390_));
 OAI21_X1 _37828_ (.A(_14390_),
    .B1(_14216_),
    .B2(_12532_),
    .ZN(_01675_));
 NAND2_X1 _37829_ (.A1(\core.keymem.key_mem[1][49] ),
    .A2(_14385_),
    .ZN(_14391_));
 NAND2_X2 _37830_ (.A1(_00058_),
    .A2(_14206_),
    .ZN(_14392_));
 NAND3_X1 _37831_ (.A1(_11986_),
    .A2(_14235_),
    .A3(_14392_),
    .ZN(_14393_));
 OAI21_X1 _37832_ (.A(_14391_),
    .B1(_14393_),
    .B2(_13529_),
    .ZN(_01676_));
 NAND2_X1 _37833_ (.A1(\core.keymem.key_mem[1][4] ),
    .A2(_14385_),
    .ZN(_14394_));
 NOR2_X1 _37834_ (.A1(_00375_),
    .A2(_11863_),
    .ZN(_14395_));
 AOI21_X1 _37835_ (.A(_14395_),
    .B1(_13415_),
    .B2(\core.key[4] ),
    .ZN(_14396_));
 NAND3_X1 _37836_ (.A1(_14274_),
    .A2(_13536_),
    .A3(_14396_),
    .ZN(_14397_));
 NAND2_X1 _37837_ (.A1(_12262_),
    .A2(_13533_),
    .ZN(_14398_));
 NAND2_X1 _37838_ (.A1(_00375_),
    .A2(_14282_),
    .ZN(_14399_));
 NAND3_X1 _37839_ (.A1(_14397_),
    .A2(_14398_),
    .A3(_14399_),
    .ZN(_14400_));
 OAI21_X1 _37840_ (.A(_14394_),
    .B1(_14400_),
    .B2(_14315_),
    .ZN(_01677_));
 NAND2_X1 _37841_ (.A1(\core.keymem.key_mem[1][50] ),
    .A2(_14385_),
    .ZN(_14401_));
 OAI21_X4 _37842_ (.A(_13556_),
    .B1(_14248_),
    .B2(_12536_),
    .ZN(_14402_));
 OAI21_X1 _37843_ (.A(_14401_),
    .B1(_14402_),
    .B2(_14315_),
    .ZN(_01678_));
 NAND2_X1 _37844_ (.A1(\core.keymem.key_mem[1][51] ),
    .A2(_14385_),
    .ZN(_14403_));
 BUF_X4 _37845_ (.A(_11936_),
    .Z(_14404_));
 MUX2_X1 _37846_ (.A(\core.key[51] ),
    .B(_13561_),
    .S(_12365_),
    .Z(_14405_));
 AOI221_X2 _37847_ (.A(_13558_),
    .B1(_13101_),
    .B2(_12028_),
    .C1(_14404_),
    .C2(_14405_),
    .ZN(_14406_));
 OAI21_X1 _37848_ (.A(_14403_),
    .B1(_14216_),
    .B2(_14406_),
    .ZN(_01679_));
 NAND2_X1 _37849_ (.A1(\core.keymem.key_mem[1][52] ),
    .A2(_14385_),
    .ZN(_14407_));
 BUF_X4 _37850_ (.A(_14200_),
    .Z(_14408_));
 OAI21_X1 _37851_ (.A(_14407_),
    .B1(_14408_),
    .B2(_12568_),
    .ZN(_01680_));
 NAND2_X1 _37852_ (.A1(\core.keymem.key_mem[1][53] ),
    .A2(_14385_),
    .ZN(_14409_));
 OAI21_X1 _37853_ (.A(_14409_),
    .B1(_14408_),
    .B2(_12584_),
    .ZN(_01681_));
 INV_X1 _37854_ (.A(\core.keymem.key_mem[1][54] ),
    .ZN(_14410_));
 OAI22_X1 _37855_ (.A1(_14410_),
    .A2(_14199_),
    .B1(_14200_),
    .B2(_13574_),
    .ZN(_01682_));
 NAND2_X2 _37856_ (.A1(_00064_),
    .A2(_14206_),
    .ZN(_14411_));
 NAND4_X1 _37857_ (.A1(_14211_),
    .A2(_13581_),
    .A3(_14227_),
    .A4(_14411_),
    .ZN(_14412_));
 INV_X1 _37858_ (.A(\core.keymem.key_mem[1][55] ),
    .ZN(_14413_));
 OAI21_X1 _37859_ (.A(_14412_),
    .B1(_14375_),
    .B2(_14413_),
    .ZN(_01683_));
 NOR2_X2 _37860_ (.A1(_12588_),
    .A2(_13875_),
    .ZN(_14414_));
 NOR4_X1 _37861_ (.A1(_11805_),
    .A2(_13583_),
    .A3(_13587_),
    .A4(_14414_),
    .ZN(_14415_));
 MUX2_X1 _37862_ (.A(\core.keymem.key_mem[1][56] ),
    .B(_14415_),
    .S(_14262_),
    .Z(_01684_));
 NAND2_X2 _37863_ (.A1(_00067_),
    .A2(_14212_),
    .ZN(_14416_));
 NAND3_X1 _37864_ (.A1(_13604_),
    .A2(_14193_),
    .A3(_14416_),
    .ZN(_14417_));
 INV_X1 _37865_ (.A(\core.keymem.key_mem[1][57] ),
    .ZN(_14418_));
 OAI21_X1 _37866_ (.A(_14417_),
    .B1(_14375_),
    .B2(_14418_),
    .ZN(_01685_));
 NOR2_X4 _37867_ (.A1(_00069_),
    .A2(_13331_),
    .ZN(_14419_));
 OAI21_X1 _37868_ (.A(_14217_),
    .B1(_14419_),
    .B2(_13611_),
    .ZN(_14420_));
 INV_X1 _37869_ (.A(\core.keymem.key_mem[1][58] ),
    .ZN(_14421_));
 OAI21_X1 _37870_ (.A(_14420_),
    .B1(_14375_),
    .B2(_14421_),
    .ZN(_01686_));
 NAND2_X1 _37871_ (.A1(\core.keymem.key_mem[1][59] ),
    .A2(_14385_),
    .ZN(_14422_));
 NOR2_X4 _37872_ (.A1(_00071_),
    .A2(_12871_),
    .ZN(_14423_));
 AOI21_X2 _37873_ (.A(_14423_),
    .B1(_13615_),
    .B2(_14201_),
    .ZN(_14424_));
 OAI21_X1 _37874_ (.A(_14422_),
    .B1(_14408_),
    .B2(_14424_),
    .ZN(_01687_));
 AOI22_X1 _37875_ (.A1(\core.keymem.key_mem[1][5] ),
    .A2(_14224_),
    .B1(_14193_),
    .B2(_12606_),
    .ZN(_14425_));
 INV_X1 _37876_ (.A(_14425_),
    .ZN(_01688_));
 NAND4_X1 _37877_ (.A1(_16285_),
    .A2(_14248_),
    .A3(_13621_),
    .A4(_14198_),
    .ZN(_14426_));
 NOR2_X2 _37878_ (.A1(_00073_),
    .A2(_14222_),
    .ZN(_14427_));
 NAND2_X1 _37879_ (.A1(_14427_),
    .A2(_14198_),
    .ZN(_14428_));
 INV_X1 _37880_ (.A(\core.keymem.key_mem[1][60] ),
    .ZN(_14429_));
 OAI221_X1 _37881_ (.A(_14426_),
    .B1(_14428_),
    .B2(_11930_),
    .C1(_14429_),
    .C2(_14199_),
    .ZN(_01689_));
 BUF_X4 _37882_ (.A(_14190_),
    .Z(_14430_));
 NAND2_X1 _37883_ (.A1(\core.keymem.key_mem[1][61] ),
    .A2(_14430_),
    .ZN(_14431_));
 NAND2_X2 _37884_ (.A1(_00075_),
    .A2(_14264_),
    .ZN(_14432_));
 NAND3_X1 _37885_ (.A1(_11986_),
    .A2(_14235_),
    .A3(_14432_),
    .ZN(_14433_));
 OR4_X4 _37886_ (.A1(_13624_),
    .A2(_13627_),
    .A3(_13629_),
    .A4(_13630_),
    .ZN(_14434_));
 OAI21_X1 _37887_ (.A(_14431_),
    .B1(_14433_),
    .B2(_14434_),
    .ZN(_01690_));
 NAND2_X1 _37888_ (.A1(\core.keymem.key_mem[1][62] ),
    .A2(_14430_),
    .ZN(_14435_));
 OAI22_X2 _37889_ (.A1(_00077_),
    .A2(_14245_),
    .B1(_12884_),
    .B2(_13635_),
    .ZN(_14436_));
 OR2_X1 _37890_ (.A1(_00078_),
    .A2(_12844_),
    .ZN(_14437_));
 OAI21_X1 _37891_ (.A(_14437_),
    .B1(_13633_),
    .B2(_14278_),
    .ZN(_14438_));
 BUF_X4 _37892_ (.A(_12336_),
    .Z(_14439_));
 AOI21_X2 _37893_ (.A(_14436_),
    .B1(_14438_),
    .B2(_14439_),
    .ZN(_14440_));
 OAI21_X1 _37894_ (.A(_14435_),
    .B1(_14408_),
    .B2(_14440_),
    .ZN(_01691_));
 NOR2_X4 _37895_ (.A1(_00079_),
    .A2(_13331_),
    .ZN(_14441_));
 OAI21_X1 _37896_ (.A(_14217_),
    .B1(_14441_),
    .B2(_13659_),
    .ZN(_14442_));
 INV_X1 _37897_ (.A(\core.keymem.key_mem[1][63] ),
    .ZN(_14443_));
 OAI21_X1 _37898_ (.A(_14442_),
    .B1(_14375_),
    .B2(_14443_),
    .ZN(_01692_));
 NAND2_X1 _37899_ (.A1(_12622_),
    .A2(_14217_),
    .ZN(_14444_));
 INV_X1 _37900_ (.A(\core.keymem.key_mem[1][64] ),
    .ZN(_14445_));
 OAI21_X1 _37901_ (.A(_14444_),
    .B1(_14375_),
    .B2(_14445_),
    .ZN(_01693_));
 NAND2_X1 _37902_ (.A1(\core.keymem.key_mem[1][65] ),
    .A2(_14430_),
    .ZN(_14446_));
 OAI21_X1 _37903_ (.A(_14446_),
    .B1(_14232_),
    .B2(_13673_),
    .ZN(_01694_));
 BUF_X4 _37904_ (.A(_11875_),
    .Z(_14447_));
 NOR2_X2 _37905_ (.A1(_00083_),
    .A2(_14447_),
    .ZN(_14448_));
 NOR2_X1 _37906_ (.A1(_14448_),
    .A2(_14189_),
    .ZN(_14449_));
 OR2_X1 _37907_ (.A1(_13677_),
    .A2(_13679_),
    .ZN(_14450_));
 INV_X1 _37908_ (.A(\core.keymem.key_mem[1][66] ),
    .ZN(_14451_));
 AOI221_X1 _37909_ (.A(_14335_),
    .B1(_14449_),
    .B2(_14450_),
    .C1(_14190_),
    .C2(_14451_),
    .ZN(_01695_));
 NAND2_X1 _37910_ (.A1(\core.keymem.key_mem[1][67] ),
    .A2(_14430_),
    .ZN(_14452_));
 OAI21_X1 _37911_ (.A(_11986_),
    .B1(_13687_),
    .B2(_13688_),
    .ZN(_14453_));
 OAI21_X1 _37912_ (.A(_14452_),
    .B1(_14453_),
    .B2(_14209_),
    .ZN(_01696_));
 NAND2_X1 _37913_ (.A1(\core.keymem.key_mem[1][68] ),
    .A2(_14430_),
    .ZN(_14454_));
 OAI21_X1 _37914_ (.A(_14454_),
    .B1(_14408_),
    .B2(_12635_),
    .ZN(_01697_));
 NAND2_X1 _37915_ (.A1(\core.keymem.key_mem[1][69] ),
    .A2(_14430_),
    .ZN(_14455_));
 OAI21_X1 _37916_ (.A(_14455_),
    .B1(_14408_),
    .B2(_13700_),
    .ZN(_01698_));
 AOI22_X1 _37917_ (.A1(\core.keymem.key_mem[1][6] ),
    .A2(_14224_),
    .B1(_14193_),
    .B2(_13711_),
    .ZN(_14456_));
 INV_X1 _37918_ (.A(_14456_),
    .ZN(_01699_));
 NAND2_X1 _37919_ (.A1(\core.keymem.key_mem[1][70] ),
    .A2(_14430_),
    .ZN(_14457_));
 OAI21_X1 _37920_ (.A(_14457_),
    .B1(_14408_),
    .B2(_12648_),
    .ZN(_01700_));
 NAND2_X1 _37921_ (.A1(\core.keymem.key_mem[1][71] ),
    .A2(_14430_),
    .ZN(_14458_));
 OAI21_X1 _37922_ (.A(_14458_),
    .B1(_14408_),
    .B2(_12659_),
    .ZN(_01701_));
 NAND2_X1 _37923_ (.A1(\core.keymem.key_mem[1][72] ),
    .A2(_14430_),
    .ZN(_14459_));
 OAI21_X1 _37924_ (.A(_14459_),
    .B1(_14232_),
    .B2(_12674_),
    .ZN(_01702_));
 NAND2_X1 _37925_ (.A1(\core.keymem.key_mem[1][73] ),
    .A2(_14430_),
    .ZN(_14460_));
 OAI21_X1 _37926_ (.A(_14460_),
    .B1(_14408_),
    .B2(_12688_),
    .ZN(_01703_));
 BUF_X4 _37927_ (.A(_14190_),
    .Z(_14461_));
 NAND2_X1 _37928_ (.A1(\core.keymem.key_mem[1][74] ),
    .A2(_14461_),
    .ZN(_14462_));
 NOR2_X2 _37929_ (.A1(_00091_),
    .A2(_14245_),
    .ZN(_14463_));
 BUF_X4 _37930_ (.A(_13415_),
    .Z(_14464_));
 AOI21_X1 _37931_ (.A(_13441_),
    .B1(\core.key[74] ),
    .B2(_14464_),
    .ZN(_14465_));
 OAI21_X2 _37932_ (.A(_14465_),
    .B1(_13723_),
    .B2(_14278_),
    .ZN(_14466_));
 AOI21_X4 _37933_ (.A(_11800_),
    .B1(_12854_),
    .B2(_12292_),
    .ZN(_14467_));
 AOI21_X4 _37934_ (.A(_14463_),
    .B1(_14466_),
    .B2(_14467_),
    .ZN(_14468_));
 OAI21_X1 _37935_ (.A(_14462_),
    .B1(_14468_),
    .B2(_14315_),
    .ZN(_01704_));
 NAND2_X1 _37936_ (.A1(\core.keymem.key_mem[1][75] ),
    .A2(_14461_),
    .ZN(_14469_));
 OAI21_X1 _37937_ (.A(_14469_),
    .B1(_14408_),
    .B2(_13733_),
    .ZN(_01705_));
 AOI22_X1 _37938_ (.A1(\core.keymem.key_mem[1][76] ),
    .A2(_14224_),
    .B1(_14192_),
    .B2(_13741_),
    .ZN(_14470_));
 INV_X1 _37939_ (.A(_14470_),
    .ZN(_01706_));
 NAND2_X1 _37940_ (.A1(\core.keymem.key_mem[1][77] ),
    .A2(_14461_),
    .ZN(_14471_));
 MUX2_X2 _37941_ (.A(_00094_),
    .B(_13749_),
    .S(_14245_),
    .Z(_14472_));
 OAI21_X1 _37942_ (.A(_14471_),
    .B1(_14472_),
    .B2(_14315_),
    .ZN(_01707_));
 NAND2_X1 _37943_ (.A1(\core.keymem.key_mem[1][78] ),
    .A2(_14461_),
    .ZN(_14473_));
 OAI21_X1 _37944_ (.A(_14473_),
    .B1(_14250_),
    .B2(_12708_),
    .ZN(_01708_));
 INV_X1 _37945_ (.A(\core.keymem.key_mem[1][79] ),
    .ZN(_14474_));
 NOR2_X2 _37946_ (.A1(_00096_),
    .A2(_12035_),
    .ZN(_14475_));
 AOI21_X4 _37947_ (.A(_14475_),
    .B1(_13756_),
    .B2(_13754_),
    .ZN(_14476_));
 OAI22_X1 _37948_ (.A1(_14474_),
    .A2(_14199_),
    .B1(_14200_),
    .B2(_14476_),
    .ZN(_01709_));
 NAND2_X1 _37949_ (.A1(\core.keymem.key_mem[1][7] ),
    .A2(_14461_),
    .ZN(_14477_));
 OAI21_X1 _37950_ (.A(_14477_),
    .B1(_14250_),
    .B2(_13767_),
    .ZN(_01710_));
 NAND2_X1 _37951_ (.A1(\core.keymem.key_mem[1][80] ),
    .A2(_14461_),
    .ZN(_14478_));
 OAI21_X1 _37952_ (.A(_14478_),
    .B1(_14250_),
    .B2(_12716_),
    .ZN(_01711_));
 NAND2_X1 _37953_ (.A1(\core.keymem.key_mem[1][81] ),
    .A2(_14461_),
    .ZN(_14479_));
 OAI21_X1 _37954_ (.A(_14479_),
    .B1(_14250_),
    .B2(_13775_),
    .ZN(_01712_));
 NAND2_X1 _37955_ (.A1(\core.keymem.key_mem[1][82] ),
    .A2(_14461_),
    .ZN(_14480_));
 OAI21_X1 _37956_ (.A(_14480_),
    .B1(_14250_),
    .B2(_13783_),
    .ZN(_01713_));
 NAND2_X1 _37957_ (.A1(\core.keymem.key_mem[1][83] ),
    .A2(_14461_),
    .ZN(_14481_));
 OAI21_X1 _37958_ (.A(_14481_),
    .B1(_14250_),
    .B2(_13791_),
    .ZN(_01714_));
 NAND2_X1 _37959_ (.A1(\core.keymem.key_mem[1][84] ),
    .A2(_14461_),
    .ZN(_14482_));
 OAI21_X1 _37960_ (.A(_14482_),
    .B1(_14250_),
    .B2(_12725_),
    .ZN(_01715_));
 NAND2_X1 _37961_ (.A1(\core.keymem.key_mem[1][85] ),
    .A2(_14191_),
    .ZN(_14483_));
 AOI21_X4 _37962_ (.A(_13793_),
    .B1(_13796_),
    .B2(_14248_),
    .ZN(_14484_));
 OAI21_X1 _37963_ (.A(_14483_),
    .B1(_14484_),
    .B2(_14315_),
    .ZN(_01716_));
 AOI22_X1 _37964_ (.A1(\core.keymem.key_mem[1][86] ),
    .A2(_14224_),
    .B1(_14192_),
    .B2(_12741_),
    .ZN(_14485_));
 INV_X1 _37965_ (.A(_14485_),
    .ZN(_01717_));
 INV_X1 _37966_ (.A(\core.keymem.key_mem[1][87] ),
    .ZN(_14486_));
 NOR2_X2 _37967_ (.A1(_00104_),
    .A2(_12002_),
    .ZN(_14487_));
 BUF_X8 _37968_ (.A(_12262_),
    .Z(_14488_));
 AOI21_X2 _37969_ (.A(_14487_),
    .B1(_13803_),
    .B2(_14488_),
    .ZN(_14489_));
 OAI22_X1 _37970_ (.A1(_14486_),
    .A2(_14199_),
    .B1(_14200_),
    .B2(_14489_),
    .ZN(_01718_));
 NAND2_X1 _37971_ (.A1(_00105_),
    .A2(_14212_),
    .ZN(_14490_));
 NAND4_X1 _37972_ (.A1(_14211_),
    .A2(_13810_),
    .A3(_14227_),
    .A4(_14490_),
    .ZN(_14491_));
 INV_X1 _37973_ (.A(\core.keymem.key_mem[1][88] ),
    .ZN(_14492_));
 OAI21_X1 _37974_ (.A(_14491_),
    .B1(_14375_),
    .B2(_14492_),
    .ZN(_01719_));
 NAND2_X1 _37975_ (.A1(\core.keymem.key_mem[1][89] ),
    .A2(_14191_),
    .ZN(_14493_));
 NAND2_X1 _37976_ (.A1(_00107_),
    .A2(_14206_),
    .ZN(_14494_));
 NAND3_X1 _37977_ (.A1(_11986_),
    .A2(_13818_),
    .A3(_14494_),
    .ZN(_14495_));
 OAI21_X1 _37978_ (.A(_14493_),
    .B1(_14495_),
    .B2(_14209_),
    .ZN(_01720_));
 NAND2_X1 _37979_ (.A1(\core.keymem.key_mem[1][8] ),
    .A2(_14191_),
    .ZN(_14496_));
 NAND2_X1 _37980_ (.A1(_00381_),
    .A2(_14206_),
    .ZN(_14497_));
 NAND3_X1 _37981_ (.A1(_11986_),
    .A2(_14227_),
    .A3(_14497_),
    .ZN(_14498_));
 NAND3_X2 _37982_ (.A1(_13819_),
    .A2(_13826_),
    .A3(_13833_),
    .ZN(_14499_));
 NOR2_X1 _37983_ (.A1(_13839_),
    .A2(_13842_),
    .ZN(_14500_));
 AND2_X1 _37984_ (.A1(_13846_),
    .A2(_13849_),
    .ZN(_14501_));
 AOI21_X2 _37985_ (.A(_14277_),
    .B1(_14500_),
    .B2(_14501_),
    .ZN(_14502_));
 XNOR2_X2 _37986_ (.A(_07262_),
    .B(_13455_),
    .ZN(_14503_));
 OAI22_X4 _37987_ (.A1(_14499_),
    .A2(_14502_),
    .B1(_14503_),
    .B2(_12884_),
    .ZN(_14504_));
 OAI21_X1 _37988_ (.A(_14496_),
    .B1(_14498_),
    .B2(_14504_),
    .ZN(_01721_));
 NAND2_X2 _37989_ (.A1(_00109_),
    .A2(_14212_),
    .ZN(_14505_));
 NAND4_X1 _37990_ (.A1(_14211_),
    .A2(_13860_),
    .A3(_14227_),
    .A4(_14505_),
    .ZN(_14506_));
 INV_X1 _37991_ (.A(\core.keymem.key_mem[1][90] ),
    .ZN(_14507_));
 OAI21_X1 _37992_ (.A(_14506_),
    .B1(_14375_),
    .B2(_14507_),
    .ZN(_01722_));
 NAND2_X1 _37993_ (.A1(\core.keymem.key_mem[1][91] ),
    .A2(_14191_),
    .ZN(_14508_));
 NAND2_X1 _37994_ (.A1(_00111_),
    .A2(_14242_),
    .ZN(_14509_));
 NAND3_X4 _37995_ (.A1(_13864_),
    .A2(_13868_),
    .A3(_14509_),
    .ZN(_14510_));
 OAI21_X1 _37996_ (.A(_14508_),
    .B1(_14510_),
    .B2(_14315_),
    .ZN(_01723_));
 NAND2_X1 _37997_ (.A1(\core.keymem.key_mem[1][92] ),
    .A2(_14191_),
    .ZN(_14511_));
 OAI22_X4 _37998_ (.A1(_12752_),
    .A2(_14201_),
    .B1(_13874_),
    .B2(_13878_),
    .ZN(_14512_));
 OAI21_X1 _37999_ (.A(_14511_),
    .B1(_14512_),
    .B2(_14315_),
    .ZN(_01724_));
 NAND2_X1 _38000_ (.A1(\core.keymem.key_mem[1][93] ),
    .A2(_14191_),
    .ZN(_14513_));
 NAND2_X2 _38001_ (.A1(_00115_),
    .A2(_14264_),
    .ZN(_14514_));
 NAND3_X1 _38002_ (.A1(_11986_),
    .A2(_14227_),
    .A3(_14514_),
    .ZN(_14515_));
 OR2_X1 _38003_ (.A1(_12307_),
    .A2(_11892_),
    .ZN(_14516_));
 NAND2_X1 _38004_ (.A1(_12307_),
    .A2(_12099_),
    .ZN(_14517_));
 MUX2_X1 _38005_ (.A(_14516_),
    .B(_14517_),
    .S(_12306_),
    .Z(_14518_));
 AOI21_X1 _38006_ (.A(_11847_),
    .B1(_00116_),
    .B2(_13415_),
    .ZN(_14519_));
 AOI221_X2 _38007_ (.A(_14205_),
    .B1(_14518_),
    .B2(_14519_),
    .C1(_13881_),
    .C2(_13441_),
    .ZN(_14520_));
 OAI21_X1 _38008_ (.A(_14513_),
    .B1(_14515_),
    .B2(_14520_),
    .ZN(_01725_));
 NAND2_X2 _38009_ (.A1(_00117_),
    .A2(_14205_),
    .ZN(_14521_));
 NAND4_X1 _38010_ (.A1(_14211_),
    .A2(_13896_),
    .A3(_14521_),
    .A4(_14227_),
    .ZN(_14522_));
 INV_X1 _38011_ (.A(\core.keymem.key_mem[1][94] ),
    .ZN(_14523_));
 OAI21_X1 _38012_ (.A(_14522_),
    .B1(_14375_),
    .B2(_14523_),
    .ZN(_01726_));
 NAND2_X2 _38013_ (.A1(_00119_),
    .A2(_14212_),
    .ZN(_14524_));
 NAND3_X1 _38014_ (.A1(_13903_),
    .A2(_14193_),
    .A3(_14524_),
    .ZN(_14525_));
 INV_X1 _38015_ (.A(\core.keymem.key_mem[1][95] ),
    .ZN(_14526_));
 OAI21_X1 _38016_ (.A(_14525_),
    .B1(_14375_),
    .B2(_14526_),
    .ZN(_01727_));
 NOR2_X1 _38017_ (.A1(_14304_),
    .A2(_13905_),
    .ZN(_14527_));
 NOR2_X1 _38018_ (.A1(_12758_),
    .A2(_12871_),
    .ZN(_14528_));
 NOR3_X1 _38019_ (.A1(_12183_),
    .A2(_14527_),
    .A3(_14528_),
    .ZN(_14529_));
 MUX2_X1 _38020_ (.A(\core.keymem.key_mem[1][96] ),
    .B(_14529_),
    .S(_14198_),
    .Z(_01728_));
 NAND2_X1 _38021_ (.A1(\core.keymem.key_mem[1][97] ),
    .A2(_14191_),
    .ZN(_14530_));
 OAI21_X1 _38022_ (.A(_14530_),
    .B1(_14232_),
    .B2(_12777_),
    .ZN(_01729_));
 NAND2_X1 _38023_ (.A1(\core.keymem.key_mem[1][98] ),
    .A2(_14191_),
    .ZN(_14531_));
 OAI21_X1 _38024_ (.A(_14531_),
    .B1(_14232_),
    .B2(_12788_),
    .ZN(_01730_));
 MUX2_X1 _38025_ (.A(\core.keymem.key_mem[1][99] ),
    .B(_12800_),
    .S(_14198_),
    .Z(_01731_));
 NOR2_X4 _38026_ (.A1(_00404_),
    .A2(_12185_),
    .ZN(_14532_));
 OAI21_X1 _38027_ (.A(_14217_),
    .B1(_14532_),
    .B2(_13919_),
    .ZN(_14533_));
 INV_X1 _38028_ (.A(\core.keymem.key_mem[1][9] ),
    .ZN(_14534_));
 OAI21_X1 _38029_ (.A(_14533_),
    .B1(_14199_),
    .B2(_14534_),
    .ZN(_01732_));
 NOR3_X1 _38030_ (.A1(_11794_),
    .A2(_16218_),
    .A3(_12804_),
    .ZN(_14535_));
 BUF_X4 _38031_ (.A(_14535_),
    .Z(_14536_));
 BUF_X4 _38032_ (.A(_14536_),
    .Z(_14537_));
 MUX2_X1 _38033_ (.A(\core.keymem.key_mem[2][0] ),
    .B(_11844_),
    .S(_14537_),
    .Z(_01733_));
 MUX2_X1 _38034_ (.A(\core.keymem.key_mem[2][100] ),
    .B(_11873_),
    .S(_14537_),
    .Z(_01734_));
 NAND3_X4 _38035_ (.A1(_16228_),
    .A2(_16216_),
    .A3(_11812_),
    .ZN(_14538_));
 BUF_X4 _38036_ (.A(_14538_),
    .Z(_14539_));
 BUF_X4 _38037_ (.A(_14539_),
    .Z(_14540_));
 NAND2_X1 _38038_ (.A1(\core.keymem.key_mem[2][101] ),
    .A2(_14540_),
    .ZN(_14541_));
 BUF_X4 _38039_ (.A(_14539_),
    .Z(_14542_));
 OAI21_X1 _38040_ (.A(_14541_),
    .B1(_14542_),
    .B2(_14202_),
    .ZN(_01735_));
 MUX2_X1 _38041_ (.A(\core.keymem.key_mem[2][102] ),
    .B(_11906_),
    .S(_14537_),
    .Z(_01736_));
 MUX2_X1 _38042_ (.A(\core.keymem.key_mem[2][103] ),
    .B(_11929_),
    .S(_14537_),
    .Z(_01737_));
 AOI21_X1 _38043_ (.A(_12821_),
    .B1(_14206_),
    .B2(_00133_),
    .ZN(_14543_));
 MUX2_X1 _38044_ (.A(\core.keymem.key_mem[2][104] ),
    .B(_14543_),
    .S(_14537_),
    .Z(_01738_));
 AND2_X1 _38045_ (.A1(_12829_),
    .A2(_14213_),
    .ZN(_14544_));
 MUX2_X1 _38046_ (.A(\core.keymem.key_mem[2][105] ),
    .B(_14544_),
    .S(_14537_),
    .Z(_01739_));
 MUX2_X1 _38047_ (.A(\core.keymem.key_mem[2][106] ),
    .B(_12832_),
    .S(_14537_),
    .Z(_01740_));
 MUX2_X1 _38048_ (.A(\core.keymem.key_mem[2][107] ),
    .B(_11967_),
    .S(_14537_),
    .Z(_01741_));
 MUX2_X1 _38049_ (.A(\core.keymem.key_mem[2][108] ),
    .B(_11981_),
    .S(_14537_),
    .Z(_01742_));
 AND2_X1 _38050_ (.A1(_12841_),
    .A2(_14218_),
    .ZN(_14545_));
 MUX2_X1 _38051_ (.A(\core.keymem.key_mem[2][109] ),
    .B(_14545_),
    .S(_14537_),
    .Z(_01743_));
 AOI21_X2 _38052_ (.A(_14229_),
    .B1(_12849_),
    .B2(_14367_),
    .ZN(_14546_));
 OAI21_X2 _38053_ (.A(_12871_),
    .B1(_12856_),
    .B2(_14274_),
    .ZN(_14547_));
 OAI22_X4 _38054_ (.A1(_11983_),
    .A2(_14488_),
    .B1(_14546_),
    .B2(_14547_),
    .ZN(_14548_));
 BUF_X4 _38055_ (.A(_14536_),
    .Z(_14549_));
 MUX2_X1 _38056_ (.A(\core.keymem.key_mem[2][10] ),
    .B(_14548_),
    .S(_14549_),
    .Z(_01744_));
 MUX2_X1 _38057_ (.A(\core.keymem.key_mem[2][110] ),
    .B(_12859_),
    .S(_14549_),
    .Z(_01745_));
 MUX2_X1 _38058_ (.A(\core.keymem.key_mem[2][111] ),
    .B(_12017_),
    .S(_14549_),
    .Z(_01746_));
 MUX2_X1 _38059_ (.A(\core.keymem.key_mem[2][112] ),
    .B(_12031_),
    .S(_14549_),
    .Z(_01747_));
 NAND2_X1 _38060_ (.A1(\core.keymem.key_mem[2][113] ),
    .A2(_14540_),
    .ZN(_14550_));
 BUF_X4 _38061_ (.A(_14536_),
    .Z(_14551_));
 NAND2_X1 _38062_ (.A1(_14236_),
    .A2(_14551_),
    .ZN(_14552_));
 OAI21_X1 _38063_ (.A(_14550_),
    .B1(_14552_),
    .B2(_14239_),
    .ZN(_01748_));
 MUX2_X1 _38064_ (.A(\core.keymem.key_mem[2][114] ),
    .B(_12869_),
    .S(_14549_),
    .Z(_01749_));
 MUX2_X1 _38065_ (.A(\core.keymem.key_mem[2][115] ),
    .B(_12059_),
    .S(_14549_),
    .Z(_01750_));
 MUX2_X1 _38066_ (.A(\core.keymem.key_mem[2][116] ),
    .B(_12077_),
    .S(_14549_),
    .Z(_01751_));
 INV_X1 _38067_ (.A(\core.keymem.key_mem[2][117] ),
    .ZN(_14553_));
 NAND2_X1 _38068_ (.A1(_14243_),
    .A2(_14551_),
    .ZN(_14554_));
 OAI22_X1 _38069_ (.A1(_14553_),
    .A2(_14551_),
    .B1(_14554_),
    .B2(_14246_),
    .ZN(_01752_));
 BUF_X4 _38070_ (.A(_14538_),
    .Z(_14555_));
 NAND2_X1 _38071_ (.A1(\core.keymem.key_mem[2][118] ),
    .A2(_14555_),
    .ZN(_14556_));
 OAI21_X1 _38072_ (.A(_14556_),
    .B1(_14542_),
    .B2(_14249_),
    .ZN(_01753_));
 MUX2_X1 _38073_ (.A(\core.keymem.key_mem[2][119] ),
    .B(_12096_),
    .S(_14549_),
    .Z(_01754_));
 NAND2_X1 _38074_ (.A1(\core.keymem.key_mem[2][11] ),
    .A2(_14555_),
    .ZN(_14557_));
 OAI21_X1 _38075_ (.A(_14557_),
    .B1(_14542_),
    .B2(_14255_),
    .ZN(_01755_));
 MUX2_X1 _38076_ (.A(\core.keymem.key_mem[2][120] ),
    .B(_12124_),
    .S(_14549_),
    .Z(_01756_));
 MUX2_X1 _38077_ (.A(\core.keymem.key_mem[2][121] ),
    .B(_12160_),
    .S(_14549_),
    .Z(_01757_));
 BUF_X4 _38078_ (.A(_14536_),
    .Z(_14558_));
 MUX2_X1 _38079_ (.A(\core.keymem.key_mem[2][122] ),
    .B(_12903_),
    .S(_14558_),
    .Z(_01758_));
 NAND2_X1 _38080_ (.A1(\core.keymem.key_mem[2][123] ),
    .A2(_14555_),
    .ZN(_14559_));
 OAI21_X1 _38081_ (.A(_14559_),
    .B1(_14542_),
    .B2(_12182_),
    .ZN(_01759_));
 NAND2_X1 _38082_ (.A1(\core.keymem.key_mem[2][124] ),
    .A2(_14555_),
    .ZN(_14560_));
 OAI21_X1 _38083_ (.A(_14560_),
    .B1(_14542_),
    .B2(_12926_),
    .ZN(_01760_));
 MUX2_X1 _38084_ (.A(\core.keymem.key_mem[2][125] ),
    .B(_12932_),
    .S(_14558_),
    .Z(_01761_));
 NAND2_X1 _38085_ (.A1(\core.keymem.key_mem[2][126] ),
    .A2(_14555_),
    .ZN(_14561_));
 OAI21_X1 _38086_ (.A(_14561_),
    .B1(_14542_),
    .B2(_12207_),
    .ZN(_01762_));
 MUX2_X1 _38087_ (.A(\core.keymem.key_mem[2][127] ),
    .B(_12945_),
    .S(_14558_),
    .Z(_01763_));
 NAND2_X1 _38088_ (.A1(\core.keymem.key_mem[2][12] ),
    .A2(_14555_),
    .ZN(_14562_));
 OAI21_X1 _38089_ (.A(_14562_),
    .B1(_14542_),
    .B2(_14281_),
    .ZN(_01764_));
 NAND2_X1 _38090_ (.A1(\core.keymem.key_mem[2][13] ),
    .A2(_14539_),
    .ZN(_14563_));
 NAND2_X1 _38091_ (.A1(_14226_),
    .A2(_14551_),
    .ZN(_14564_));
 OAI221_X1 _38092_ (.A(_14563_),
    .B1(_14539_),
    .B2(_14283_),
    .C1(_14290_),
    .C2(_14564_),
    .ZN(_01765_));
 NAND3_X1 _38093_ (.A1(_12978_),
    .A2(_11996_),
    .A3(_12980_),
    .ZN(_14565_));
 XOR2_X1 _38094_ (.A(_12978_),
    .B(_11992_),
    .Z(_14566_));
 MUX2_X1 _38095_ (.A(_14566_),
    .B(_14295_),
    .S(_12980_),
    .Z(_14567_));
 NOR2_X1 _38096_ (.A1(net11),
    .A2(_14567_),
    .ZN(_14568_));
 NOR3_X1 _38097_ (.A1(_12979_),
    .A2(_12698_),
    .A3(_14295_),
    .ZN(_14569_));
 AOI21_X1 _38098_ (.A(_14568_),
    .B1(_14569_),
    .B2(net11),
    .ZN(_14570_));
 AND4_X1 _38099_ (.A1(_14298_),
    .A2(_14299_),
    .A3(_14565_),
    .A4(_14570_),
    .ZN(_14571_));
 OAI21_X1 _38100_ (.A(_12951_),
    .B1(\core.key[14] ),
    .B2(_12302_),
    .ZN(_14572_));
 OAI22_X2 _38101_ (.A1(_13132_),
    .A2(_13004_),
    .B1(_14571_),
    .B2(_14572_),
    .ZN(_14573_));
 AND3_X1 _38102_ (.A1(_11952_),
    .A2(_14302_),
    .A3(_14573_),
    .ZN(_14574_));
 MUX2_X1 _38103_ (.A(\core.keymem.key_mem[2][14] ),
    .B(_14574_),
    .S(_14558_),
    .Z(_01766_));
 MUX2_X1 _38104_ (.A(\core.keymem.key_mem[2][15] ),
    .B(_14306_),
    .S(_14558_),
    .Z(_01767_));
 AND2_X1 _38105_ (.A1(_13028_),
    .A2(_14307_),
    .ZN(_14575_));
 MUX2_X1 _38106_ (.A(\core.keymem.key_mem[2][16] ),
    .B(_14575_),
    .S(_14558_),
    .Z(_01768_));
 NAND2_X1 _38107_ (.A1(\core.keymem.key_mem[2][17] ),
    .A2(_14555_),
    .ZN(_14576_));
 OAI21_X1 _38108_ (.A(_14576_),
    .B1(_14542_),
    .B2(_14314_),
    .ZN(_01769_));
 AND2_X1 _38109_ (.A1(_13093_),
    .A2(_14316_),
    .ZN(_14577_));
 MUX2_X1 _38110_ (.A(\core.keymem.key_mem[2][18] ),
    .B(_14577_),
    .S(_14558_),
    .Z(_01770_));
 NAND2_X1 _38111_ (.A1(\core.keymem.key_mem[2][19] ),
    .A2(_14555_),
    .ZN(_14578_));
 OAI21_X1 _38112_ (.A(_14578_),
    .B1(_14542_),
    .B2(_14322_),
    .ZN(_01771_));
 MUX2_X1 _38113_ (.A(\core.keymem.key_mem[2][1] ),
    .B(_14324_),
    .S(_14558_),
    .Z(_01772_));
 MUX2_X1 _38114_ (.A(\core.keymem.key_mem[2][20] ),
    .B(_14326_),
    .S(_14558_),
    .Z(_01773_));
 OR2_X1 _38115_ (.A1(_14328_),
    .A2(_14329_),
    .ZN(_14579_));
 MUX2_X1 _38116_ (.A(\core.keymem.key_mem[2][21] ),
    .B(_14579_),
    .S(_14558_),
    .Z(_01774_));
 NAND2_X1 _38117_ (.A1(_13190_),
    .A2(_14332_),
    .ZN(_14580_));
 BUF_X8 _38118_ (.A(_14536_),
    .Z(_14581_));
 MUX2_X1 _38119_ (.A(\core.keymem.key_mem[2][22] ),
    .B(_14580_),
    .S(_14581_),
    .Z(_01775_));
 NAND2_X1 _38120_ (.A1(\core.keymem.key_mem[2][23] ),
    .A2(_14555_),
    .ZN(_14582_));
 OAI21_X1 _38121_ (.A(_14582_),
    .B1(_14542_),
    .B2(_12272_),
    .ZN(_01776_));
 NAND2_X1 _38122_ (.A1(\core.keymem.key_mem[2][24] ),
    .A2(_14555_),
    .ZN(_14583_));
 BUF_X4 _38123_ (.A(_14539_),
    .Z(_14584_));
 OAI21_X1 _38124_ (.A(_14583_),
    .B1(_14584_),
    .B2(_13212_),
    .ZN(_01777_));
 AND2_X1 _38125_ (.A1(_13232_),
    .A2(_14338_),
    .ZN(_14585_));
 MUX2_X1 _38126_ (.A(\core.keymem.key_mem[2][25] ),
    .B(_14585_),
    .S(_14581_),
    .Z(_01778_));
 MUX2_X1 _38127_ (.A(\core.keymem.key_mem[2][26] ),
    .B(_13241_),
    .S(_14581_),
    .Z(_01779_));
 MUX2_X1 _38128_ (.A(\core.keymem.key_mem[2][27] ),
    .B(_13284_),
    .S(_14581_),
    .Z(_01780_));
 MUX2_X1 _38129_ (.A(\core.keymem.key_mem[2][28] ),
    .B(_13325_),
    .S(_14581_),
    .Z(_01781_));
 MUX2_X1 _38130_ (.A(\core.keymem.key_mem[2][29] ),
    .B(_13329_),
    .S(_14581_),
    .Z(_01782_));
 BUF_X4 _38131_ (.A(_14538_),
    .Z(_14586_));
 NAND2_X1 _38132_ (.A1(\core.keymem.key_mem[2][2] ),
    .A2(_14586_),
    .ZN(_14587_));
 OAI21_X1 _38133_ (.A(_14587_),
    .B1(_14584_),
    .B2(_12337_),
    .ZN(_01783_));
 MUX2_X1 _38134_ (.A(\core.keymem.key_mem[2][30] ),
    .B(_13379_),
    .S(_14581_),
    .Z(_01784_));
 MUX2_X1 _38135_ (.A(\core.keymem.key_mem[2][31] ),
    .B(_13395_),
    .S(_14581_),
    .Z(_01785_));
 MUX2_X1 _38136_ (.A(\core.keymem.key_mem[2][32] ),
    .B(_13396_),
    .S(_14581_),
    .Z(_01786_));
 MUX2_X1 _38137_ (.A(\core.keymem.key_mem[2][33] ),
    .B(_13402_),
    .S(_14581_),
    .Z(_01787_));
 BUF_X4 _38138_ (.A(_14536_),
    .Z(_14588_));
 MUX2_X1 _38139_ (.A(\core.keymem.key_mem[2][34] ),
    .B(_13403_),
    .S(_14588_),
    .Z(_01788_));
 MUX2_X1 _38140_ (.A(\core.keymem.key_mem[2][35] ),
    .B(_13405_),
    .S(_14588_),
    .Z(_01789_));
 NAND2_X1 _38141_ (.A1(\core.keymem.key_mem[2][36] ),
    .A2(_14586_),
    .ZN(_14589_));
 OAI21_X1 _38142_ (.A(_14589_),
    .B1(_14584_),
    .B2(_13407_),
    .ZN(_01790_));
 NAND2_X1 _38143_ (.A1(\core.keymem.key_mem[2][37] ),
    .A2(_14586_),
    .ZN(_14590_));
 OAI21_X1 _38144_ (.A(_14590_),
    .B1(_14584_),
    .B2(_12439_),
    .ZN(_01791_));
 MUX2_X1 _38145_ (.A(\core.keymem.key_mem[2][38] ),
    .B(_13410_),
    .S(_14588_),
    .Z(_01792_));
 NAND2_X1 _38146_ (.A1(\core.keymem.key_mem[2][39] ),
    .A2(_14586_),
    .ZN(_14591_));
 NAND2_X1 _38147_ (.A1(_14360_),
    .A2(_14551_),
    .ZN(_14592_));
 OAI21_X1 _38148_ (.A(_14591_),
    .B1(_14592_),
    .B2(_13435_),
    .ZN(_01793_));
 MUX2_X1 _38149_ (.A(\core.keymem.key_mem[2][3] ),
    .B(_14370_),
    .S(_14588_),
    .Z(_01794_));
 NAND2_X1 _38150_ (.A1(\core.keymem.key_mem[2][40] ),
    .A2(_14586_),
    .ZN(_14593_));
 NAND2_X1 _38151_ (.A1(_14372_),
    .A2(_14551_),
    .ZN(_14594_));
 OAI21_X1 _38152_ (.A(_14593_),
    .B1(_14594_),
    .B2(_13457_),
    .ZN(_01795_));
 MUX2_X1 _38153_ (.A(\core.keymem.key_mem[2][41] ),
    .B(_13467_),
    .S(_14588_),
    .Z(_01796_));
 NAND2_X1 _38154_ (.A1(\core.keymem.key_mem[2][42] ),
    .A2(_14586_),
    .ZN(_14595_));
 OAI21_X1 _38155_ (.A(_14595_),
    .B1(_14584_),
    .B2(_14378_),
    .ZN(_01797_));
 AOI21_X1 _38156_ (.A(_13495_),
    .B1(_14206_),
    .B2(_00052_),
    .ZN(_14596_));
 MUX2_X1 _38157_ (.A(\core.keymem.key_mem[2][43] ),
    .B(_14596_),
    .S(_14588_),
    .Z(_01798_));
 MUX2_X1 _38158_ (.A(\core.keymem.key_mem[2][44] ),
    .B(_13497_),
    .S(_14588_),
    .Z(_01799_));
 NAND2_X1 _38159_ (.A1(\core.keymem.key_mem[2][45] ),
    .A2(_14586_),
    .ZN(_14597_));
 OR2_X1 _38160_ (.A1(_14383_),
    .A2(_13509_),
    .ZN(_14598_));
 OAI21_X1 _38161_ (.A(_14597_),
    .B1(_14584_),
    .B2(_14598_),
    .ZN(_01800_));
 AOI21_X1 _38162_ (.A(_13516_),
    .B1(_14206_),
    .B2(_00055_),
    .ZN(_14599_));
 MUX2_X1 _38163_ (.A(\core.keymem.key_mem[2][46] ),
    .B(_14599_),
    .S(_14588_),
    .Z(_01801_));
 NAND2_X1 _38164_ (.A1(\core.keymem.key_mem[2][47] ),
    .A2(_14586_),
    .ZN(_14600_));
 OAI21_X1 _38165_ (.A(_14600_),
    .B1(_14584_),
    .B2(_12520_),
    .ZN(_01802_));
 NAND2_X1 _38166_ (.A1(\core.keymem.key_mem[2][48] ),
    .A2(_14586_),
    .ZN(_14601_));
 OAI21_X1 _38167_ (.A(_14601_),
    .B1(_14584_),
    .B2(_12532_),
    .ZN(_01803_));
 NAND2_X1 _38168_ (.A1(\core.keymem.key_mem[2][49] ),
    .A2(_14586_),
    .ZN(_14602_));
 NAND2_X1 _38169_ (.A1(_14392_),
    .A2(_14551_),
    .ZN(_14603_));
 OAI21_X1 _38170_ (.A(_14602_),
    .B1(_14603_),
    .B2(_13529_),
    .ZN(_01804_));
 AND3_X1 _38171_ (.A1(_14397_),
    .A2(_14398_),
    .A3(_14399_),
    .ZN(_14604_));
 MUX2_X1 _38172_ (.A(\core.keymem.key_mem[2][4] ),
    .B(_14604_),
    .S(_14588_),
    .Z(_01805_));
 BUF_X4 _38173_ (.A(_14538_),
    .Z(_14605_));
 NAND2_X1 _38174_ (.A1(\core.keymem.key_mem[2][50] ),
    .A2(_14605_),
    .ZN(_14606_));
 OAI21_X1 _38175_ (.A(_14606_),
    .B1(_14584_),
    .B2(_14402_),
    .ZN(_01806_));
 MUX2_X1 _38176_ (.A(\core.keymem.key_mem[2][51] ),
    .B(_13564_),
    .S(_14588_),
    .Z(_01807_));
 NAND2_X1 _38177_ (.A1(\core.keymem.key_mem[2][52] ),
    .A2(_14605_),
    .ZN(_14607_));
 OAI21_X1 _38178_ (.A(_14607_),
    .B1(_14584_),
    .B2(_12568_),
    .ZN(_01808_));
 NAND2_X1 _38179_ (.A1(\core.keymem.key_mem[2][53] ),
    .A2(_14605_),
    .ZN(_14608_));
 BUF_X4 _38180_ (.A(_14539_),
    .Z(_14609_));
 OAI21_X1 _38181_ (.A(_14608_),
    .B1(_14609_),
    .B2(_12584_),
    .ZN(_01809_));
 NAND2_X1 _38182_ (.A1(\core.keymem.key_mem[2][54] ),
    .A2(_14605_),
    .ZN(_14610_));
 OAI21_X1 _38183_ (.A(_14610_),
    .B1(_14609_),
    .B2(_13575_),
    .ZN(_01810_));
 NAND2_X1 _38184_ (.A1(\core.keymem.key_mem[2][55] ),
    .A2(_14605_),
    .ZN(_14611_));
 NAND2_X1 _38185_ (.A1(_13580_),
    .A2(_14411_),
    .ZN(_14612_));
 OAI21_X1 _38186_ (.A(_14611_),
    .B1(_14609_),
    .B2(_14612_),
    .ZN(_01811_));
 NOR3_X4 _38187_ (.A1(_13583_),
    .A2(_13587_),
    .A3(_14414_),
    .ZN(_14613_));
 BUF_X4 _38188_ (.A(_14536_),
    .Z(_14614_));
 MUX2_X1 _38189_ (.A(\core.keymem.key_mem[2][56] ),
    .B(_14613_),
    .S(_14614_),
    .Z(_01812_));
 AND2_X1 _38190_ (.A1(_13603_),
    .A2(_14416_),
    .ZN(_14615_));
 MUX2_X1 _38191_ (.A(\core.keymem.key_mem[2][57] ),
    .B(_14615_),
    .S(_14614_),
    .Z(_01813_));
 OR2_X1 _38192_ (.A1(_13610_),
    .A2(_14419_),
    .ZN(_14616_));
 MUX2_X1 _38193_ (.A(\core.keymem.key_mem[2][58] ),
    .B(_14616_),
    .S(_14614_),
    .Z(_01814_));
 NAND2_X1 _38194_ (.A1(\core.keymem.key_mem[2][59] ),
    .A2(_14605_),
    .ZN(_14617_));
 OAI21_X1 _38195_ (.A(_14617_),
    .B1(_14609_),
    .B2(_14424_),
    .ZN(_01815_));
 MUX2_X1 _38196_ (.A(\core.keymem.key_mem[2][5] ),
    .B(_12606_),
    .S(_14614_),
    .Z(_01816_));
 NAND2_X1 _38197_ (.A1(\core.keymem.key_mem[2][60] ),
    .A2(_14605_),
    .ZN(_14618_));
 AOI21_X1 _38198_ (.A(_14427_),
    .B1(_13621_),
    .B2(_14248_),
    .ZN(_14619_));
 OAI21_X1 _38199_ (.A(_14618_),
    .B1(_14609_),
    .B2(_14619_),
    .ZN(_01817_));
 NAND2_X1 _38200_ (.A1(\core.keymem.key_mem[2][61] ),
    .A2(_14605_),
    .ZN(_14620_));
 NAND2_X1 _38201_ (.A1(_14432_),
    .A2(_14551_),
    .ZN(_14621_));
 OAI21_X1 _38202_ (.A(_14620_),
    .B1(_14621_),
    .B2(_14434_),
    .ZN(_01818_));
 MUX2_X1 _38203_ (.A(\core.keymem.key_mem[2][62] ),
    .B(_13637_),
    .S(_14614_),
    .Z(_01819_));
 OR2_X1 _38204_ (.A1(_13658_),
    .A2(_14441_),
    .ZN(_14622_));
 MUX2_X1 _38205_ (.A(\core.keymem.key_mem[2][63] ),
    .B(_14622_),
    .S(_14614_),
    .Z(_01820_));
 MUX2_X1 _38206_ (.A(\core.keymem.key_mem[2][64] ),
    .B(_12622_),
    .S(_14614_),
    .Z(_01821_));
 NAND2_X1 _38207_ (.A1(\core.keymem.key_mem[2][65] ),
    .A2(_14605_),
    .ZN(_14623_));
 OAI21_X1 _38208_ (.A(_14623_),
    .B1(_14609_),
    .B2(_13673_),
    .ZN(_01822_));
 MUX2_X1 _38209_ (.A(\core.keymem.key_mem[2][66] ),
    .B(_13681_),
    .S(_14614_),
    .Z(_01823_));
 NAND2_X1 _38210_ (.A1(\core.keymem.key_mem[2][67] ),
    .A2(_14605_),
    .ZN(_14624_));
 OAI21_X1 _38211_ (.A(_14624_),
    .B1(_14609_),
    .B2(_13690_),
    .ZN(_01824_));
 BUF_X4 _38212_ (.A(_14538_),
    .Z(_14625_));
 NAND2_X1 _38213_ (.A1(\core.keymem.key_mem[2][68] ),
    .A2(_14625_),
    .ZN(_14626_));
 OAI21_X1 _38214_ (.A(_14626_),
    .B1(_14609_),
    .B2(_12635_),
    .ZN(_01825_));
 NAND2_X1 _38215_ (.A1(\core.keymem.key_mem[2][69] ),
    .A2(_14625_),
    .ZN(_14627_));
 OAI21_X1 _38216_ (.A(_14627_),
    .B1(_14609_),
    .B2(_13700_),
    .ZN(_01826_));
 MUX2_X1 _38217_ (.A(\core.keymem.key_mem[2][6] ),
    .B(_13711_),
    .S(_14614_),
    .Z(_01827_));
 MUX2_X1 _38218_ (.A(\core.keymem.key_mem[2][70] ),
    .B(_13713_),
    .S(_14614_),
    .Z(_01828_));
 NAND2_X1 _38219_ (.A1(\core.keymem.key_mem[2][71] ),
    .A2(_14625_),
    .ZN(_14628_));
 OAI21_X1 _38220_ (.A(_14628_),
    .B1(_14609_),
    .B2(_12659_),
    .ZN(_01829_));
 NAND2_X1 _38221_ (.A1(\core.keymem.key_mem[2][72] ),
    .A2(_14625_),
    .ZN(_14629_));
 BUF_X4 _38222_ (.A(_14539_),
    .Z(_14630_));
 OAI21_X1 _38223_ (.A(_14629_),
    .B1(_14630_),
    .B2(_13716_),
    .ZN(_01830_));
 NAND2_X1 _38224_ (.A1(\core.keymem.key_mem[2][73] ),
    .A2(_14625_),
    .ZN(_14631_));
 OAI21_X1 _38225_ (.A(_14631_),
    .B1(_14630_),
    .B2(_12688_),
    .ZN(_01831_));
 NAND2_X1 _38226_ (.A1(_06678_),
    .A2(_13722_),
    .ZN(_14632_));
 XNOR2_X2 _38227_ (.A(_13470_),
    .B(_11944_),
    .ZN(_14633_));
 AOI21_X2 _38228_ (.A(_14632_),
    .B1(_14633_),
    .B2(_14367_),
    .ZN(_14634_));
 INV_X1 _38229_ (.A(_14467_),
    .ZN(_14635_));
 OAI22_X4 _38230_ (.A1(_00091_),
    .A2(_14488_),
    .B1(_14634_),
    .B2(_14635_),
    .ZN(_14636_));
 BUF_X4 _38231_ (.A(_14536_),
    .Z(_14637_));
 MUX2_X1 _38232_ (.A(\core.keymem.key_mem[2][74] ),
    .B(_14636_),
    .S(_14637_),
    .Z(_01832_));
 NAND2_X1 _38233_ (.A1(\core.keymem.key_mem[2][75] ),
    .A2(_14625_),
    .ZN(_14638_));
 OAI21_X1 _38234_ (.A(_14638_),
    .B1(_14630_),
    .B2(_13733_),
    .ZN(_01833_));
 MUX2_X1 _38235_ (.A(\core.keymem.key_mem[2][76] ),
    .B(_13741_),
    .S(_14637_),
    .Z(_01834_));
 OAI21_X4 _38236_ (.A(_13744_),
    .B1(_13749_),
    .B2(_14264_),
    .ZN(_14639_));
 MUX2_X1 _38237_ (.A(\core.keymem.key_mem[2][77] ),
    .B(_14639_),
    .S(_14637_),
    .Z(_01835_));
 NAND2_X1 _38238_ (.A1(\core.keymem.key_mem[2][78] ),
    .A2(_14625_),
    .ZN(_14640_));
 OAI21_X1 _38239_ (.A(_14640_),
    .B1(_14630_),
    .B2(_12708_),
    .ZN(_01836_));
 NAND2_X1 _38240_ (.A1(\core.keymem.key_mem[2][79] ),
    .A2(_14625_),
    .ZN(_14641_));
 OAI21_X1 _38241_ (.A(_14641_),
    .B1(_14630_),
    .B2(_14476_),
    .ZN(_01837_));
 NAND2_X1 _38242_ (.A1(\core.keymem.key_mem[2][7] ),
    .A2(_14625_),
    .ZN(_14642_));
 OAI21_X1 _38243_ (.A(_14642_),
    .B1(_14630_),
    .B2(_13767_),
    .ZN(_01838_));
 MUX2_X1 _38244_ (.A(\core.keymem.key_mem[2][80] ),
    .B(_13769_),
    .S(_14637_),
    .Z(_01839_));
 NAND2_X1 _38245_ (.A1(\core.keymem.key_mem[2][81] ),
    .A2(_14625_),
    .ZN(_14643_));
 OAI21_X1 _38246_ (.A(_14643_),
    .B1(_14630_),
    .B2(_13775_),
    .ZN(_01840_));
 BUF_X4 _38247_ (.A(_14538_),
    .Z(_14644_));
 NAND2_X1 _38248_ (.A1(\core.keymem.key_mem[2][82] ),
    .A2(_14644_),
    .ZN(_14645_));
 OAI21_X1 _38249_ (.A(_14645_),
    .B1(_14630_),
    .B2(_13783_),
    .ZN(_01841_));
 NAND2_X1 _38250_ (.A1(\core.keymem.key_mem[2][83] ),
    .A2(_14644_),
    .ZN(_14646_));
 OAI21_X1 _38251_ (.A(_14646_),
    .B1(_14630_),
    .B2(_13791_),
    .ZN(_01842_));
 NAND2_X1 _38252_ (.A1(\core.keymem.key_mem[2][84] ),
    .A2(_14644_),
    .ZN(_14647_));
 OAI21_X1 _38253_ (.A(_14647_),
    .B1(_14630_),
    .B2(_12725_),
    .ZN(_01843_));
 NAND2_X1 _38254_ (.A1(\core.keymem.key_mem[2][85] ),
    .A2(_14644_),
    .ZN(_14648_));
 OAI21_X1 _38255_ (.A(_14648_),
    .B1(_14540_),
    .B2(_14484_),
    .ZN(_01844_));
 MUX2_X1 _38256_ (.A(\core.keymem.key_mem[2][86] ),
    .B(_12741_),
    .S(_14637_),
    .Z(_01845_));
 NAND2_X1 _38257_ (.A1(\core.keymem.key_mem[2][87] ),
    .A2(_14644_),
    .ZN(_14649_));
 OAI21_X1 _38258_ (.A(_14649_),
    .B1(_14540_),
    .B2(_14489_),
    .ZN(_01846_));
 AND2_X1 _38259_ (.A1(_13809_),
    .A2(_14490_),
    .ZN(_14650_));
 MUX2_X1 _38260_ (.A(\core.keymem.key_mem[2][88] ),
    .B(_14650_),
    .S(_14637_),
    .Z(_01847_));
 NAND2_X1 _38261_ (.A1(\core.keymem.key_mem[2][89] ),
    .A2(_14644_),
    .ZN(_14651_));
 NAND2_X1 _38262_ (.A1(_13817_),
    .A2(_14494_),
    .ZN(_14652_));
 OAI21_X1 _38263_ (.A(_14651_),
    .B1(_14540_),
    .B2(_14652_),
    .ZN(_01848_));
 NAND2_X1 _38264_ (.A1(\core.keymem.key_mem[2][8] ),
    .A2(_14644_),
    .ZN(_14653_));
 NAND2_X1 _38265_ (.A1(_14497_),
    .A2(_14551_),
    .ZN(_14654_));
 OAI21_X1 _38266_ (.A(_14653_),
    .B1(_14654_),
    .B2(_14504_),
    .ZN(_01849_));
 AND2_X1 _38267_ (.A1(_13859_),
    .A2(_14505_),
    .ZN(_14655_));
 MUX2_X1 _38268_ (.A(\core.keymem.key_mem[2][90] ),
    .B(_14655_),
    .S(_14637_),
    .Z(_01850_));
 NAND2_X1 _38269_ (.A1(\core.keymem.key_mem[2][91] ),
    .A2(_14644_),
    .ZN(_14656_));
 OAI21_X1 _38270_ (.A(_14656_),
    .B1(_14540_),
    .B2(_14510_),
    .ZN(_01851_));
 NAND2_X1 _38271_ (.A1(\core.keymem.key_mem[2][92] ),
    .A2(_14644_),
    .ZN(_14657_));
 OAI21_X1 _38272_ (.A(_14657_),
    .B1(_14540_),
    .B2(_14512_),
    .ZN(_01852_));
 NAND2_X1 _38273_ (.A1(\core.keymem.key_mem[2][93] ),
    .A2(_14644_),
    .ZN(_14658_));
 NAND2_X1 _38274_ (.A1(_14514_),
    .A2(_14551_),
    .ZN(_14659_));
 OAI21_X1 _38275_ (.A(_14658_),
    .B1(_14659_),
    .B2(_14520_),
    .ZN(_01853_));
 AND2_X1 _38276_ (.A1(_13895_),
    .A2(_14521_),
    .ZN(_14660_));
 MUX2_X1 _38277_ (.A(\core.keymem.key_mem[2][94] ),
    .B(_14660_),
    .S(_14637_),
    .Z(_01854_));
 AND2_X1 _38278_ (.A1(_13902_),
    .A2(_14524_),
    .ZN(_14661_));
 MUX2_X1 _38279_ (.A(\core.keymem.key_mem[2][95] ),
    .B(_14661_),
    .S(_14637_),
    .Z(_01855_));
 NAND2_X1 _38280_ (.A1(\core.keymem.key_mem[2][96] ),
    .A2(_14539_),
    .ZN(_14662_));
 OR2_X1 _38281_ (.A1(_14527_),
    .A2(_14528_),
    .ZN(_14663_));
 OAI21_X1 _38282_ (.A(_14662_),
    .B1(_14540_),
    .B2(_14663_),
    .ZN(_01856_));
 NAND2_X1 _38283_ (.A1(\core.keymem.key_mem[2][97] ),
    .A2(_14539_),
    .ZN(_14664_));
 OAI21_X1 _38284_ (.A(_14664_),
    .B1(_14540_),
    .B2(_12777_),
    .ZN(_01857_));
 NAND2_X1 _38285_ (.A1(\core.keymem.key_mem[2][98] ),
    .A2(_14539_),
    .ZN(_14665_));
 OAI21_X1 _38286_ (.A(_14665_),
    .B1(_14540_),
    .B2(_13910_),
    .ZN(_01858_));
 MUX2_X1 _38287_ (.A(\core.keymem.key_mem[2][99] ),
    .B(_12800_),
    .S(_14637_),
    .Z(_01859_));
 OR2_X1 _38288_ (.A1(_13918_),
    .A2(_14532_),
    .ZN(_14666_));
 MUX2_X1 _38289_ (.A(\core.keymem.key_mem[2][9] ),
    .B(_14666_),
    .S(_14536_),
    .Z(_01860_));
 NOR3_X2 _38290_ (.A1(_11794_),
    .A2(_16218_),
    .A3(_13921_),
    .ZN(_14667_));
 BUF_X8 _38291_ (.A(_14667_),
    .Z(_14668_));
 BUF_X4 _38292_ (.A(_14668_),
    .Z(_14669_));
 MUX2_X1 _38293_ (.A(\core.keymem.key_mem[3][0] ),
    .B(_11844_),
    .S(_14669_),
    .Z(_01861_));
 MUX2_X1 _38294_ (.A(\core.keymem.key_mem[3][100] ),
    .B(_11873_),
    .S(_14669_),
    .Z(_01862_));
 NAND3_X4 _38295_ (.A1(_16229_),
    .A2(_13920_),
    .A3(_11812_),
    .ZN(_14670_));
 BUF_X4 _38296_ (.A(_14670_),
    .Z(_14671_));
 BUF_X4 _38297_ (.A(_14671_),
    .Z(_14672_));
 NAND2_X1 _38298_ (.A1(\core.keymem.key_mem[3][101] ),
    .A2(_14672_),
    .ZN(_14673_));
 BUF_X4 _38299_ (.A(_14671_),
    .Z(_14674_));
 OAI21_X1 _38300_ (.A(_14673_),
    .B1(_14674_),
    .B2(_14202_),
    .ZN(_01863_));
 MUX2_X1 _38301_ (.A(\core.keymem.key_mem[3][102] ),
    .B(_11906_),
    .S(_14669_),
    .Z(_01864_));
 MUX2_X1 _38302_ (.A(\core.keymem.key_mem[3][103] ),
    .B(_11929_),
    .S(_14669_),
    .Z(_01865_));
 MUX2_X1 _38303_ (.A(\core.keymem.key_mem[3][104] ),
    .B(_14543_),
    .S(_14669_),
    .Z(_01866_));
 MUX2_X1 _38304_ (.A(\core.keymem.key_mem[3][105] ),
    .B(_14544_),
    .S(_14669_),
    .Z(_01867_));
 MUX2_X1 _38305_ (.A(\core.keymem.key_mem[3][106] ),
    .B(_12832_),
    .S(_14669_),
    .Z(_01868_));
 MUX2_X1 _38306_ (.A(\core.keymem.key_mem[3][107] ),
    .B(_11967_),
    .S(_14669_),
    .Z(_01869_));
 MUX2_X1 _38307_ (.A(\core.keymem.key_mem[3][108] ),
    .B(_11981_),
    .S(_14669_),
    .Z(_01870_));
 BUF_X4 _38308_ (.A(_14668_),
    .Z(_14675_));
 MUX2_X1 _38309_ (.A(\core.keymem.key_mem[3][109] ),
    .B(_14545_),
    .S(_14675_),
    .Z(_01871_));
 MUX2_X1 _38310_ (.A(\core.keymem.key_mem[3][10] ),
    .B(_14548_),
    .S(_14675_),
    .Z(_01872_));
 MUX2_X1 _38311_ (.A(\core.keymem.key_mem[3][110] ),
    .B(_12859_),
    .S(_14675_),
    .Z(_01873_));
 MUX2_X1 _38312_ (.A(\core.keymem.key_mem[3][111] ),
    .B(_12017_),
    .S(_14675_),
    .Z(_01874_));
 MUX2_X1 _38313_ (.A(\core.keymem.key_mem[3][112] ),
    .B(_12031_),
    .S(_14675_),
    .Z(_01875_));
 NAND2_X1 _38314_ (.A1(\core.keymem.key_mem[3][113] ),
    .A2(_14672_),
    .ZN(_14676_));
 BUF_X4 _38315_ (.A(_14668_),
    .Z(_14677_));
 NAND2_X1 _38316_ (.A1(_14236_),
    .A2(_14677_),
    .ZN(_14678_));
 OAI21_X1 _38317_ (.A(_14676_),
    .B1(_14678_),
    .B2(_14239_),
    .ZN(_01876_));
 MUX2_X1 _38318_ (.A(\core.keymem.key_mem[3][114] ),
    .B(_12869_),
    .S(_14675_),
    .Z(_01877_));
 MUX2_X1 _38319_ (.A(\core.keymem.key_mem[3][115] ),
    .B(_12059_),
    .S(_14675_),
    .Z(_01878_));
 MUX2_X1 _38320_ (.A(\core.keymem.key_mem[3][116] ),
    .B(_12077_),
    .S(_14675_),
    .Z(_01879_));
 BUF_X4 _38321_ (.A(_14671_),
    .Z(_14679_));
 NAND2_X1 _38322_ (.A1(\core.keymem.key_mem[3][117] ),
    .A2(_14679_),
    .ZN(_14680_));
 NAND2_X1 _38323_ (.A1(_14243_),
    .A2(_14677_),
    .ZN(_14681_));
 OAI21_X1 _38324_ (.A(_14680_),
    .B1(_14681_),
    .B2(_14246_),
    .ZN(_01880_));
 NAND2_X1 _38325_ (.A1(\core.keymem.key_mem[3][118] ),
    .A2(_14679_),
    .ZN(_14682_));
 OAI21_X1 _38326_ (.A(_14682_),
    .B1(_14674_),
    .B2(_14249_),
    .ZN(_01881_));
 MUX2_X1 _38327_ (.A(\core.keymem.key_mem[3][119] ),
    .B(_12096_),
    .S(_14675_),
    .Z(_01882_));
 NAND2_X1 _38328_ (.A1(\core.keymem.key_mem[3][11] ),
    .A2(_14679_),
    .ZN(_14683_));
 OAI21_X1 _38329_ (.A(_14683_),
    .B1(_14674_),
    .B2(_14255_),
    .ZN(_01883_));
 MUX2_X1 _38330_ (.A(\core.keymem.key_mem[3][120] ),
    .B(_12124_),
    .S(_14675_),
    .Z(_01884_));
 BUF_X8 _38331_ (.A(_14668_),
    .Z(_14684_));
 MUX2_X1 _38332_ (.A(\core.keymem.key_mem[3][121] ),
    .B(_12160_),
    .S(_14684_),
    .Z(_01885_));
 MUX2_X1 _38333_ (.A(\core.keymem.key_mem[3][122] ),
    .B(_12903_),
    .S(_14684_),
    .Z(_01886_));
 NAND2_X1 _38334_ (.A1(\core.keymem.key_mem[3][123] ),
    .A2(_14679_),
    .ZN(_14685_));
 OAI21_X1 _38335_ (.A(_14685_),
    .B1(_14674_),
    .B2(_12182_),
    .ZN(_01887_));
 NAND2_X1 _38336_ (.A1(\core.keymem.key_mem[3][124] ),
    .A2(_14679_),
    .ZN(_14686_));
 OAI21_X1 _38337_ (.A(_14686_),
    .B1(_14674_),
    .B2(_12926_),
    .ZN(_01888_));
 MUX2_X1 _38338_ (.A(\core.keymem.key_mem[3][125] ),
    .B(_12932_),
    .S(_14684_),
    .Z(_01889_));
 NAND2_X1 _38339_ (.A1(\core.keymem.key_mem[3][126] ),
    .A2(_14679_),
    .ZN(_14687_));
 OAI21_X1 _38340_ (.A(_14687_),
    .B1(_14674_),
    .B2(_12207_),
    .ZN(_01890_));
 MUX2_X1 _38341_ (.A(\core.keymem.key_mem[3][127] ),
    .B(_12945_),
    .S(_14684_),
    .Z(_01891_));
 NAND2_X1 _38342_ (.A1(\core.keymem.key_mem[3][12] ),
    .A2(_14679_),
    .ZN(_14688_));
 OAI21_X1 _38343_ (.A(_14688_),
    .B1(_14674_),
    .B2(_14281_),
    .ZN(_01892_));
 NAND2_X1 _38344_ (.A1(\core.keymem.key_mem[3][13] ),
    .A2(_14671_),
    .ZN(_14689_));
 NAND2_X1 _38345_ (.A1(_14226_),
    .A2(_14669_),
    .ZN(_14690_));
 OAI221_X1 _38346_ (.A(_14689_),
    .B1(_14671_),
    .B2(_14283_),
    .C1(_14290_),
    .C2(_14690_),
    .ZN(_01893_));
 MUX2_X1 _38347_ (.A(\core.keymem.key_mem[3][14] ),
    .B(_14574_),
    .S(_14684_),
    .Z(_01894_));
 MUX2_X1 _38348_ (.A(\core.keymem.key_mem[3][15] ),
    .B(_14306_),
    .S(_14684_),
    .Z(_01895_));
 MUX2_X1 _38349_ (.A(\core.keymem.key_mem[3][16] ),
    .B(_14575_),
    .S(_14684_),
    .Z(_01896_));
 NAND2_X1 _38350_ (.A1(\core.keymem.key_mem[3][17] ),
    .A2(_14679_),
    .ZN(_14691_));
 OAI21_X1 _38351_ (.A(_14691_),
    .B1(_14674_),
    .B2(_14314_),
    .ZN(_01897_));
 MUX2_X1 _38352_ (.A(\core.keymem.key_mem[3][18] ),
    .B(_14577_),
    .S(_14684_),
    .Z(_01898_));
 NAND2_X1 _38353_ (.A1(\core.keymem.key_mem[3][19] ),
    .A2(_14679_),
    .ZN(_14692_));
 OAI21_X1 _38354_ (.A(_14692_),
    .B1(_14674_),
    .B2(_14322_),
    .ZN(_01899_));
 MUX2_X1 _38355_ (.A(\core.keymem.key_mem[3][1] ),
    .B(_14324_),
    .S(_14684_),
    .Z(_01900_));
 MUX2_X1 _38356_ (.A(\core.keymem.key_mem[3][20] ),
    .B(_14326_),
    .S(_14684_),
    .Z(_01901_));
 BUF_X8 _38357_ (.A(_14668_),
    .Z(_14693_));
 MUX2_X1 _38358_ (.A(\core.keymem.key_mem[3][21] ),
    .B(_14579_),
    .S(_14693_),
    .Z(_01902_));
 MUX2_X1 _38359_ (.A(\core.keymem.key_mem[3][22] ),
    .B(_14580_),
    .S(_14693_),
    .Z(_01903_));
 NAND2_X1 _38360_ (.A1(\core.keymem.key_mem[3][23] ),
    .A2(_14679_),
    .ZN(_14694_));
 OAI21_X1 _38361_ (.A(_14694_),
    .B1(_14674_),
    .B2(_12272_),
    .ZN(_01904_));
 BUF_X4 _38362_ (.A(_14670_),
    .Z(_14695_));
 NAND2_X1 _38363_ (.A1(\core.keymem.key_mem[3][24] ),
    .A2(_14695_),
    .ZN(_14696_));
 BUF_X4 _38364_ (.A(_14671_),
    .Z(_14697_));
 OAI21_X1 _38365_ (.A(_14696_),
    .B1(_14697_),
    .B2(_13212_),
    .ZN(_01905_));
 MUX2_X1 _38366_ (.A(\core.keymem.key_mem[3][25] ),
    .B(_14585_),
    .S(_14693_),
    .Z(_01906_));
 MUX2_X1 _38367_ (.A(\core.keymem.key_mem[3][26] ),
    .B(_13241_),
    .S(_14693_),
    .Z(_01907_));
 MUX2_X1 _38368_ (.A(\core.keymem.key_mem[3][27] ),
    .B(_13284_),
    .S(_14693_),
    .Z(_01908_));
 MUX2_X1 _38369_ (.A(\core.keymem.key_mem[3][28] ),
    .B(_13325_),
    .S(_14693_),
    .Z(_01909_));
 MUX2_X1 _38370_ (.A(\core.keymem.key_mem[3][29] ),
    .B(_13329_),
    .S(_14693_),
    .Z(_01910_));
 NAND2_X1 _38371_ (.A1(\core.keymem.key_mem[3][2] ),
    .A2(_14695_),
    .ZN(_14698_));
 OAI21_X1 _38372_ (.A(_14698_),
    .B1(_14697_),
    .B2(_12337_),
    .ZN(_01911_));
 MUX2_X1 _38373_ (.A(\core.keymem.key_mem[3][30] ),
    .B(_13379_),
    .S(_14693_),
    .Z(_01912_));
 MUX2_X1 _38374_ (.A(\core.keymem.key_mem[3][31] ),
    .B(_13395_),
    .S(_14693_),
    .Z(_01913_));
 MUX2_X1 _38375_ (.A(\core.keymem.key_mem[3][32] ),
    .B(_13396_),
    .S(_14693_),
    .Z(_01914_));
 BUF_X4 _38376_ (.A(_14668_),
    .Z(_14699_));
 MUX2_X1 _38377_ (.A(\core.keymem.key_mem[3][33] ),
    .B(_13402_),
    .S(_14699_),
    .Z(_01915_));
 MUX2_X1 _38378_ (.A(\core.keymem.key_mem[3][34] ),
    .B(_13403_),
    .S(_14699_),
    .Z(_01916_));
 MUX2_X1 _38379_ (.A(\core.keymem.key_mem[3][35] ),
    .B(_13405_),
    .S(_14699_),
    .Z(_01917_));
 NAND2_X1 _38380_ (.A1(\core.keymem.key_mem[3][36] ),
    .A2(_14695_),
    .ZN(_14700_));
 OAI21_X1 _38381_ (.A(_14700_),
    .B1(_14697_),
    .B2(_13407_),
    .ZN(_01918_));
 NAND2_X1 _38382_ (.A1(\core.keymem.key_mem[3][37] ),
    .A2(_14695_),
    .ZN(_14701_));
 OAI21_X1 _38383_ (.A(_14701_),
    .B1(_14697_),
    .B2(_12439_),
    .ZN(_01919_));
 MUX2_X1 _38384_ (.A(\core.keymem.key_mem[3][38] ),
    .B(_13410_),
    .S(_14699_),
    .Z(_01920_));
 INV_X1 _38385_ (.A(\core.keymem.key_mem[3][39] ),
    .ZN(_14702_));
 NAND2_X1 _38386_ (.A1(_14360_),
    .A2(_14677_),
    .ZN(_14703_));
 OAI22_X1 _38387_ (.A1(_14702_),
    .A2(_14677_),
    .B1(_14703_),
    .B2(_13434_),
    .ZN(_01921_));
 MUX2_X1 _38388_ (.A(\core.keymem.key_mem[3][3] ),
    .B(_14370_),
    .S(_14699_),
    .Z(_01922_));
 NAND2_X1 _38389_ (.A1(\core.keymem.key_mem[3][40] ),
    .A2(_14695_),
    .ZN(_14704_));
 NAND2_X1 _38390_ (.A1(_14372_),
    .A2(_14677_),
    .ZN(_14705_));
 OAI21_X1 _38391_ (.A(_14704_),
    .B1(_14705_),
    .B2(_13457_),
    .ZN(_01923_));
 MUX2_X1 _38392_ (.A(\core.keymem.key_mem[3][41] ),
    .B(_13467_),
    .S(_14699_),
    .Z(_01924_));
 NAND2_X1 _38393_ (.A1(\core.keymem.key_mem[3][42] ),
    .A2(_14695_),
    .ZN(_14706_));
 OAI21_X1 _38394_ (.A(_14706_),
    .B1(_14697_),
    .B2(_14378_),
    .ZN(_01925_));
 MUX2_X1 _38395_ (.A(\core.keymem.key_mem[3][43] ),
    .B(_14596_),
    .S(_14699_),
    .Z(_01926_));
 MUX2_X1 _38396_ (.A(\core.keymem.key_mem[3][44] ),
    .B(_13497_),
    .S(_14699_),
    .Z(_01927_));
 NAND2_X1 _38397_ (.A1(\core.keymem.key_mem[3][45] ),
    .A2(_14695_),
    .ZN(_14707_));
 OAI21_X1 _38398_ (.A(_14707_),
    .B1(_14697_),
    .B2(_14598_),
    .ZN(_01928_));
 MUX2_X1 _38399_ (.A(\core.keymem.key_mem[3][46] ),
    .B(_14599_),
    .S(_14699_),
    .Z(_01929_));
 NAND2_X1 _38400_ (.A1(\core.keymem.key_mem[3][47] ),
    .A2(_14695_),
    .ZN(_14708_));
 OAI21_X1 _38401_ (.A(_14708_),
    .B1(_14697_),
    .B2(_12520_),
    .ZN(_01930_));
 NAND2_X1 _38402_ (.A1(\core.keymem.key_mem[3][48] ),
    .A2(_14695_),
    .ZN(_14709_));
 OAI21_X1 _38403_ (.A(_14709_),
    .B1(_14697_),
    .B2(_12532_),
    .ZN(_01931_));
 NAND2_X1 _38404_ (.A1(\core.keymem.key_mem[3][49] ),
    .A2(_14695_),
    .ZN(_14710_));
 NAND2_X1 _38405_ (.A1(_14392_),
    .A2(_14677_),
    .ZN(_14711_));
 OAI21_X1 _38406_ (.A(_14710_),
    .B1(_14711_),
    .B2(_13529_),
    .ZN(_01932_));
 MUX2_X1 _38407_ (.A(\core.keymem.key_mem[3][4] ),
    .B(_14604_),
    .S(_14699_),
    .Z(_01933_));
 BUF_X4 _38408_ (.A(_14670_),
    .Z(_14712_));
 NAND2_X1 _38409_ (.A1(\core.keymem.key_mem[3][50] ),
    .A2(_14712_),
    .ZN(_14713_));
 OAI21_X1 _38410_ (.A(_14713_),
    .B1(_14697_),
    .B2(_14402_),
    .ZN(_01934_));
 BUF_X4 _38411_ (.A(_14668_),
    .Z(_14714_));
 MUX2_X1 _38412_ (.A(\core.keymem.key_mem[3][51] ),
    .B(_13564_),
    .S(_14714_),
    .Z(_01935_));
 NAND2_X1 _38413_ (.A1(\core.keymem.key_mem[3][52] ),
    .A2(_14712_),
    .ZN(_14715_));
 OAI21_X1 _38414_ (.A(_14715_),
    .B1(_14697_),
    .B2(_12568_),
    .ZN(_01936_));
 NAND2_X1 _38415_ (.A1(\core.keymem.key_mem[3][53] ),
    .A2(_14712_),
    .ZN(_14716_));
 BUF_X4 _38416_ (.A(_14671_),
    .Z(_14717_));
 OAI21_X1 _38417_ (.A(_14716_),
    .B1(_14717_),
    .B2(_12584_),
    .ZN(_01937_));
 NAND2_X1 _38418_ (.A1(\core.keymem.key_mem[3][54] ),
    .A2(_14712_),
    .ZN(_14718_));
 OAI21_X1 _38419_ (.A(_14718_),
    .B1(_14717_),
    .B2(_13575_),
    .ZN(_01938_));
 NAND2_X1 _38420_ (.A1(\core.keymem.key_mem[3][55] ),
    .A2(_14712_),
    .ZN(_14719_));
 OAI21_X1 _38421_ (.A(_14719_),
    .B1(_14717_),
    .B2(_14612_),
    .ZN(_01939_));
 MUX2_X1 _38422_ (.A(\core.keymem.key_mem[3][56] ),
    .B(_14613_),
    .S(_14714_),
    .Z(_01940_));
 MUX2_X1 _38423_ (.A(\core.keymem.key_mem[3][57] ),
    .B(_14615_),
    .S(_14714_),
    .Z(_01941_));
 MUX2_X1 _38424_ (.A(\core.keymem.key_mem[3][58] ),
    .B(_14616_),
    .S(_14714_),
    .Z(_01942_));
 NAND2_X1 _38425_ (.A1(\core.keymem.key_mem[3][59] ),
    .A2(_14712_),
    .ZN(_14720_));
 OAI21_X1 _38426_ (.A(_14720_),
    .B1(_14717_),
    .B2(_14424_),
    .ZN(_01943_));
 MUX2_X1 _38427_ (.A(\core.keymem.key_mem[3][5] ),
    .B(_12606_),
    .S(_14714_),
    .Z(_01944_));
 NAND2_X1 _38428_ (.A1(\core.keymem.key_mem[3][60] ),
    .A2(_14712_),
    .ZN(_14721_));
 OAI21_X1 _38429_ (.A(_14721_),
    .B1(_14717_),
    .B2(_14619_),
    .ZN(_01945_));
 INV_X1 _38430_ (.A(\core.keymem.key_mem[3][61] ),
    .ZN(_14722_));
 NAND2_X1 _38431_ (.A1(_14432_),
    .A2(_14677_),
    .ZN(_14723_));
 OAI22_X1 _38432_ (.A1(_14722_),
    .A2(_14677_),
    .B1(_14723_),
    .B2(_14434_),
    .ZN(_01946_));
 MUX2_X1 _38433_ (.A(\core.keymem.key_mem[3][62] ),
    .B(_13637_),
    .S(_14714_),
    .Z(_01947_));
 MUX2_X1 _38434_ (.A(\core.keymem.key_mem[3][63] ),
    .B(_14622_),
    .S(_14714_),
    .Z(_01948_));
 MUX2_X1 _38435_ (.A(\core.keymem.key_mem[3][64] ),
    .B(_12622_),
    .S(_14714_),
    .Z(_01949_));
 NAND2_X1 _38436_ (.A1(\core.keymem.key_mem[3][65] ),
    .A2(_14712_),
    .ZN(_14724_));
 OAI21_X1 _38437_ (.A(_14724_),
    .B1(_14717_),
    .B2(_13673_),
    .ZN(_01950_));
 MUX2_X1 _38438_ (.A(\core.keymem.key_mem[3][66] ),
    .B(_13681_),
    .S(_14714_),
    .Z(_01951_));
 NAND2_X1 _38439_ (.A1(\core.keymem.key_mem[3][67] ),
    .A2(_14712_),
    .ZN(_14725_));
 OAI21_X1 _38440_ (.A(_14725_),
    .B1(_14717_),
    .B2(_13690_),
    .ZN(_01952_));
 NAND2_X1 _38441_ (.A1(\core.keymem.key_mem[3][68] ),
    .A2(_14712_),
    .ZN(_14726_));
 OAI21_X1 _38442_ (.A(_14726_),
    .B1(_14717_),
    .B2(_12635_),
    .ZN(_01953_));
 BUF_X4 _38443_ (.A(_14670_),
    .Z(_14727_));
 NAND2_X1 _38444_ (.A1(\core.keymem.key_mem[3][69] ),
    .A2(_14727_),
    .ZN(_14728_));
 OAI21_X1 _38445_ (.A(_14728_),
    .B1(_14717_),
    .B2(_13700_),
    .ZN(_01954_));
 MUX2_X1 _38446_ (.A(\core.keymem.key_mem[3][6] ),
    .B(_13711_),
    .S(_14714_),
    .Z(_01955_));
 BUF_X8 _38447_ (.A(_14668_),
    .Z(_14729_));
 MUX2_X1 _38448_ (.A(\core.keymem.key_mem[3][70] ),
    .B(_13713_),
    .S(_14729_),
    .Z(_01956_));
 NAND2_X1 _38449_ (.A1(\core.keymem.key_mem[3][71] ),
    .A2(_14727_),
    .ZN(_14730_));
 OAI21_X1 _38450_ (.A(_14730_),
    .B1(_14717_),
    .B2(_12659_),
    .ZN(_01957_));
 NAND2_X1 _38451_ (.A1(\core.keymem.key_mem[3][72] ),
    .A2(_14727_),
    .ZN(_14731_));
 BUF_X4 _38452_ (.A(_14671_),
    .Z(_14732_));
 OAI21_X1 _38453_ (.A(_14731_),
    .B1(_14732_),
    .B2(_13716_),
    .ZN(_01958_));
 NAND2_X1 _38454_ (.A1(\core.keymem.key_mem[3][73] ),
    .A2(_14727_),
    .ZN(_14733_));
 OAI21_X1 _38455_ (.A(_14733_),
    .B1(_14732_),
    .B2(_12688_),
    .ZN(_01959_));
 MUX2_X1 _38456_ (.A(\core.keymem.key_mem[3][74] ),
    .B(_14636_),
    .S(_14729_),
    .Z(_01960_));
 NAND2_X1 _38457_ (.A1(\core.keymem.key_mem[3][75] ),
    .A2(_14727_),
    .ZN(_14734_));
 OAI21_X1 _38458_ (.A(_14734_),
    .B1(_14732_),
    .B2(_13733_),
    .ZN(_01961_));
 MUX2_X1 _38459_ (.A(\core.keymem.key_mem[3][76] ),
    .B(_13741_),
    .S(_14729_),
    .Z(_01962_));
 MUX2_X1 _38460_ (.A(\core.keymem.key_mem[3][77] ),
    .B(_14639_),
    .S(_14729_),
    .Z(_01963_));
 NAND2_X1 _38461_ (.A1(\core.keymem.key_mem[3][78] ),
    .A2(_14727_),
    .ZN(_14735_));
 OAI21_X1 _38462_ (.A(_14735_),
    .B1(_14732_),
    .B2(_12708_),
    .ZN(_01964_));
 NAND2_X1 _38463_ (.A1(\core.keymem.key_mem[3][79] ),
    .A2(_14727_),
    .ZN(_14736_));
 OAI21_X1 _38464_ (.A(_14736_),
    .B1(_14732_),
    .B2(_14476_),
    .ZN(_01965_));
 NAND2_X1 _38465_ (.A1(\core.keymem.key_mem[3][7] ),
    .A2(_14727_),
    .ZN(_14737_));
 OAI21_X1 _38466_ (.A(_14737_),
    .B1(_14732_),
    .B2(_13767_),
    .ZN(_01966_));
 MUX2_X1 _38467_ (.A(\core.keymem.key_mem[3][80] ),
    .B(_13769_),
    .S(_14729_),
    .Z(_01967_));
 NAND2_X1 _38468_ (.A1(\core.keymem.key_mem[3][81] ),
    .A2(_14727_),
    .ZN(_14738_));
 OAI21_X1 _38469_ (.A(_14738_),
    .B1(_14732_),
    .B2(_13775_),
    .ZN(_01968_));
 NAND2_X1 _38470_ (.A1(\core.keymem.key_mem[3][82] ),
    .A2(_14727_),
    .ZN(_14739_));
 OAI21_X1 _38471_ (.A(_14739_),
    .B1(_14732_),
    .B2(_13783_),
    .ZN(_01969_));
 BUF_X4 _38472_ (.A(_14670_),
    .Z(_14740_));
 NAND2_X1 _38473_ (.A1(\core.keymem.key_mem[3][83] ),
    .A2(_14740_),
    .ZN(_14741_));
 OAI21_X1 _38474_ (.A(_14741_),
    .B1(_14732_),
    .B2(_13791_),
    .ZN(_01970_));
 NAND2_X1 _38475_ (.A1(\core.keymem.key_mem[3][84] ),
    .A2(_14740_),
    .ZN(_14742_));
 OAI21_X1 _38476_ (.A(_14742_),
    .B1(_14732_),
    .B2(_12725_),
    .ZN(_01971_));
 NAND2_X1 _38477_ (.A1(\core.keymem.key_mem[3][85] ),
    .A2(_14740_),
    .ZN(_14743_));
 OAI21_X1 _38478_ (.A(_14743_),
    .B1(_14672_),
    .B2(_14484_),
    .ZN(_01972_));
 MUX2_X1 _38479_ (.A(\core.keymem.key_mem[3][86] ),
    .B(_12741_),
    .S(_14729_),
    .Z(_01973_));
 NAND2_X1 _38480_ (.A1(\core.keymem.key_mem[3][87] ),
    .A2(_14740_),
    .ZN(_14744_));
 OAI21_X1 _38481_ (.A(_14744_),
    .B1(_14672_),
    .B2(_14489_),
    .ZN(_01974_));
 MUX2_X1 _38482_ (.A(\core.keymem.key_mem[3][88] ),
    .B(_14650_),
    .S(_14729_),
    .Z(_01975_));
 NAND2_X1 _38483_ (.A1(\core.keymem.key_mem[3][89] ),
    .A2(_14740_),
    .ZN(_14745_));
 OAI21_X1 _38484_ (.A(_14745_),
    .B1(_14672_),
    .B2(_14652_),
    .ZN(_01976_));
 NAND2_X1 _38485_ (.A1(\core.keymem.key_mem[3][8] ),
    .A2(_14740_),
    .ZN(_14746_));
 NAND2_X1 _38486_ (.A1(_14497_),
    .A2(_14677_),
    .ZN(_14747_));
 OAI21_X1 _38487_ (.A(_14746_),
    .B1(_14747_),
    .B2(_14504_),
    .ZN(_01977_));
 MUX2_X1 _38488_ (.A(\core.keymem.key_mem[3][90] ),
    .B(_14655_),
    .S(_14729_),
    .Z(_01978_));
 NAND2_X1 _38489_ (.A1(\core.keymem.key_mem[3][91] ),
    .A2(_14740_),
    .ZN(_14748_));
 OAI21_X1 _38490_ (.A(_14748_),
    .B1(_14672_),
    .B2(_14510_),
    .ZN(_01979_));
 NAND2_X1 _38491_ (.A1(\core.keymem.key_mem[3][92] ),
    .A2(_14740_),
    .ZN(_14749_));
 OAI21_X1 _38492_ (.A(_14749_),
    .B1(_14672_),
    .B2(_14512_),
    .ZN(_01980_));
 NAND2_X1 _38493_ (.A1(\core.keymem.key_mem[3][93] ),
    .A2(_14740_),
    .ZN(_14750_));
 NAND2_X1 _38494_ (.A1(_14514_),
    .A2(_14677_),
    .ZN(_14751_));
 OAI21_X1 _38495_ (.A(_14750_),
    .B1(_14751_),
    .B2(_14520_),
    .ZN(_01981_));
 MUX2_X1 _38496_ (.A(\core.keymem.key_mem[3][94] ),
    .B(_14660_),
    .S(_14729_),
    .Z(_01982_));
 MUX2_X1 _38497_ (.A(\core.keymem.key_mem[3][95] ),
    .B(_14661_),
    .S(_14729_),
    .Z(_01983_));
 NAND2_X1 _38498_ (.A1(\core.keymem.key_mem[3][96] ),
    .A2(_14740_),
    .ZN(_14752_));
 OAI21_X1 _38499_ (.A(_14752_),
    .B1(_14672_),
    .B2(_14663_),
    .ZN(_01984_));
 NAND2_X1 _38500_ (.A1(\core.keymem.key_mem[3][97] ),
    .A2(_14671_),
    .ZN(_14753_));
 OAI21_X1 _38501_ (.A(_14753_),
    .B1(_14672_),
    .B2(_12777_),
    .ZN(_01985_));
 NAND2_X1 _38502_ (.A1(\core.keymem.key_mem[3][98] ),
    .A2(_14671_),
    .ZN(_14754_));
 OAI21_X1 _38503_ (.A(_14754_),
    .B1(_14672_),
    .B2(_13910_),
    .ZN(_01986_));
 MUX2_X1 _38504_ (.A(\core.keymem.key_mem[3][99] ),
    .B(_12800_),
    .S(_14668_),
    .Z(_01987_));
 MUX2_X1 _38505_ (.A(\core.keymem.key_mem[3][9] ),
    .B(_14666_),
    .S(_14668_),
    .Z(_01988_));
 OR2_X1 _38506_ (.A1(_11794_),
    .A2(_12802_),
    .ZN(_14755_));
 BUF_X4 _38507_ (.A(_14755_),
    .Z(_14756_));
 NOR2_X4 _38508_ (.A1(_13989_),
    .A2(_14756_),
    .ZN(_14757_));
 BUF_X4 _38509_ (.A(_14757_),
    .Z(_14758_));
 BUF_X4 _38510_ (.A(_14758_),
    .Z(_14759_));
 MUX2_X1 _38511_ (.A(\core.keymem.key_mem[4][0] ),
    .B(_11844_),
    .S(_14759_),
    .Z(_01989_));
 MUX2_X1 _38512_ (.A(\core.keymem.key_mem[4][100] ),
    .B(_11873_),
    .S(_14759_),
    .Z(_01990_));
 MUX2_X1 _38513_ (.A(\core.keymem.key_mem[4][101] ),
    .B(_12813_),
    .S(_14759_),
    .Z(_01991_));
 MUX2_X1 _38514_ (.A(\core.keymem.key_mem[4][102] ),
    .B(_11906_),
    .S(_14759_),
    .Z(_01992_));
 MUX2_X1 _38515_ (.A(\core.keymem.key_mem[4][103] ),
    .B(_11929_),
    .S(_14759_),
    .Z(_01993_));
 OR2_X1 _38516_ (.A1(_13989_),
    .A2(_14756_),
    .ZN(_14760_));
 CLKBUF_X3 _38517_ (.A(_14760_),
    .Z(_14761_));
 BUF_X4 _38518_ (.A(_14761_),
    .Z(_14762_));
 NAND2_X1 _38519_ (.A1(\core.keymem.key_mem[4][104] ),
    .A2(_14762_),
    .ZN(_14763_));
 BUF_X4 _38520_ (.A(_14761_),
    .Z(_14764_));
 BUF_X4 _38521_ (.A(_14764_),
    .Z(_14765_));
 OAI21_X1 _38522_ (.A(_14763_),
    .B1(_14765_),
    .B2(_12822_),
    .ZN(_01994_));
 MUX2_X1 _38523_ (.A(\core.keymem.key_mem[4][105] ),
    .B(_12830_),
    .S(_14759_),
    .Z(_01995_));
 BUF_X4 _38524_ (.A(_14758_),
    .Z(_14766_));
 MUX2_X1 _38525_ (.A(\core.keymem.key_mem[4][106] ),
    .B(_12832_),
    .S(_14766_),
    .Z(_01996_));
 MUX2_X1 _38526_ (.A(\core.keymem.key_mem[4][107] ),
    .B(_11967_),
    .S(_14766_),
    .Z(_01997_));
 MUX2_X1 _38527_ (.A(\core.keymem.key_mem[4][108] ),
    .B(_11981_),
    .S(_14766_),
    .Z(_01998_));
 MUX2_X1 _38528_ (.A(\core.keymem.key_mem[4][109] ),
    .B(_12842_),
    .S(_14766_),
    .Z(_01999_));
 NAND2_X1 _38529_ (.A1(\core.keymem.key_mem[4][10] ),
    .A2(_14762_),
    .ZN(_14767_));
 OAI21_X1 _38530_ (.A(_14767_),
    .B1(_14765_),
    .B2(_12858_),
    .ZN(_02000_));
 MUX2_X1 _38531_ (.A(\core.keymem.key_mem[4][110] ),
    .B(_12859_),
    .S(_14766_),
    .Z(_02001_));
 MUX2_X1 _38532_ (.A(\core.keymem.key_mem[4][111] ),
    .B(_12017_),
    .S(_14766_),
    .Z(_02002_));
 MUX2_X1 _38533_ (.A(\core.keymem.key_mem[4][112] ),
    .B(_12031_),
    .S(_14766_),
    .Z(_02003_));
 MUX2_X1 _38534_ (.A(\core.keymem.key_mem[4][113] ),
    .B(_12868_),
    .S(_14766_),
    .Z(_02004_));
 MUX2_X1 _38535_ (.A(\core.keymem.key_mem[4][114] ),
    .B(_12869_),
    .S(_14766_),
    .Z(_02005_));
 MUX2_X1 _38536_ (.A(\core.keymem.key_mem[4][115] ),
    .B(_12059_),
    .S(_14766_),
    .Z(_02006_));
 BUF_X4 _38537_ (.A(_14758_),
    .Z(_14768_));
 MUX2_X1 _38538_ (.A(\core.keymem.key_mem[4][116] ),
    .B(_12077_),
    .S(_14768_),
    .Z(_02007_));
 MUX2_X1 _38539_ (.A(\core.keymem.key_mem[4][117] ),
    .B(_12877_),
    .S(_14768_),
    .Z(_02008_));
 MUX2_X1 _38540_ (.A(\core.keymem.key_mem[4][118] ),
    .B(_12882_),
    .S(_14768_),
    .Z(_02009_));
 MUX2_X1 _38541_ (.A(\core.keymem.key_mem[4][119] ),
    .B(_12096_),
    .S(_14768_),
    .Z(_02010_));
 NAND2_X1 _38542_ (.A1(\core.keymem.key_mem[4][11] ),
    .A2(_14762_),
    .ZN(_14769_));
 OAI21_X1 _38543_ (.A(_14769_),
    .B1(_14765_),
    .B2(_12895_),
    .ZN(_02011_));
 MUX2_X1 _38544_ (.A(\core.keymem.key_mem[4][120] ),
    .B(_12124_),
    .S(_14768_),
    .Z(_02012_));
 MUX2_X1 _38545_ (.A(\core.keymem.key_mem[4][121] ),
    .B(_12160_),
    .S(_14768_),
    .Z(_02013_));
 MUX2_X1 _38546_ (.A(\core.keymem.key_mem[4][122] ),
    .B(_12903_),
    .S(_14768_),
    .Z(_02014_));
 NAND2_X1 _38547_ (.A1(\core.keymem.key_mem[4][123] ),
    .A2(_14762_),
    .ZN(_14770_));
 OAI21_X1 _38548_ (.A(_14770_),
    .B1(_14765_),
    .B2(_12182_),
    .ZN(_02015_));
 NAND2_X1 _38549_ (.A1(\core.keymem.key_mem[4][124] ),
    .A2(_14762_),
    .ZN(_14771_));
 OAI21_X1 _38550_ (.A(_14771_),
    .B1(_14765_),
    .B2(_12926_),
    .ZN(_02016_));
 MUX2_X1 _38551_ (.A(\core.keymem.key_mem[4][125] ),
    .B(_12932_),
    .S(_14768_),
    .Z(_02017_));
 NAND2_X1 _38552_ (.A1(\core.keymem.key_mem[4][126] ),
    .A2(_14762_),
    .ZN(_14772_));
 OAI21_X1 _38553_ (.A(_14772_),
    .B1(_14765_),
    .B2(_12207_),
    .ZN(_02018_));
 MUX2_X1 _38554_ (.A(\core.keymem.key_mem[4][127] ),
    .B(_12945_),
    .S(_14768_),
    .Z(_02019_));
 MUX2_X1 _38555_ (.A(\core.keymem.key_mem[4][12] ),
    .B(_12958_),
    .S(_14768_),
    .Z(_02020_));
 BUF_X4 _38556_ (.A(_14757_),
    .Z(_14773_));
 MUX2_X1 _38557_ (.A(\core.keymem.key_mem[4][13] ),
    .B(_12974_),
    .S(_14773_),
    .Z(_02021_));
 NOR2_X1 _38558_ (.A1(\core.keymem.key_mem[4][14] ),
    .A2(_14759_),
    .ZN(_14774_));
 AOI21_X1 _38559_ (.A(_14774_),
    .B1(_14759_),
    .B2(_13007_),
    .ZN(_02022_));
 MUX2_X1 _38560_ (.A(\core.keymem.key_mem[4][15] ),
    .B(_13017_),
    .S(_14773_),
    .Z(_02023_));
 MUX2_X1 _38561_ (.A(\core.keymem.key_mem[4][16] ),
    .B(_13029_),
    .S(_14773_),
    .Z(_02024_));
 NAND2_X1 _38562_ (.A1(\core.keymem.key_mem[4][17] ),
    .A2(_14762_),
    .ZN(_14775_));
 OAI21_X1 _38563_ (.A(_14775_),
    .B1(_14765_),
    .B2(_13042_),
    .ZN(_02025_));
 MUX2_X1 _38564_ (.A(\core.keymem.key_mem[4][18] ),
    .B(_13094_),
    .S(_14773_),
    .Z(_02026_));
 BUF_X4 _38565_ (.A(_14761_),
    .Z(_14776_));
 NAND2_X1 _38566_ (.A1(\core.keymem.key_mem[4][19] ),
    .A2(_14776_),
    .ZN(_14777_));
 OAI21_X1 _38567_ (.A(_14777_),
    .B1(_14765_),
    .B2(_13109_),
    .ZN(_02027_));
 MUX2_X1 _38568_ (.A(\core.keymem.key_mem[4][1] ),
    .B(_13134_),
    .S(_14773_),
    .Z(_02028_));
 MUX2_X1 _38569_ (.A(\core.keymem.key_mem[4][20] ),
    .B(_13146_),
    .S(_14773_),
    .Z(_02029_));
 MUX2_X1 _38570_ (.A(\core.keymem.key_mem[4][21] ),
    .B(_13155_),
    .S(_14773_),
    .Z(_02030_));
 NOR2_X1 _38571_ (.A1(\core.keymem.key_mem[4][22] ),
    .A2(_14759_),
    .ZN(_14778_));
 AOI21_X1 _38572_ (.A(_14778_),
    .B1(_14759_),
    .B2(_13191_),
    .ZN(_02031_));
 MUX2_X1 _38573_ (.A(\core.keymem.key_mem[4][23] ),
    .B(_13196_),
    .S(_14773_),
    .Z(_02032_));
 NAND2_X1 _38574_ (.A1(\core.keymem.key_mem[4][24] ),
    .A2(_14776_),
    .ZN(_14779_));
 OAI21_X1 _38575_ (.A(_14779_),
    .B1(_14765_),
    .B2(_13212_),
    .ZN(_02033_));
 MUX2_X1 _38576_ (.A(\core.keymem.key_mem[4][25] ),
    .B(_13233_),
    .S(_14773_),
    .Z(_02034_));
 MUX2_X1 _38577_ (.A(\core.keymem.key_mem[4][26] ),
    .B(_13241_),
    .S(_14773_),
    .Z(_02035_));
 BUF_X4 _38578_ (.A(_14757_),
    .Z(_14780_));
 MUX2_X1 _38579_ (.A(\core.keymem.key_mem[4][27] ),
    .B(_13284_),
    .S(_14780_),
    .Z(_02036_));
 MUX2_X1 _38580_ (.A(\core.keymem.key_mem[4][28] ),
    .B(_13325_),
    .S(_14780_),
    .Z(_02037_));
 MUX2_X1 _38581_ (.A(\core.keymem.key_mem[4][29] ),
    .B(_13329_),
    .S(_14780_),
    .Z(_02038_));
 NAND2_X1 _38582_ (.A1(\core.keymem.key_mem[4][2] ),
    .A2(_14776_),
    .ZN(_14781_));
 OAI21_X1 _38583_ (.A(_14781_),
    .B1(_14765_),
    .B2(_13335_),
    .ZN(_02039_));
 MUX2_X1 _38584_ (.A(\core.keymem.key_mem[4][30] ),
    .B(_13379_),
    .S(_14780_),
    .Z(_02040_));
 MUX2_X1 _38585_ (.A(\core.keymem.key_mem[4][31] ),
    .B(_13395_),
    .S(_14780_),
    .Z(_02041_));
 MUX2_X1 _38586_ (.A(\core.keymem.key_mem[4][32] ),
    .B(_13396_),
    .S(_14780_),
    .Z(_02042_));
 MUX2_X1 _38587_ (.A(\core.keymem.key_mem[4][33] ),
    .B(_13402_),
    .S(_14780_),
    .Z(_02043_));
 MUX2_X1 _38588_ (.A(\core.keymem.key_mem[4][34] ),
    .B(_13403_),
    .S(_14780_),
    .Z(_02044_));
 MUX2_X1 _38589_ (.A(\core.keymem.key_mem[4][35] ),
    .B(_13405_),
    .S(_14780_),
    .Z(_02045_));
 NAND2_X1 _38590_ (.A1(\core.keymem.key_mem[4][36] ),
    .A2(_14776_),
    .ZN(_14782_));
 BUF_X4 _38591_ (.A(_14764_),
    .Z(_14783_));
 OAI21_X1 _38592_ (.A(_14782_),
    .B1(_14783_),
    .B2(_13407_),
    .ZN(_02046_));
 NAND2_X1 _38593_ (.A1(\core.keymem.key_mem[4][37] ),
    .A2(_14776_),
    .ZN(_14784_));
 OAI21_X1 _38594_ (.A(_14784_),
    .B1(_14783_),
    .B2(_12439_),
    .ZN(_02047_));
 MUX2_X1 _38595_ (.A(\core.keymem.key_mem[4][38] ),
    .B(_13410_),
    .S(_14780_),
    .Z(_02048_));
 NAND2_X1 _38596_ (.A1(\core.keymem.key_mem[4][39] ),
    .A2(_14776_),
    .ZN(_14785_));
 OAI21_X1 _38597_ (.A(_14785_),
    .B1(_14783_),
    .B2(_13435_),
    .ZN(_02049_));
 NAND2_X1 _38598_ (.A1(\core.keymem.key_mem[4][3] ),
    .A2(_14776_),
    .ZN(_14786_));
 OAI21_X1 _38599_ (.A(_14786_),
    .B1(_14783_),
    .B2(_13448_),
    .ZN(_02050_));
 NAND2_X1 _38600_ (.A1(\core.keymem.key_mem[4][40] ),
    .A2(_14776_),
    .ZN(_14787_));
 OAI21_X1 _38601_ (.A(_14787_),
    .B1(_14783_),
    .B2(_13457_),
    .ZN(_02051_));
 BUF_X4 _38602_ (.A(_14757_),
    .Z(_14788_));
 MUX2_X1 _38603_ (.A(\core.keymem.key_mem[4][41] ),
    .B(_13467_),
    .S(_14788_),
    .Z(_02052_));
 MUX2_X1 _38604_ (.A(\core.keymem.key_mem[4][42] ),
    .B(_13490_),
    .S(_14788_),
    .Z(_02053_));
 NAND2_X1 _38605_ (.A1(\core.keymem.key_mem[4][43] ),
    .A2(_14776_),
    .ZN(_14789_));
 OAI21_X1 _38606_ (.A(_14789_),
    .B1(_14783_),
    .B2(_13496_),
    .ZN(_02054_));
 MUX2_X1 _38607_ (.A(\core.keymem.key_mem[4][44] ),
    .B(_13497_),
    .S(_14788_),
    .Z(_02055_));
 NAND2_X1 _38608_ (.A1(\core.keymem.key_mem[4][45] ),
    .A2(_14776_),
    .ZN(_14790_));
 OAI21_X1 _38609_ (.A(_14790_),
    .B1(_14783_),
    .B2(_13510_),
    .ZN(_02056_));
 BUF_X4 _38610_ (.A(_14761_),
    .Z(_14791_));
 NAND2_X1 _38611_ (.A1(\core.keymem.key_mem[4][46] ),
    .A2(_14791_),
    .ZN(_14792_));
 OAI21_X1 _38612_ (.A(_14792_),
    .B1(_14783_),
    .B2(_13517_),
    .ZN(_02057_));
 NAND2_X1 _38613_ (.A1(\core.keymem.key_mem[4][47] ),
    .A2(_14791_),
    .ZN(_14793_));
 OAI21_X1 _38614_ (.A(_14793_),
    .B1(_14783_),
    .B2(_12520_),
    .ZN(_02058_));
 NAND2_X1 _38615_ (.A1(\core.keymem.key_mem[4][48] ),
    .A2(_14791_),
    .ZN(_14794_));
 OAI21_X1 _38616_ (.A(_14794_),
    .B1(_14783_),
    .B2(_12532_),
    .ZN(_02059_));
 NAND2_X1 _38617_ (.A1(\core.keymem.key_mem[4][49] ),
    .A2(_14791_),
    .ZN(_14795_));
 BUF_X4 _38618_ (.A(_14764_),
    .Z(_14796_));
 OAI21_X1 _38619_ (.A(_14795_),
    .B1(_14796_),
    .B2(_13529_),
    .ZN(_02060_));
 MUX2_X1 _38620_ (.A(\core.keymem.key_mem[4][4] ),
    .B(_13538_),
    .S(_14788_),
    .Z(_02061_));
 MUX2_X1 _38621_ (.A(\core.keymem.key_mem[4][50] ),
    .B(_13557_),
    .S(_14788_),
    .Z(_02062_));
 MUX2_X1 _38622_ (.A(\core.keymem.key_mem[4][51] ),
    .B(_13564_),
    .S(_14788_),
    .Z(_02063_));
 NAND2_X1 _38623_ (.A1(\core.keymem.key_mem[4][52] ),
    .A2(_14791_),
    .ZN(_14797_));
 OAI21_X1 _38624_ (.A(_14797_),
    .B1(_14796_),
    .B2(_12568_),
    .ZN(_02064_));
 NAND2_X1 _38625_ (.A1(\core.keymem.key_mem[4][53] ),
    .A2(_14791_),
    .ZN(_14798_));
 OAI21_X1 _38626_ (.A(_14798_),
    .B1(_14796_),
    .B2(_12584_),
    .ZN(_02065_));
 NAND2_X1 _38627_ (.A1(\core.keymem.key_mem[4][54] ),
    .A2(_14791_),
    .ZN(_14799_));
 OAI21_X1 _38628_ (.A(_14799_),
    .B1(_14796_),
    .B2(_13575_),
    .ZN(_02066_));
 MUX2_X1 _38629_ (.A(\core.keymem.key_mem[4][55] ),
    .B(_13581_),
    .S(_14788_),
    .Z(_02067_));
 MUX2_X1 _38630_ (.A(\core.keymem.key_mem[4][56] ),
    .B(_13589_),
    .S(_14788_),
    .Z(_02068_));
 MUX2_X1 _38631_ (.A(\core.keymem.key_mem[4][57] ),
    .B(_13604_),
    .S(_14788_),
    .Z(_02069_));
 MUX2_X1 _38632_ (.A(\core.keymem.key_mem[4][58] ),
    .B(_13611_),
    .S(_14788_),
    .Z(_02070_));
 BUF_X4 _38633_ (.A(_14757_),
    .Z(_14800_));
 MUX2_X1 _38634_ (.A(\core.keymem.key_mem[4][59] ),
    .B(_13616_),
    .S(_14800_),
    .Z(_02071_));
 MUX2_X1 _38635_ (.A(\core.keymem.key_mem[4][5] ),
    .B(_12606_),
    .S(_14800_),
    .Z(_02072_));
 MUX2_X1 _38636_ (.A(\core.keymem.key_mem[4][60] ),
    .B(_13622_),
    .S(_14800_),
    .Z(_02073_));
 MUX2_X1 _38637_ (.A(\core.keymem.key_mem[4][61] ),
    .B(_13632_),
    .S(_14800_),
    .Z(_02074_));
 MUX2_X1 _38638_ (.A(\core.keymem.key_mem[4][62] ),
    .B(_13637_),
    .S(_14800_),
    .Z(_02075_));
 MUX2_X1 _38639_ (.A(\core.keymem.key_mem[4][63] ),
    .B(_13659_),
    .S(_14800_),
    .Z(_02076_));
 MUX2_X1 _38640_ (.A(\core.keymem.key_mem[4][64] ),
    .B(_12622_),
    .S(_14800_),
    .Z(_02077_));
 NAND2_X1 _38641_ (.A1(\core.keymem.key_mem[4][65] ),
    .A2(_14791_),
    .ZN(_14801_));
 OAI21_X1 _38642_ (.A(_14801_),
    .B1(_14796_),
    .B2(_13673_),
    .ZN(_02078_));
 MUX2_X1 _38643_ (.A(\core.keymem.key_mem[4][66] ),
    .B(_13681_),
    .S(_14800_),
    .Z(_02079_));
 NAND2_X1 _38644_ (.A1(\core.keymem.key_mem[4][67] ),
    .A2(_14791_),
    .ZN(_14802_));
 OAI21_X1 _38645_ (.A(_14802_),
    .B1(_14796_),
    .B2(_13690_),
    .ZN(_02080_));
 NAND2_X1 _38646_ (.A1(\core.keymem.key_mem[4][68] ),
    .A2(_14791_),
    .ZN(_14803_));
 OAI21_X1 _38647_ (.A(_14803_),
    .B1(_14796_),
    .B2(_12635_),
    .ZN(_02081_));
 BUF_X4 _38648_ (.A(_14761_),
    .Z(_14804_));
 NAND2_X1 _38649_ (.A1(\core.keymem.key_mem[4][69] ),
    .A2(_14804_),
    .ZN(_14805_));
 OAI21_X1 _38650_ (.A(_14805_),
    .B1(_14796_),
    .B2(_13700_),
    .ZN(_02082_));
 MUX2_X1 _38651_ (.A(\core.keymem.key_mem[4][6] ),
    .B(_13711_),
    .S(_14800_),
    .Z(_02083_));
 MUX2_X1 _38652_ (.A(\core.keymem.key_mem[4][70] ),
    .B(_13713_),
    .S(_14800_),
    .Z(_02084_));
 NAND2_X1 _38653_ (.A1(\core.keymem.key_mem[4][71] ),
    .A2(_14804_),
    .ZN(_14806_));
 OAI21_X1 _38654_ (.A(_14806_),
    .B1(_14796_),
    .B2(_12659_),
    .ZN(_02085_));
 NAND2_X1 _38655_ (.A1(\core.keymem.key_mem[4][72] ),
    .A2(_14804_),
    .ZN(_14807_));
 OAI21_X1 _38656_ (.A(_14807_),
    .B1(_14796_),
    .B2(_13716_),
    .ZN(_02086_));
 NAND2_X1 _38657_ (.A1(\core.keymem.key_mem[4][73] ),
    .A2(_14804_),
    .ZN(_14808_));
 BUF_X4 _38658_ (.A(_14764_),
    .Z(_14809_));
 OAI21_X1 _38659_ (.A(_14808_),
    .B1(_14809_),
    .B2(_12688_),
    .ZN(_02087_));
 NAND2_X1 _38660_ (.A1(\core.keymem.key_mem[4][74] ),
    .A2(_14804_),
    .ZN(_14810_));
 OAI21_X1 _38661_ (.A(_14810_),
    .B1(_14809_),
    .B2(_13726_),
    .ZN(_02088_));
 NAND2_X1 _38662_ (.A1(\core.keymem.key_mem[4][75] ),
    .A2(_14804_),
    .ZN(_14811_));
 OAI21_X1 _38663_ (.A(_14811_),
    .B1(_14809_),
    .B2(_13733_),
    .ZN(_02089_));
 BUF_X4 _38664_ (.A(_14757_),
    .Z(_14812_));
 MUX2_X1 _38665_ (.A(\core.keymem.key_mem[4][76] ),
    .B(_13741_),
    .S(_14812_),
    .Z(_02090_));
 MUX2_X1 _38666_ (.A(\core.keymem.key_mem[4][77] ),
    .B(_13751_),
    .S(_14812_),
    .Z(_02091_));
 NAND2_X1 _38667_ (.A1(\core.keymem.key_mem[4][78] ),
    .A2(_14804_),
    .ZN(_14813_));
 OAI21_X1 _38668_ (.A(_14813_),
    .B1(_14809_),
    .B2(_12708_),
    .ZN(_02092_));
 MUX2_X1 _38669_ (.A(\core.keymem.key_mem[4][79] ),
    .B(_13758_),
    .S(_14812_),
    .Z(_02093_));
 NAND2_X1 _38670_ (.A1(\core.keymem.key_mem[4][7] ),
    .A2(_14804_),
    .ZN(_14814_));
 OAI21_X1 _38671_ (.A(_14814_),
    .B1(_14809_),
    .B2(_13767_),
    .ZN(_02094_));
 MUX2_X1 _38672_ (.A(\core.keymem.key_mem[4][80] ),
    .B(_13769_),
    .S(_14812_),
    .Z(_02095_));
 NAND2_X1 _38673_ (.A1(\core.keymem.key_mem[4][81] ),
    .A2(_14804_),
    .ZN(_14815_));
 OAI21_X1 _38674_ (.A(_14815_),
    .B1(_14809_),
    .B2(_13775_),
    .ZN(_02096_));
 NAND2_X1 _38675_ (.A1(\core.keymem.key_mem[4][82] ),
    .A2(_14804_),
    .ZN(_14816_));
 OAI21_X1 _38676_ (.A(_14816_),
    .B1(_14809_),
    .B2(_13783_),
    .ZN(_02097_));
 NAND2_X1 _38677_ (.A1(\core.keymem.key_mem[4][83] ),
    .A2(_14764_),
    .ZN(_14817_));
 OAI21_X1 _38678_ (.A(_14817_),
    .B1(_14809_),
    .B2(_13791_),
    .ZN(_02098_));
 NAND2_X1 _38679_ (.A1(\core.keymem.key_mem[4][84] ),
    .A2(_14764_),
    .ZN(_14818_));
 OAI21_X1 _38680_ (.A(_14818_),
    .B1(_14809_),
    .B2(_12725_),
    .ZN(_02099_));
 MUX2_X1 _38681_ (.A(\core.keymem.key_mem[4][85] ),
    .B(_13798_),
    .S(_14812_),
    .Z(_02100_));
 MUX2_X1 _38682_ (.A(\core.keymem.key_mem[4][86] ),
    .B(_12741_),
    .S(_14812_),
    .Z(_02101_));
 MUX2_X1 _38683_ (.A(\core.keymem.key_mem[4][87] ),
    .B(_13804_),
    .S(_14812_),
    .Z(_02102_));
 MUX2_X1 _38684_ (.A(\core.keymem.key_mem[4][88] ),
    .B(_13810_),
    .S(_14812_),
    .Z(_02103_));
 MUX2_X1 _38685_ (.A(\core.keymem.key_mem[4][89] ),
    .B(_13818_),
    .S(_14812_),
    .Z(_02104_));
 MUX2_X1 _38686_ (.A(\core.keymem.key_mem[4][8] ),
    .B(_13854_),
    .S(_14812_),
    .Z(_02105_));
 MUX2_X1 _38687_ (.A(\core.keymem.key_mem[4][90] ),
    .B(_13860_),
    .S(_14758_),
    .Z(_02106_));
 NAND2_X1 _38688_ (.A1(\core.keymem.key_mem[4][91] ),
    .A2(_14764_),
    .ZN(_14819_));
 OAI21_X1 _38689_ (.A(_14819_),
    .B1(_14809_),
    .B2(_13870_),
    .ZN(_02107_));
 NAND2_X1 _38690_ (.A1(\core.keymem.key_mem[4][92] ),
    .A2(_14764_),
    .ZN(_14820_));
 OAI21_X1 _38691_ (.A(_14820_),
    .B1(_14762_),
    .B2(_13880_),
    .ZN(_02108_));
 MUX2_X1 _38692_ (.A(\core.keymem.key_mem[4][93] ),
    .B(_13889_),
    .S(_14758_),
    .Z(_02109_));
 MUX2_X1 _38693_ (.A(\core.keymem.key_mem[4][94] ),
    .B(_13896_),
    .S(_14758_),
    .Z(_02110_));
 MUX2_X1 _38694_ (.A(\core.keymem.key_mem[4][95] ),
    .B(_13903_),
    .S(_14758_),
    .Z(_02111_));
 MUX2_X1 _38695_ (.A(\core.keymem.key_mem[4][96] ),
    .B(_13907_),
    .S(_14758_),
    .Z(_02112_));
 NAND2_X1 _38696_ (.A1(\core.keymem.key_mem[4][97] ),
    .A2(_14764_),
    .ZN(_14821_));
 OAI21_X1 _38697_ (.A(_14821_),
    .B1(_14762_),
    .B2(_12777_),
    .ZN(_02113_));
 NAND2_X1 _38698_ (.A1(\core.keymem.key_mem[4][98] ),
    .A2(_14764_),
    .ZN(_14822_));
 OAI21_X1 _38699_ (.A(_14822_),
    .B1(_14762_),
    .B2(_13910_),
    .ZN(_02114_));
 MUX2_X1 _38700_ (.A(\core.keymem.key_mem[4][99] ),
    .B(_12800_),
    .S(_14758_),
    .Z(_02115_));
 MUX2_X1 _38701_ (.A(\core.keymem.key_mem[4][9] ),
    .B(_13919_),
    .S(_14758_),
    .Z(_02116_));
 NOR2_X4 _38702_ (.A1(_14056_),
    .A2(_14756_),
    .ZN(_14823_));
 BUF_X4 _38703_ (.A(_14823_),
    .Z(_14824_));
 BUF_X4 _38704_ (.A(_14824_),
    .Z(_14825_));
 MUX2_X1 _38705_ (.A(\core.keymem.key_mem[5][0] ),
    .B(_11843_),
    .S(_14825_),
    .Z(_02117_));
 MUX2_X1 _38706_ (.A(\core.keymem.key_mem[5][100] ),
    .B(_11872_),
    .S(_14825_),
    .Z(_02118_));
 MUX2_X1 _38707_ (.A(\core.keymem.key_mem[5][101] ),
    .B(_12813_),
    .S(_14825_),
    .Z(_02119_));
 MUX2_X1 _38708_ (.A(\core.keymem.key_mem[5][102] ),
    .B(_11905_),
    .S(_14825_),
    .Z(_02120_));
 MUX2_X1 _38709_ (.A(\core.keymem.key_mem[5][103] ),
    .B(_11928_),
    .S(_14825_),
    .Z(_02121_));
 OR2_X1 _38710_ (.A1(_14056_),
    .A2(_14756_),
    .ZN(_14826_));
 CLKBUF_X3 _38711_ (.A(_14826_),
    .Z(_14827_));
 BUF_X4 _38712_ (.A(_14827_),
    .Z(_14828_));
 NAND2_X1 _38713_ (.A1(\core.keymem.key_mem[5][104] ),
    .A2(_14828_),
    .ZN(_14829_));
 BUF_X4 _38714_ (.A(_14827_),
    .Z(_14830_));
 BUF_X4 _38715_ (.A(_14830_),
    .Z(_14831_));
 OAI21_X1 _38716_ (.A(_14829_),
    .B1(_14831_),
    .B2(_12822_),
    .ZN(_02122_));
 MUX2_X1 _38717_ (.A(\core.keymem.key_mem[5][105] ),
    .B(_12830_),
    .S(_14825_),
    .Z(_02123_));
 BUF_X4 _38718_ (.A(_14824_),
    .Z(_14832_));
 MUX2_X1 _38719_ (.A(\core.keymem.key_mem[5][106] ),
    .B(_12832_),
    .S(_14832_),
    .Z(_02124_));
 MUX2_X1 _38720_ (.A(\core.keymem.key_mem[5][107] ),
    .B(_11966_),
    .S(_14832_),
    .Z(_02125_));
 MUX2_X1 _38721_ (.A(\core.keymem.key_mem[5][108] ),
    .B(_11980_),
    .S(_14832_),
    .Z(_02126_));
 MUX2_X1 _38722_ (.A(\core.keymem.key_mem[5][109] ),
    .B(_12842_),
    .S(_14832_),
    .Z(_02127_));
 NAND2_X1 _38723_ (.A1(\core.keymem.key_mem[5][10] ),
    .A2(_14828_),
    .ZN(_14833_));
 OAI21_X1 _38724_ (.A(_14833_),
    .B1(_14831_),
    .B2(_12858_),
    .ZN(_02128_));
 MUX2_X1 _38725_ (.A(\core.keymem.key_mem[5][110] ),
    .B(_12859_),
    .S(_14832_),
    .Z(_02129_));
 MUX2_X1 _38726_ (.A(\core.keymem.key_mem[5][111] ),
    .B(_12016_),
    .S(_14832_),
    .Z(_02130_));
 MUX2_X1 _38727_ (.A(\core.keymem.key_mem[5][112] ),
    .B(_12030_),
    .S(_14832_),
    .Z(_02131_));
 MUX2_X1 _38728_ (.A(\core.keymem.key_mem[5][113] ),
    .B(_12868_),
    .S(_14832_),
    .Z(_02132_));
 MUX2_X1 _38729_ (.A(\core.keymem.key_mem[5][114] ),
    .B(_12869_),
    .S(_14832_),
    .Z(_02133_));
 MUX2_X1 _38730_ (.A(\core.keymem.key_mem[5][115] ),
    .B(_12058_),
    .S(_14832_),
    .Z(_02134_));
 BUF_X4 _38731_ (.A(_14824_),
    .Z(_14834_));
 MUX2_X1 _38732_ (.A(\core.keymem.key_mem[5][116] ),
    .B(_12076_),
    .S(_14834_),
    .Z(_02135_));
 MUX2_X1 _38733_ (.A(\core.keymem.key_mem[5][117] ),
    .B(_12877_),
    .S(_14834_),
    .Z(_02136_));
 MUX2_X1 _38734_ (.A(\core.keymem.key_mem[5][118] ),
    .B(_12882_),
    .S(_14834_),
    .Z(_02137_));
 MUX2_X1 _38735_ (.A(\core.keymem.key_mem[5][119] ),
    .B(_12095_),
    .S(_14834_),
    .Z(_02138_));
 NAND2_X1 _38736_ (.A1(\core.keymem.key_mem[5][11] ),
    .A2(_14828_),
    .ZN(_14835_));
 OAI21_X1 _38737_ (.A(_14835_),
    .B1(_14831_),
    .B2(_12895_),
    .ZN(_02139_));
 MUX2_X1 _38738_ (.A(\core.keymem.key_mem[5][120] ),
    .B(_12123_),
    .S(_14834_),
    .Z(_02140_));
 MUX2_X1 _38739_ (.A(\core.keymem.key_mem[5][121] ),
    .B(_12159_),
    .S(_14834_),
    .Z(_02141_));
 MUX2_X1 _38740_ (.A(\core.keymem.key_mem[5][122] ),
    .B(_12903_),
    .S(_14834_),
    .Z(_02142_));
 NAND2_X1 _38741_ (.A1(\core.keymem.key_mem[5][123] ),
    .A2(_14828_),
    .ZN(_14836_));
 OAI21_X1 _38742_ (.A(_14836_),
    .B1(_14831_),
    .B2(_12181_),
    .ZN(_02143_));
 NAND2_X1 _38743_ (.A1(\core.keymem.key_mem[5][124] ),
    .A2(_14828_),
    .ZN(_14837_));
 OAI21_X1 _38744_ (.A(_14837_),
    .B1(_14831_),
    .B2(_12926_),
    .ZN(_02144_));
 MUX2_X1 _38745_ (.A(\core.keymem.key_mem[5][125] ),
    .B(_12932_),
    .S(_14834_),
    .Z(_02145_));
 NAND2_X1 _38746_ (.A1(\core.keymem.key_mem[5][126] ),
    .A2(_14828_),
    .ZN(_14838_));
 OAI21_X1 _38747_ (.A(_14838_),
    .B1(_14831_),
    .B2(_12206_),
    .ZN(_02146_));
 MUX2_X1 _38748_ (.A(\core.keymem.key_mem[5][127] ),
    .B(_12945_),
    .S(_14834_),
    .Z(_02147_));
 MUX2_X1 _38749_ (.A(\core.keymem.key_mem[5][12] ),
    .B(_12958_),
    .S(_14834_),
    .Z(_02148_));
 BUF_X4 _38750_ (.A(_14823_),
    .Z(_14839_));
 MUX2_X1 _38751_ (.A(\core.keymem.key_mem[5][13] ),
    .B(_12974_),
    .S(_14839_),
    .Z(_02149_));
 NOR2_X1 _38752_ (.A1(\core.keymem.key_mem[5][14] ),
    .A2(_14825_),
    .ZN(_14840_));
 AOI21_X1 _38753_ (.A(_14840_),
    .B1(_14825_),
    .B2(_13007_),
    .ZN(_02150_));
 MUX2_X1 _38754_ (.A(\core.keymem.key_mem[5][15] ),
    .B(_13017_),
    .S(_14839_),
    .Z(_02151_));
 MUX2_X1 _38755_ (.A(\core.keymem.key_mem[5][16] ),
    .B(_13029_),
    .S(_14839_),
    .Z(_02152_));
 NAND2_X1 _38756_ (.A1(\core.keymem.key_mem[5][17] ),
    .A2(_14828_),
    .ZN(_14841_));
 OAI21_X1 _38757_ (.A(_14841_),
    .B1(_14831_),
    .B2(_13042_),
    .ZN(_02153_));
 MUX2_X1 _38758_ (.A(\core.keymem.key_mem[5][18] ),
    .B(_13094_),
    .S(_14839_),
    .Z(_02154_));
 BUF_X4 _38759_ (.A(_14827_),
    .Z(_14842_));
 NAND2_X1 _38760_ (.A1(\core.keymem.key_mem[5][19] ),
    .A2(_14842_),
    .ZN(_14843_));
 OAI21_X1 _38761_ (.A(_14843_),
    .B1(_14831_),
    .B2(_13109_),
    .ZN(_02155_));
 MUX2_X1 _38762_ (.A(\core.keymem.key_mem[5][1] ),
    .B(_13134_),
    .S(_14839_),
    .Z(_02156_));
 MUX2_X1 _38763_ (.A(\core.keymem.key_mem[5][20] ),
    .B(_13146_),
    .S(_14839_),
    .Z(_02157_));
 MUX2_X1 _38764_ (.A(\core.keymem.key_mem[5][21] ),
    .B(_13155_),
    .S(_14839_),
    .Z(_02158_));
 NOR2_X1 _38765_ (.A1(\core.keymem.key_mem[5][22] ),
    .A2(_14825_),
    .ZN(_14844_));
 AOI21_X1 _38766_ (.A(_14844_),
    .B1(_14825_),
    .B2(_13191_),
    .ZN(_02159_));
 MUX2_X1 _38767_ (.A(\core.keymem.key_mem[5][23] ),
    .B(_13196_),
    .S(_14839_),
    .Z(_02160_));
 NAND2_X1 _38768_ (.A1(\core.keymem.key_mem[5][24] ),
    .A2(_14842_),
    .ZN(_14845_));
 OAI21_X1 _38769_ (.A(_14845_),
    .B1(_14831_),
    .B2(_13212_),
    .ZN(_02161_));
 MUX2_X1 _38770_ (.A(\core.keymem.key_mem[5][25] ),
    .B(_13233_),
    .S(_14839_),
    .Z(_02162_));
 MUX2_X1 _38771_ (.A(\core.keymem.key_mem[5][26] ),
    .B(_13241_),
    .S(_14839_),
    .Z(_02163_));
 BUF_X4 _38772_ (.A(_14823_),
    .Z(_14846_));
 MUX2_X1 _38773_ (.A(\core.keymem.key_mem[5][27] ),
    .B(_13284_),
    .S(_14846_),
    .Z(_02164_));
 MUX2_X1 _38774_ (.A(\core.keymem.key_mem[5][28] ),
    .B(_13325_),
    .S(_14846_),
    .Z(_02165_));
 MUX2_X1 _38775_ (.A(\core.keymem.key_mem[5][29] ),
    .B(_13329_),
    .S(_14846_),
    .Z(_02166_));
 NAND2_X1 _38776_ (.A1(\core.keymem.key_mem[5][2] ),
    .A2(_14842_),
    .ZN(_14847_));
 OAI21_X1 _38777_ (.A(_14847_),
    .B1(_14831_),
    .B2(_13335_),
    .ZN(_02167_));
 MUX2_X1 _38778_ (.A(\core.keymem.key_mem[5][30] ),
    .B(_13379_),
    .S(_14846_),
    .Z(_02168_));
 MUX2_X1 _38779_ (.A(\core.keymem.key_mem[5][31] ),
    .B(_13395_),
    .S(_14846_),
    .Z(_02169_));
 MUX2_X1 _38780_ (.A(\core.keymem.key_mem[5][32] ),
    .B(_13396_),
    .S(_14846_),
    .Z(_02170_));
 MUX2_X1 _38781_ (.A(\core.keymem.key_mem[5][33] ),
    .B(_13402_),
    .S(_14846_),
    .Z(_02171_));
 MUX2_X1 _38782_ (.A(\core.keymem.key_mem[5][34] ),
    .B(_13403_),
    .S(_14846_),
    .Z(_02172_));
 MUX2_X1 _38783_ (.A(\core.keymem.key_mem[5][35] ),
    .B(_13405_),
    .S(_14846_),
    .Z(_02173_));
 NAND2_X1 _38784_ (.A1(\core.keymem.key_mem[5][36] ),
    .A2(_14842_),
    .ZN(_14848_));
 BUF_X4 _38785_ (.A(_14830_),
    .Z(_14849_));
 OAI21_X1 _38786_ (.A(_14848_),
    .B1(_14849_),
    .B2(_13407_),
    .ZN(_02174_));
 NAND2_X1 _38787_ (.A1(\core.keymem.key_mem[5][37] ),
    .A2(_14842_),
    .ZN(_14850_));
 OAI21_X1 _38788_ (.A(_14850_),
    .B1(_14849_),
    .B2(_12438_),
    .ZN(_02175_));
 MUX2_X1 _38789_ (.A(\core.keymem.key_mem[5][38] ),
    .B(_13410_),
    .S(_14846_),
    .Z(_02176_));
 NAND2_X1 _38790_ (.A1(\core.keymem.key_mem[5][39] ),
    .A2(_14842_),
    .ZN(_14851_));
 OAI21_X1 _38791_ (.A(_14851_),
    .B1(_14849_),
    .B2(_13435_),
    .ZN(_02177_));
 NAND2_X1 _38792_ (.A1(\core.keymem.key_mem[5][3] ),
    .A2(_14842_),
    .ZN(_14852_));
 OAI21_X1 _38793_ (.A(_14852_),
    .B1(_14849_),
    .B2(_13448_),
    .ZN(_02178_));
 NAND2_X1 _38794_ (.A1(\core.keymem.key_mem[5][40] ),
    .A2(_14842_),
    .ZN(_14853_));
 OAI21_X1 _38795_ (.A(_14853_),
    .B1(_14849_),
    .B2(_13457_),
    .ZN(_02179_));
 BUF_X4 _38796_ (.A(_14823_),
    .Z(_14854_));
 MUX2_X1 _38797_ (.A(\core.keymem.key_mem[5][41] ),
    .B(_13467_),
    .S(_14854_),
    .Z(_02180_));
 MUX2_X1 _38798_ (.A(\core.keymem.key_mem[5][42] ),
    .B(_13490_),
    .S(_14854_),
    .Z(_02181_));
 NAND2_X1 _38799_ (.A1(\core.keymem.key_mem[5][43] ),
    .A2(_14842_),
    .ZN(_14855_));
 OAI21_X1 _38800_ (.A(_14855_),
    .B1(_14849_),
    .B2(_13496_),
    .ZN(_02182_));
 MUX2_X1 _38801_ (.A(\core.keymem.key_mem[5][44] ),
    .B(_13497_),
    .S(_14854_),
    .Z(_02183_));
 NAND2_X1 _38802_ (.A1(\core.keymem.key_mem[5][45] ),
    .A2(_14842_),
    .ZN(_14856_));
 OAI21_X1 _38803_ (.A(_14856_),
    .B1(_14849_),
    .B2(_13510_),
    .ZN(_02184_));
 BUF_X4 _38804_ (.A(_14827_),
    .Z(_14857_));
 NAND2_X1 _38805_ (.A1(\core.keymem.key_mem[5][46] ),
    .A2(_14857_),
    .ZN(_14858_));
 OAI21_X1 _38806_ (.A(_14858_),
    .B1(_14849_),
    .B2(_13517_),
    .ZN(_02185_));
 NAND2_X1 _38807_ (.A1(\core.keymem.key_mem[5][47] ),
    .A2(_14857_),
    .ZN(_14859_));
 OAI21_X1 _38808_ (.A(_14859_),
    .B1(_14849_),
    .B2(_12519_),
    .ZN(_02186_));
 NAND2_X1 _38809_ (.A1(\core.keymem.key_mem[5][48] ),
    .A2(_14857_),
    .ZN(_14860_));
 OAI21_X1 _38810_ (.A(_14860_),
    .B1(_14849_),
    .B2(_12531_),
    .ZN(_02187_));
 NAND2_X1 _38811_ (.A1(\core.keymem.key_mem[5][49] ),
    .A2(_14857_),
    .ZN(_14861_));
 BUF_X4 _38812_ (.A(_14830_),
    .Z(_14862_));
 OAI21_X1 _38813_ (.A(_14861_),
    .B1(_14862_),
    .B2(_13529_),
    .ZN(_02188_));
 MUX2_X1 _38814_ (.A(\core.keymem.key_mem[5][4] ),
    .B(_13538_),
    .S(_14854_),
    .Z(_02189_));
 MUX2_X1 _38815_ (.A(\core.keymem.key_mem[5][50] ),
    .B(_13557_),
    .S(_14854_),
    .Z(_02190_));
 MUX2_X1 _38816_ (.A(\core.keymem.key_mem[5][51] ),
    .B(_13564_),
    .S(_14854_),
    .Z(_02191_));
 NAND2_X1 _38817_ (.A1(\core.keymem.key_mem[5][52] ),
    .A2(_14857_),
    .ZN(_14863_));
 OAI21_X1 _38818_ (.A(_14863_),
    .B1(_14862_),
    .B2(_12567_),
    .ZN(_02192_));
 NAND2_X1 _38819_ (.A1(\core.keymem.key_mem[5][53] ),
    .A2(_14857_),
    .ZN(_14864_));
 OAI21_X1 _38820_ (.A(_14864_),
    .B1(_14862_),
    .B2(_12583_),
    .ZN(_02193_));
 NAND2_X1 _38821_ (.A1(\core.keymem.key_mem[5][54] ),
    .A2(_14857_),
    .ZN(_14865_));
 OAI21_X1 _38822_ (.A(_14865_),
    .B1(_14862_),
    .B2(_13575_),
    .ZN(_02194_));
 MUX2_X1 _38823_ (.A(\core.keymem.key_mem[5][55] ),
    .B(_13581_),
    .S(_14854_),
    .Z(_02195_));
 MUX2_X1 _38824_ (.A(\core.keymem.key_mem[5][56] ),
    .B(_13589_),
    .S(_14854_),
    .Z(_02196_));
 MUX2_X1 _38825_ (.A(\core.keymem.key_mem[5][57] ),
    .B(_13604_),
    .S(_14854_),
    .Z(_02197_));
 MUX2_X1 _38826_ (.A(\core.keymem.key_mem[5][58] ),
    .B(_13611_),
    .S(_14854_),
    .Z(_02198_));
 BUF_X4 _38827_ (.A(_14823_),
    .Z(_14866_));
 MUX2_X1 _38828_ (.A(\core.keymem.key_mem[5][59] ),
    .B(_13616_),
    .S(_14866_),
    .Z(_02199_));
 MUX2_X1 _38829_ (.A(\core.keymem.key_mem[5][5] ),
    .B(_12605_),
    .S(_14866_),
    .Z(_02200_));
 MUX2_X1 _38830_ (.A(\core.keymem.key_mem[5][60] ),
    .B(_13622_),
    .S(_14866_),
    .Z(_02201_));
 MUX2_X1 _38831_ (.A(\core.keymem.key_mem[5][61] ),
    .B(_13632_),
    .S(_14866_),
    .Z(_02202_));
 MUX2_X1 _38832_ (.A(\core.keymem.key_mem[5][62] ),
    .B(_13637_),
    .S(_14866_),
    .Z(_02203_));
 MUX2_X1 _38833_ (.A(\core.keymem.key_mem[5][63] ),
    .B(_13659_),
    .S(_14866_),
    .Z(_02204_));
 MUX2_X1 _38834_ (.A(\core.keymem.key_mem[5][64] ),
    .B(_12621_),
    .S(_14866_),
    .Z(_02205_));
 NAND2_X1 _38835_ (.A1(\core.keymem.key_mem[5][65] ),
    .A2(_14857_),
    .ZN(_14867_));
 OAI21_X1 _38836_ (.A(_14867_),
    .B1(_14862_),
    .B2(_13673_),
    .ZN(_02206_));
 MUX2_X1 _38837_ (.A(\core.keymem.key_mem[5][66] ),
    .B(_13681_),
    .S(_14866_),
    .Z(_02207_));
 NAND2_X1 _38838_ (.A1(\core.keymem.key_mem[5][67] ),
    .A2(_14857_),
    .ZN(_14868_));
 OAI21_X1 _38839_ (.A(_14868_),
    .B1(_14862_),
    .B2(_13690_),
    .ZN(_02208_));
 NAND2_X1 _38840_ (.A1(\core.keymem.key_mem[5][68] ),
    .A2(_14857_),
    .ZN(_14869_));
 OAI21_X1 _38841_ (.A(_14869_),
    .B1(_14862_),
    .B2(_12634_),
    .ZN(_02209_));
 BUF_X4 _38842_ (.A(_14827_),
    .Z(_14870_));
 NAND2_X1 _38843_ (.A1(\core.keymem.key_mem[5][69] ),
    .A2(_14870_),
    .ZN(_14871_));
 OAI21_X1 _38844_ (.A(_14871_),
    .B1(_14862_),
    .B2(_13700_),
    .ZN(_02210_));
 MUX2_X1 _38845_ (.A(\core.keymem.key_mem[5][6] ),
    .B(_13711_),
    .S(_14866_),
    .Z(_02211_));
 MUX2_X1 _38846_ (.A(\core.keymem.key_mem[5][70] ),
    .B(_13713_),
    .S(_14866_),
    .Z(_02212_));
 NAND2_X1 _38847_ (.A1(\core.keymem.key_mem[5][71] ),
    .A2(_14870_),
    .ZN(_14872_));
 OAI21_X1 _38848_ (.A(_14872_),
    .B1(_14862_),
    .B2(_12658_),
    .ZN(_02213_));
 NAND2_X1 _38849_ (.A1(\core.keymem.key_mem[5][72] ),
    .A2(_14870_),
    .ZN(_14873_));
 OAI21_X1 _38850_ (.A(_14873_),
    .B1(_14862_),
    .B2(_13716_),
    .ZN(_02214_));
 NAND2_X1 _38851_ (.A1(\core.keymem.key_mem[5][73] ),
    .A2(_14870_),
    .ZN(_14874_));
 BUF_X4 _38852_ (.A(_14830_),
    .Z(_14875_));
 OAI21_X1 _38853_ (.A(_14874_),
    .B1(_14875_),
    .B2(_12687_),
    .ZN(_02215_));
 NAND2_X1 _38854_ (.A1(\core.keymem.key_mem[5][74] ),
    .A2(_14870_),
    .ZN(_14876_));
 OAI21_X1 _38855_ (.A(_14876_),
    .B1(_14875_),
    .B2(_13726_),
    .ZN(_02216_));
 NAND2_X1 _38856_ (.A1(\core.keymem.key_mem[5][75] ),
    .A2(_14870_),
    .ZN(_14877_));
 OAI21_X1 _38857_ (.A(_14877_),
    .B1(_14875_),
    .B2(_13733_),
    .ZN(_02217_));
 BUF_X4 _38858_ (.A(_14823_),
    .Z(_14878_));
 MUX2_X1 _38859_ (.A(\core.keymem.key_mem[5][76] ),
    .B(_13741_),
    .S(_14878_),
    .Z(_02218_));
 MUX2_X1 _38860_ (.A(\core.keymem.key_mem[5][77] ),
    .B(_13751_),
    .S(_14878_),
    .Z(_02219_));
 NAND2_X1 _38861_ (.A1(\core.keymem.key_mem[5][78] ),
    .A2(_14870_),
    .ZN(_14879_));
 OAI21_X1 _38862_ (.A(_14879_),
    .B1(_14875_),
    .B2(_12707_),
    .ZN(_02220_));
 MUX2_X1 _38863_ (.A(\core.keymem.key_mem[5][79] ),
    .B(_13758_),
    .S(_14878_),
    .Z(_02221_));
 NAND2_X1 _38864_ (.A1(\core.keymem.key_mem[5][7] ),
    .A2(_14870_),
    .ZN(_14880_));
 OAI21_X1 _38865_ (.A(_14880_),
    .B1(_14875_),
    .B2(_13767_),
    .ZN(_02222_));
 MUX2_X1 _38866_ (.A(\core.keymem.key_mem[5][80] ),
    .B(_13769_),
    .S(_14878_),
    .Z(_02223_));
 NAND2_X1 _38867_ (.A1(\core.keymem.key_mem[5][81] ),
    .A2(_14870_),
    .ZN(_14881_));
 OAI21_X1 _38868_ (.A(_14881_),
    .B1(_14875_),
    .B2(_13775_),
    .ZN(_02224_));
 NAND2_X1 _38869_ (.A1(\core.keymem.key_mem[5][82] ),
    .A2(_14870_),
    .ZN(_14882_));
 OAI21_X1 _38870_ (.A(_14882_),
    .B1(_14875_),
    .B2(_13783_),
    .ZN(_02225_));
 NAND2_X1 _38871_ (.A1(\core.keymem.key_mem[5][83] ),
    .A2(_14830_),
    .ZN(_14883_));
 OAI21_X1 _38872_ (.A(_14883_),
    .B1(_14875_),
    .B2(_13791_),
    .ZN(_02226_));
 NAND2_X1 _38873_ (.A1(\core.keymem.key_mem[5][84] ),
    .A2(_14830_),
    .ZN(_14884_));
 OAI21_X1 _38874_ (.A(_14884_),
    .B1(_14875_),
    .B2(_12724_),
    .ZN(_02227_));
 MUX2_X1 _38875_ (.A(\core.keymem.key_mem[5][85] ),
    .B(_13798_),
    .S(_14878_),
    .Z(_02228_));
 MUX2_X1 _38876_ (.A(\core.keymem.key_mem[5][86] ),
    .B(_12740_),
    .S(_14878_),
    .Z(_02229_));
 MUX2_X1 _38877_ (.A(\core.keymem.key_mem[5][87] ),
    .B(_13804_),
    .S(_14878_),
    .Z(_02230_));
 MUX2_X1 _38878_ (.A(\core.keymem.key_mem[5][88] ),
    .B(_13810_),
    .S(_14878_),
    .Z(_02231_));
 MUX2_X1 _38879_ (.A(\core.keymem.key_mem[5][89] ),
    .B(_13818_),
    .S(_14878_),
    .Z(_02232_));
 MUX2_X1 _38880_ (.A(\core.keymem.key_mem[5][8] ),
    .B(_13854_),
    .S(_14878_),
    .Z(_02233_));
 MUX2_X1 _38881_ (.A(\core.keymem.key_mem[5][90] ),
    .B(_13860_),
    .S(_14824_),
    .Z(_02234_));
 NAND2_X1 _38882_ (.A1(\core.keymem.key_mem[5][91] ),
    .A2(_14830_),
    .ZN(_14885_));
 OAI21_X1 _38883_ (.A(_14885_),
    .B1(_14875_),
    .B2(_13870_),
    .ZN(_02235_));
 NAND2_X1 _38884_ (.A1(\core.keymem.key_mem[5][92] ),
    .A2(_14830_),
    .ZN(_14886_));
 OAI21_X1 _38885_ (.A(_14886_),
    .B1(_14828_),
    .B2(_13880_),
    .ZN(_02236_));
 MUX2_X1 _38886_ (.A(\core.keymem.key_mem[5][93] ),
    .B(_13889_),
    .S(_14824_),
    .Z(_02237_));
 MUX2_X1 _38887_ (.A(\core.keymem.key_mem[5][94] ),
    .B(_13896_),
    .S(_14824_),
    .Z(_02238_));
 MUX2_X1 _38888_ (.A(\core.keymem.key_mem[5][95] ),
    .B(_13903_),
    .S(_14824_),
    .Z(_02239_));
 MUX2_X1 _38889_ (.A(\core.keymem.key_mem[5][96] ),
    .B(_13907_),
    .S(_14824_),
    .Z(_02240_));
 NAND2_X1 _38890_ (.A1(\core.keymem.key_mem[5][97] ),
    .A2(_14830_),
    .ZN(_14887_));
 OAI21_X1 _38891_ (.A(_14887_),
    .B1(_14828_),
    .B2(_12776_),
    .ZN(_02241_));
 NAND2_X1 _38892_ (.A1(\core.keymem.key_mem[5][98] ),
    .A2(_14830_),
    .ZN(_14888_));
 OAI21_X1 _38893_ (.A(_14888_),
    .B1(_14828_),
    .B2(_13910_),
    .ZN(_02242_));
 MUX2_X1 _38894_ (.A(\core.keymem.key_mem[5][99] ),
    .B(_12799_),
    .S(_14824_),
    .Z(_02243_));
 MUX2_X1 _38895_ (.A(\core.keymem.key_mem[5][9] ),
    .B(_13919_),
    .S(_14824_),
    .Z(_02244_));
 NOR2_X4 _38896_ (.A1(_12804_),
    .A2(_14756_),
    .ZN(_14889_));
 BUF_X4 _38897_ (.A(_14889_),
    .Z(_14890_));
 BUF_X4 _38898_ (.A(_14890_),
    .Z(_14891_));
 MUX2_X1 _38899_ (.A(\core.keymem.key_mem[6][0] ),
    .B(_11843_),
    .S(_14891_),
    .Z(_02245_));
 MUX2_X1 _38900_ (.A(\core.keymem.key_mem[6][100] ),
    .B(_11872_),
    .S(_14891_),
    .Z(_02246_));
 MUX2_X1 _38901_ (.A(\core.keymem.key_mem[6][101] ),
    .B(_12813_),
    .S(_14891_),
    .Z(_02247_));
 MUX2_X1 _38902_ (.A(\core.keymem.key_mem[6][102] ),
    .B(_11905_),
    .S(_14891_),
    .Z(_02248_));
 MUX2_X1 _38903_ (.A(\core.keymem.key_mem[6][103] ),
    .B(_11928_),
    .S(_14891_),
    .Z(_02249_));
 OR2_X1 _38904_ (.A1(_12804_),
    .A2(_14756_),
    .ZN(_14892_));
 CLKBUF_X3 _38905_ (.A(_14892_),
    .Z(_14893_));
 BUF_X4 _38906_ (.A(_14893_),
    .Z(_14894_));
 NAND2_X1 _38907_ (.A1(\core.keymem.key_mem[6][104] ),
    .A2(_14894_),
    .ZN(_14895_));
 BUF_X4 _38908_ (.A(_14893_),
    .Z(_14896_));
 BUF_X4 _38909_ (.A(_14896_),
    .Z(_14897_));
 OAI21_X1 _38910_ (.A(_14895_),
    .B1(_14897_),
    .B2(_12822_),
    .ZN(_02250_));
 MUX2_X1 _38911_ (.A(\core.keymem.key_mem[6][105] ),
    .B(_12830_),
    .S(_14891_),
    .Z(_02251_));
 BUF_X4 _38912_ (.A(_14890_),
    .Z(_14898_));
 MUX2_X1 _38913_ (.A(\core.keymem.key_mem[6][106] ),
    .B(_12832_),
    .S(_14898_),
    .Z(_02252_));
 MUX2_X1 _38914_ (.A(\core.keymem.key_mem[6][107] ),
    .B(_11966_),
    .S(_14898_),
    .Z(_02253_));
 MUX2_X1 _38915_ (.A(\core.keymem.key_mem[6][108] ),
    .B(_11980_),
    .S(_14898_),
    .Z(_02254_));
 MUX2_X1 _38916_ (.A(\core.keymem.key_mem[6][109] ),
    .B(_12842_),
    .S(_14898_),
    .Z(_02255_));
 NAND2_X1 _38917_ (.A1(\core.keymem.key_mem[6][10] ),
    .A2(_14894_),
    .ZN(_14899_));
 OAI21_X1 _38918_ (.A(_14899_),
    .B1(_14897_),
    .B2(_12858_),
    .ZN(_02256_));
 MUX2_X1 _38919_ (.A(\core.keymem.key_mem[6][110] ),
    .B(_12859_),
    .S(_14898_),
    .Z(_02257_));
 MUX2_X1 _38920_ (.A(\core.keymem.key_mem[6][111] ),
    .B(_12016_),
    .S(_14898_),
    .Z(_02258_));
 MUX2_X1 _38921_ (.A(\core.keymem.key_mem[6][112] ),
    .B(_12030_),
    .S(_14898_),
    .Z(_02259_));
 MUX2_X1 _38922_ (.A(\core.keymem.key_mem[6][113] ),
    .B(_12868_),
    .S(_14898_),
    .Z(_02260_));
 MUX2_X1 _38923_ (.A(\core.keymem.key_mem[6][114] ),
    .B(_12869_),
    .S(_14898_),
    .Z(_02261_));
 MUX2_X1 _38924_ (.A(\core.keymem.key_mem[6][115] ),
    .B(_12058_),
    .S(_14898_),
    .Z(_02262_));
 BUF_X4 _38925_ (.A(_14890_),
    .Z(_14900_));
 MUX2_X1 _38926_ (.A(\core.keymem.key_mem[6][116] ),
    .B(_12076_),
    .S(_14900_),
    .Z(_02263_));
 MUX2_X1 _38927_ (.A(\core.keymem.key_mem[6][117] ),
    .B(_12877_),
    .S(_14900_),
    .Z(_02264_));
 MUX2_X1 _38928_ (.A(\core.keymem.key_mem[6][118] ),
    .B(_12882_),
    .S(_14900_),
    .Z(_02265_));
 MUX2_X1 _38929_ (.A(\core.keymem.key_mem[6][119] ),
    .B(_12095_),
    .S(_14900_),
    .Z(_02266_));
 NAND2_X1 _38930_ (.A1(\core.keymem.key_mem[6][11] ),
    .A2(_14894_),
    .ZN(_14901_));
 OAI21_X1 _38931_ (.A(_14901_),
    .B1(_14897_),
    .B2(_12895_),
    .ZN(_02267_));
 MUX2_X1 _38932_ (.A(\core.keymem.key_mem[6][120] ),
    .B(_12123_),
    .S(_14900_),
    .Z(_02268_));
 MUX2_X1 _38933_ (.A(\core.keymem.key_mem[6][121] ),
    .B(_12159_),
    .S(_14900_),
    .Z(_02269_));
 MUX2_X1 _38934_ (.A(\core.keymem.key_mem[6][122] ),
    .B(_12902_),
    .S(_14900_),
    .Z(_02270_));
 NAND2_X1 _38935_ (.A1(\core.keymem.key_mem[6][123] ),
    .A2(_14894_),
    .ZN(_14902_));
 OAI21_X1 _38936_ (.A(_14902_),
    .B1(_14897_),
    .B2(_12181_),
    .ZN(_02271_));
 NAND2_X1 _38937_ (.A1(\core.keymem.key_mem[6][124] ),
    .A2(_14894_),
    .ZN(_14903_));
 OAI21_X1 _38938_ (.A(_14903_),
    .B1(_14897_),
    .B2(_12926_),
    .ZN(_02272_));
 MUX2_X1 _38939_ (.A(\core.keymem.key_mem[6][125] ),
    .B(_12932_),
    .S(_14900_),
    .Z(_02273_));
 NAND2_X1 _38940_ (.A1(\core.keymem.key_mem[6][126] ),
    .A2(_14894_),
    .ZN(_14904_));
 OAI21_X1 _38941_ (.A(_14904_),
    .B1(_14897_),
    .B2(_12206_),
    .ZN(_02274_));
 MUX2_X1 _38942_ (.A(\core.keymem.key_mem[6][127] ),
    .B(_12944_),
    .S(_14900_),
    .Z(_02275_));
 MUX2_X1 _38943_ (.A(\core.keymem.key_mem[6][12] ),
    .B(_12958_),
    .S(_14900_),
    .Z(_02276_));
 BUF_X4 _38944_ (.A(_14889_),
    .Z(_14905_));
 MUX2_X1 _38945_ (.A(\core.keymem.key_mem[6][13] ),
    .B(_12974_),
    .S(_14905_),
    .Z(_02277_));
 NOR2_X1 _38946_ (.A1(\core.keymem.key_mem[6][14] ),
    .A2(_14891_),
    .ZN(_14906_));
 AOI21_X1 _38947_ (.A(_14906_),
    .B1(_14891_),
    .B2(_13007_),
    .ZN(_02278_));
 MUX2_X1 _38948_ (.A(\core.keymem.key_mem[6][15] ),
    .B(_13017_),
    .S(_14905_),
    .Z(_02279_));
 MUX2_X1 _38949_ (.A(\core.keymem.key_mem[6][16] ),
    .B(_13029_),
    .S(_14905_),
    .Z(_02280_));
 NAND2_X1 _38950_ (.A1(\core.keymem.key_mem[6][17] ),
    .A2(_14894_),
    .ZN(_14907_));
 OAI21_X1 _38951_ (.A(_14907_),
    .B1(_14897_),
    .B2(_13042_),
    .ZN(_02281_));
 MUX2_X1 _38952_ (.A(\core.keymem.key_mem[6][18] ),
    .B(_13094_),
    .S(_14905_),
    .Z(_02282_));
 BUF_X4 _38953_ (.A(_14893_),
    .Z(_14908_));
 NAND2_X1 _38954_ (.A1(\core.keymem.key_mem[6][19] ),
    .A2(_14908_),
    .ZN(_14909_));
 OAI21_X1 _38955_ (.A(_14909_),
    .B1(_14897_),
    .B2(_13109_),
    .ZN(_02283_));
 MUX2_X1 _38956_ (.A(\core.keymem.key_mem[6][1] ),
    .B(_13134_),
    .S(_14905_),
    .Z(_02284_));
 MUX2_X1 _38957_ (.A(\core.keymem.key_mem[6][20] ),
    .B(_13146_),
    .S(_14905_),
    .Z(_02285_));
 MUX2_X1 _38958_ (.A(\core.keymem.key_mem[6][21] ),
    .B(_13155_),
    .S(_14905_),
    .Z(_02286_));
 NOR2_X1 _38959_ (.A1(\core.keymem.key_mem[6][22] ),
    .A2(_14891_),
    .ZN(_14910_));
 AOI21_X1 _38960_ (.A(_14910_),
    .B1(_14891_),
    .B2(_13191_),
    .ZN(_02287_));
 MUX2_X1 _38961_ (.A(\core.keymem.key_mem[6][23] ),
    .B(_13196_),
    .S(_14905_),
    .Z(_02288_));
 NAND2_X1 _38962_ (.A1(\core.keymem.key_mem[6][24] ),
    .A2(_14908_),
    .ZN(_14911_));
 OAI21_X1 _38963_ (.A(_14911_),
    .B1(_14897_),
    .B2(_13212_),
    .ZN(_02289_));
 MUX2_X1 _38964_ (.A(\core.keymem.key_mem[6][25] ),
    .B(_13233_),
    .S(_14905_),
    .Z(_02290_));
 MUX2_X1 _38965_ (.A(\core.keymem.key_mem[6][26] ),
    .B(_13240_),
    .S(_14905_),
    .Z(_02291_));
 BUF_X4 _38966_ (.A(_14889_),
    .Z(_14912_));
 MUX2_X1 _38967_ (.A(\core.keymem.key_mem[6][27] ),
    .B(_13284_),
    .S(_14912_),
    .Z(_02292_));
 MUX2_X1 _38968_ (.A(\core.keymem.key_mem[6][28] ),
    .B(_13325_),
    .S(_14912_),
    .Z(_02293_));
 MUX2_X1 _38969_ (.A(\core.keymem.key_mem[6][29] ),
    .B(_13329_),
    .S(_14912_),
    .Z(_02294_));
 NAND2_X1 _38970_ (.A1(\core.keymem.key_mem[6][2] ),
    .A2(_14908_),
    .ZN(_14913_));
 OAI21_X1 _38971_ (.A(_14913_),
    .B1(_14897_),
    .B2(_13335_),
    .ZN(_02295_));
 MUX2_X1 _38972_ (.A(\core.keymem.key_mem[6][30] ),
    .B(_13379_),
    .S(_14912_),
    .Z(_02296_));
 MUX2_X1 _38973_ (.A(\core.keymem.key_mem[6][31] ),
    .B(_13395_),
    .S(_14912_),
    .Z(_02297_));
 MUX2_X1 _38974_ (.A(\core.keymem.key_mem[6][32] ),
    .B(_13396_),
    .S(_14912_),
    .Z(_02298_));
 MUX2_X1 _38975_ (.A(\core.keymem.key_mem[6][33] ),
    .B(_13401_),
    .S(_14912_),
    .Z(_02299_));
 MUX2_X1 _38976_ (.A(\core.keymem.key_mem[6][34] ),
    .B(_13403_),
    .S(_14912_),
    .Z(_02300_));
 MUX2_X1 _38977_ (.A(\core.keymem.key_mem[6][35] ),
    .B(_13405_),
    .S(_14912_),
    .Z(_02301_));
 NAND2_X1 _38978_ (.A1(\core.keymem.key_mem[6][36] ),
    .A2(_14908_),
    .ZN(_14914_));
 BUF_X4 _38979_ (.A(_14896_),
    .Z(_14915_));
 OAI21_X1 _38980_ (.A(_14914_),
    .B1(_14915_),
    .B2(_13407_),
    .ZN(_02302_));
 NAND2_X1 _38981_ (.A1(\core.keymem.key_mem[6][37] ),
    .A2(_14908_),
    .ZN(_14916_));
 OAI21_X1 _38982_ (.A(_14916_),
    .B1(_14915_),
    .B2(_12438_),
    .ZN(_02303_));
 MUX2_X1 _38983_ (.A(\core.keymem.key_mem[6][38] ),
    .B(_13410_),
    .S(_14912_),
    .Z(_02304_));
 NAND2_X1 _38984_ (.A1(\core.keymem.key_mem[6][39] ),
    .A2(_14908_),
    .ZN(_14917_));
 OAI21_X1 _38985_ (.A(_14917_),
    .B1(_14915_),
    .B2(_13435_),
    .ZN(_02305_));
 NAND2_X1 _38986_ (.A1(\core.keymem.key_mem[6][3] ),
    .A2(_14908_),
    .ZN(_14918_));
 OAI21_X1 _38987_ (.A(_14918_),
    .B1(_14915_),
    .B2(_13448_),
    .ZN(_02306_));
 NAND2_X1 _38988_ (.A1(\core.keymem.key_mem[6][40] ),
    .A2(_14908_),
    .ZN(_14919_));
 OAI21_X1 _38989_ (.A(_14919_),
    .B1(_14915_),
    .B2(_13456_),
    .ZN(_02307_));
 BUF_X4 _38990_ (.A(_14889_),
    .Z(_14920_));
 MUX2_X1 _38991_ (.A(\core.keymem.key_mem[6][41] ),
    .B(_13466_),
    .S(_14920_),
    .Z(_02308_));
 MUX2_X1 _38992_ (.A(\core.keymem.key_mem[6][42] ),
    .B(_13490_),
    .S(_14920_),
    .Z(_02309_));
 NAND2_X1 _38993_ (.A1(\core.keymem.key_mem[6][43] ),
    .A2(_14908_),
    .ZN(_14921_));
 OAI21_X1 _38994_ (.A(_14921_),
    .B1(_14915_),
    .B2(_13496_),
    .ZN(_02310_));
 MUX2_X1 _38995_ (.A(\core.keymem.key_mem[6][44] ),
    .B(_13497_),
    .S(_14920_),
    .Z(_02311_));
 NAND2_X1 _38996_ (.A1(\core.keymem.key_mem[6][45] ),
    .A2(_14908_),
    .ZN(_14922_));
 OAI21_X1 _38997_ (.A(_14922_),
    .B1(_14915_),
    .B2(_13510_),
    .ZN(_02312_));
 BUF_X4 _38998_ (.A(_14893_),
    .Z(_14923_));
 NAND2_X1 _38999_ (.A1(\core.keymem.key_mem[6][46] ),
    .A2(_14923_),
    .ZN(_14924_));
 OAI21_X1 _39000_ (.A(_14924_),
    .B1(_14915_),
    .B2(_13517_),
    .ZN(_02313_));
 NAND2_X1 _39001_ (.A1(\core.keymem.key_mem[6][47] ),
    .A2(_14923_),
    .ZN(_14925_));
 OAI21_X1 _39002_ (.A(_14925_),
    .B1(_14915_),
    .B2(_12519_),
    .ZN(_02314_));
 NAND2_X1 _39003_ (.A1(\core.keymem.key_mem[6][48] ),
    .A2(_14923_),
    .ZN(_14926_));
 OAI21_X1 _39004_ (.A(_14926_),
    .B1(_14915_),
    .B2(_12531_),
    .ZN(_02315_));
 NAND2_X1 _39005_ (.A1(\core.keymem.key_mem[6][49] ),
    .A2(_14923_),
    .ZN(_14927_));
 BUF_X4 _39006_ (.A(_14896_),
    .Z(_14928_));
 OAI21_X1 _39007_ (.A(_14927_),
    .B1(_14928_),
    .B2(_13528_),
    .ZN(_02316_));
 MUX2_X1 _39008_ (.A(\core.keymem.key_mem[6][4] ),
    .B(_13538_),
    .S(_14920_),
    .Z(_02317_));
 MUX2_X1 _39009_ (.A(\core.keymem.key_mem[6][50] ),
    .B(_13557_),
    .S(_14920_),
    .Z(_02318_));
 MUX2_X1 _39010_ (.A(\core.keymem.key_mem[6][51] ),
    .B(_13564_),
    .S(_14920_),
    .Z(_02319_));
 NAND2_X1 _39011_ (.A1(\core.keymem.key_mem[6][52] ),
    .A2(_14923_),
    .ZN(_14929_));
 OAI21_X1 _39012_ (.A(_14929_),
    .B1(_14928_),
    .B2(_12567_),
    .ZN(_02320_));
 NAND2_X1 _39013_ (.A1(\core.keymem.key_mem[6][53] ),
    .A2(_14923_),
    .ZN(_14930_));
 OAI21_X1 _39014_ (.A(_14930_),
    .B1(_14928_),
    .B2(_12583_),
    .ZN(_02321_));
 NAND2_X1 _39015_ (.A1(\core.keymem.key_mem[6][54] ),
    .A2(_14923_),
    .ZN(_14931_));
 OAI21_X1 _39016_ (.A(_14931_),
    .B1(_14928_),
    .B2(_13575_),
    .ZN(_02322_));
 MUX2_X1 _39017_ (.A(\core.keymem.key_mem[6][55] ),
    .B(_13581_),
    .S(_14920_),
    .Z(_02323_));
 MUX2_X1 _39018_ (.A(\core.keymem.key_mem[6][56] ),
    .B(_13589_),
    .S(_14920_),
    .Z(_02324_));
 MUX2_X1 _39019_ (.A(\core.keymem.key_mem[6][57] ),
    .B(_13604_),
    .S(_14920_),
    .Z(_02325_));
 MUX2_X1 _39020_ (.A(\core.keymem.key_mem[6][58] ),
    .B(_13611_),
    .S(_14920_),
    .Z(_02326_));
 BUF_X4 _39021_ (.A(_14889_),
    .Z(_14932_));
 MUX2_X1 _39022_ (.A(\core.keymem.key_mem[6][59] ),
    .B(_13616_),
    .S(_14932_),
    .Z(_02327_));
 MUX2_X1 _39023_ (.A(\core.keymem.key_mem[6][5] ),
    .B(_12605_),
    .S(_14932_),
    .Z(_02328_));
 MUX2_X1 _39024_ (.A(\core.keymem.key_mem[6][60] ),
    .B(_13622_),
    .S(_14932_),
    .Z(_02329_));
 MUX2_X1 _39025_ (.A(\core.keymem.key_mem[6][61] ),
    .B(_13632_),
    .S(_14932_),
    .Z(_02330_));
 MUX2_X1 _39026_ (.A(\core.keymem.key_mem[6][62] ),
    .B(_13637_),
    .S(_14932_),
    .Z(_02331_));
 MUX2_X1 _39027_ (.A(\core.keymem.key_mem[6][63] ),
    .B(_13659_),
    .S(_14932_),
    .Z(_02332_));
 MUX2_X1 _39028_ (.A(\core.keymem.key_mem[6][64] ),
    .B(_12621_),
    .S(_14932_),
    .Z(_02333_));
 NAND2_X1 _39029_ (.A1(\core.keymem.key_mem[6][65] ),
    .A2(_14923_),
    .ZN(_14933_));
 OAI21_X1 _39030_ (.A(_14933_),
    .B1(_14928_),
    .B2(_13672_),
    .ZN(_02334_));
 MUX2_X1 _39031_ (.A(\core.keymem.key_mem[6][66] ),
    .B(_13681_),
    .S(_14932_),
    .Z(_02335_));
 NAND2_X1 _39032_ (.A1(\core.keymem.key_mem[6][67] ),
    .A2(_14923_),
    .ZN(_14934_));
 OAI21_X1 _39033_ (.A(_14934_),
    .B1(_14928_),
    .B2(_13690_),
    .ZN(_02336_));
 NAND2_X1 _39034_ (.A1(\core.keymem.key_mem[6][68] ),
    .A2(_14923_),
    .ZN(_14935_));
 OAI21_X1 _39035_ (.A(_14935_),
    .B1(_14928_),
    .B2(_12634_),
    .ZN(_02337_));
 BUF_X4 _39036_ (.A(_14893_),
    .Z(_14936_));
 NAND2_X1 _39037_ (.A1(\core.keymem.key_mem[6][69] ),
    .A2(_14936_),
    .ZN(_14937_));
 OAI21_X1 _39038_ (.A(_14937_),
    .B1(_14928_),
    .B2(_13699_),
    .ZN(_02338_));
 MUX2_X1 _39039_ (.A(\core.keymem.key_mem[6][6] ),
    .B(_13710_),
    .S(_14932_),
    .Z(_02339_));
 MUX2_X1 _39040_ (.A(\core.keymem.key_mem[6][70] ),
    .B(_13713_),
    .S(_14932_),
    .Z(_02340_));
 NAND2_X1 _39041_ (.A1(\core.keymem.key_mem[6][71] ),
    .A2(_14936_),
    .ZN(_14938_));
 OAI21_X1 _39042_ (.A(_14938_),
    .B1(_14928_),
    .B2(_12658_),
    .ZN(_02341_));
 NAND2_X1 _39043_ (.A1(\core.keymem.key_mem[6][72] ),
    .A2(_14936_),
    .ZN(_14939_));
 OAI21_X1 _39044_ (.A(_14939_),
    .B1(_14928_),
    .B2(_13716_),
    .ZN(_02342_));
 NAND2_X1 _39045_ (.A1(\core.keymem.key_mem[6][73] ),
    .A2(_14936_),
    .ZN(_14940_));
 BUF_X4 _39046_ (.A(_14896_),
    .Z(_14941_));
 OAI21_X1 _39047_ (.A(_14940_),
    .B1(_14941_),
    .B2(_12687_),
    .ZN(_02343_));
 NAND2_X1 _39048_ (.A1(\core.keymem.key_mem[6][74] ),
    .A2(_14936_),
    .ZN(_14942_));
 OAI21_X1 _39049_ (.A(_14942_),
    .B1(_14941_),
    .B2(_13726_),
    .ZN(_02344_));
 NAND2_X1 _39050_ (.A1(\core.keymem.key_mem[6][75] ),
    .A2(_14936_),
    .ZN(_14943_));
 OAI21_X1 _39051_ (.A(_14943_),
    .B1(_14941_),
    .B2(_13732_),
    .ZN(_02345_));
 BUF_X4 _39052_ (.A(_14889_),
    .Z(_14944_));
 MUX2_X1 _39053_ (.A(\core.keymem.key_mem[6][76] ),
    .B(_13740_),
    .S(_14944_),
    .Z(_02346_));
 MUX2_X1 _39054_ (.A(\core.keymem.key_mem[6][77] ),
    .B(_13751_),
    .S(_14944_),
    .Z(_02347_));
 NAND2_X1 _39055_ (.A1(\core.keymem.key_mem[6][78] ),
    .A2(_14936_),
    .ZN(_14945_));
 OAI21_X1 _39056_ (.A(_14945_),
    .B1(_14941_),
    .B2(_12707_),
    .ZN(_02348_));
 MUX2_X1 _39057_ (.A(\core.keymem.key_mem[6][79] ),
    .B(_13758_),
    .S(_14944_),
    .Z(_02349_));
 NAND2_X1 _39058_ (.A1(\core.keymem.key_mem[6][7] ),
    .A2(_14936_),
    .ZN(_14946_));
 OAI21_X1 _39059_ (.A(_14946_),
    .B1(_14941_),
    .B2(_13766_),
    .ZN(_02350_));
 MUX2_X1 _39060_ (.A(\core.keymem.key_mem[6][80] ),
    .B(_13769_),
    .S(_14944_),
    .Z(_02351_));
 NAND2_X1 _39061_ (.A1(\core.keymem.key_mem[6][81] ),
    .A2(_14936_),
    .ZN(_14947_));
 OAI21_X1 _39062_ (.A(_14947_),
    .B1(_14941_),
    .B2(_13774_),
    .ZN(_02352_));
 NAND2_X1 _39063_ (.A1(\core.keymem.key_mem[6][82] ),
    .A2(_14936_),
    .ZN(_14948_));
 OAI21_X1 _39064_ (.A(_14948_),
    .B1(_14941_),
    .B2(_13782_),
    .ZN(_02353_));
 NAND2_X1 _39065_ (.A1(\core.keymem.key_mem[6][83] ),
    .A2(_14896_),
    .ZN(_14949_));
 OAI21_X1 _39066_ (.A(_14949_),
    .B1(_14941_),
    .B2(_13790_),
    .ZN(_02354_));
 NAND2_X1 _39067_ (.A1(\core.keymem.key_mem[6][84] ),
    .A2(_14896_),
    .ZN(_14950_));
 OAI21_X1 _39068_ (.A(_14950_),
    .B1(_14941_),
    .B2(_12724_),
    .ZN(_02355_));
 MUX2_X1 _39069_ (.A(\core.keymem.key_mem[6][85] ),
    .B(_13798_),
    .S(_14944_),
    .Z(_02356_));
 MUX2_X1 _39070_ (.A(\core.keymem.key_mem[6][86] ),
    .B(_12740_),
    .S(_14944_),
    .Z(_02357_));
 MUX2_X1 _39071_ (.A(\core.keymem.key_mem[6][87] ),
    .B(_13804_),
    .S(_14944_),
    .Z(_02358_));
 MUX2_X1 _39072_ (.A(\core.keymem.key_mem[6][88] ),
    .B(_13810_),
    .S(_14944_),
    .Z(_02359_));
 MUX2_X1 _39073_ (.A(\core.keymem.key_mem[6][89] ),
    .B(_13818_),
    .S(_14944_),
    .Z(_02360_));
 MUX2_X1 _39074_ (.A(\core.keymem.key_mem[6][8] ),
    .B(_13854_),
    .S(_14944_),
    .Z(_02361_));
 MUX2_X1 _39075_ (.A(\core.keymem.key_mem[6][90] ),
    .B(_13860_),
    .S(_14890_),
    .Z(_02362_));
 NAND2_X1 _39076_ (.A1(\core.keymem.key_mem[6][91] ),
    .A2(_14896_),
    .ZN(_14951_));
 OAI21_X1 _39077_ (.A(_14951_),
    .B1(_14941_),
    .B2(_13870_),
    .ZN(_02363_));
 NAND2_X1 _39078_ (.A1(\core.keymem.key_mem[6][92] ),
    .A2(_14896_),
    .ZN(_14952_));
 OAI21_X1 _39079_ (.A(_14952_),
    .B1(_14894_),
    .B2(_13880_),
    .ZN(_02364_));
 MUX2_X1 _39080_ (.A(\core.keymem.key_mem[6][93] ),
    .B(_13889_),
    .S(_14890_),
    .Z(_02365_));
 MUX2_X1 _39081_ (.A(\core.keymem.key_mem[6][94] ),
    .B(_13896_),
    .S(_14890_),
    .Z(_02366_));
 MUX2_X1 _39082_ (.A(\core.keymem.key_mem[6][95] ),
    .B(_13903_),
    .S(_14890_),
    .Z(_02367_));
 MUX2_X1 _39083_ (.A(\core.keymem.key_mem[6][96] ),
    .B(_13907_),
    .S(_14890_),
    .Z(_02368_));
 NAND2_X1 _39084_ (.A1(\core.keymem.key_mem[6][97] ),
    .A2(_14896_),
    .ZN(_14953_));
 OAI21_X1 _39085_ (.A(_14953_),
    .B1(_14894_),
    .B2(_12776_),
    .ZN(_02369_));
 NAND2_X1 _39086_ (.A1(\core.keymem.key_mem[6][98] ),
    .A2(_14896_),
    .ZN(_14954_));
 OAI21_X1 _39087_ (.A(_14954_),
    .B1(_14894_),
    .B2(_13910_),
    .ZN(_02370_));
 MUX2_X1 _39088_ (.A(\core.keymem.key_mem[6][99] ),
    .B(_12799_),
    .S(_14890_),
    .Z(_02371_));
 MUX2_X1 _39089_ (.A(\core.keymem.key_mem[6][9] ),
    .B(_13919_),
    .S(_14890_),
    .Z(_02372_));
 NOR2_X4 _39090_ (.A1(_13921_),
    .A2(_14756_),
    .ZN(_14955_));
 BUF_X4 _39091_ (.A(_14955_),
    .Z(_14956_));
 BUF_X4 _39092_ (.A(_14956_),
    .Z(_14957_));
 MUX2_X1 _39093_ (.A(\core.keymem.key_mem[7][0] ),
    .B(_11843_),
    .S(_14957_),
    .Z(_02373_));
 MUX2_X1 _39094_ (.A(\core.keymem.key_mem[7][100] ),
    .B(_11872_),
    .S(_14957_),
    .Z(_02374_));
 MUX2_X1 _39095_ (.A(\core.keymem.key_mem[7][101] ),
    .B(_12813_),
    .S(_14957_),
    .Z(_02375_));
 MUX2_X1 _39096_ (.A(\core.keymem.key_mem[7][102] ),
    .B(_11905_),
    .S(_14957_),
    .Z(_02376_));
 MUX2_X1 _39097_ (.A(\core.keymem.key_mem[7][103] ),
    .B(_11928_),
    .S(_14957_),
    .Z(_02377_));
 OR2_X1 _39098_ (.A1(_13921_),
    .A2(_14756_),
    .ZN(_14958_));
 CLKBUF_X3 _39099_ (.A(_14958_),
    .Z(_14959_));
 BUF_X4 _39100_ (.A(_14959_),
    .Z(_14960_));
 NAND2_X1 _39101_ (.A1(\core.keymem.key_mem[7][104] ),
    .A2(_14960_),
    .ZN(_14961_));
 BUF_X4 _39102_ (.A(_14959_),
    .Z(_14962_));
 BUF_X4 _39103_ (.A(_14962_),
    .Z(_14963_));
 OAI21_X1 _39104_ (.A(_14961_),
    .B1(_14963_),
    .B2(_12822_),
    .ZN(_02378_));
 MUX2_X1 _39105_ (.A(\core.keymem.key_mem[7][105] ),
    .B(_12830_),
    .S(_14957_),
    .Z(_02379_));
 BUF_X4 _39106_ (.A(_14956_),
    .Z(_14964_));
 MUX2_X1 _39107_ (.A(\core.keymem.key_mem[7][106] ),
    .B(_12831_),
    .S(_14964_),
    .Z(_02380_));
 MUX2_X1 _39108_ (.A(\core.keymem.key_mem[7][107] ),
    .B(_11966_),
    .S(_14964_),
    .Z(_02381_));
 MUX2_X1 _39109_ (.A(\core.keymem.key_mem[7][108] ),
    .B(_11980_),
    .S(_14964_),
    .Z(_02382_));
 MUX2_X1 _39110_ (.A(\core.keymem.key_mem[7][109] ),
    .B(_12842_),
    .S(_14964_),
    .Z(_02383_));
 NAND2_X1 _39111_ (.A1(\core.keymem.key_mem[7][10] ),
    .A2(_14960_),
    .ZN(_14965_));
 OAI21_X1 _39112_ (.A(_14965_),
    .B1(_14963_),
    .B2(_12858_),
    .ZN(_02384_));
 MUX2_X1 _39113_ (.A(\core.keymem.key_mem[7][110] ),
    .B(_12003_),
    .S(_14964_),
    .Z(_02385_));
 MUX2_X1 _39114_ (.A(\core.keymem.key_mem[7][111] ),
    .B(_12016_),
    .S(_14964_),
    .Z(_02386_));
 MUX2_X1 _39115_ (.A(\core.keymem.key_mem[7][112] ),
    .B(_12030_),
    .S(_14964_),
    .Z(_02387_));
 MUX2_X1 _39116_ (.A(\core.keymem.key_mem[7][113] ),
    .B(_12868_),
    .S(_14964_),
    .Z(_02388_));
 MUX2_X1 _39117_ (.A(\core.keymem.key_mem[7][114] ),
    .B(_12048_),
    .S(_14964_),
    .Z(_02389_));
 MUX2_X1 _39118_ (.A(\core.keymem.key_mem[7][115] ),
    .B(_12058_),
    .S(_14964_),
    .Z(_02390_));
 BUF_X4 _39119_ (.A(_14956_),
    .Z(_14966_));
 MUX2_X1 _39120_ (.A(\core.keymem.key_mem[7][116] ),
    .B(_12076_),
    .S(_14966_),
    .Z(_02391_));
 MUX2_X1 _39121_ (.A(\core.keymem.key_mem[7][117] ),
    .B(_12877_),
    .S(_14966_),
    .Z(_02392_));
 MUX2_X1 _39122_ (.A(\core.keymem.key_mem[7][118] ),
    .B(_12882_),
    .S(_14966_),
    .Z(_02393_));
 MUX2_X1 _39123_ (.A(\core.keymem.key_mem[7][119] ),
    .B(_12095_),
    .S(_14966_),
    .Z(_02394_));
 NAND2_X1 _39124_ (.A1(\core.keymem.key_mem[7][11] ),
    .A2(_14960_),
    .ZN(_14967_));
 OAI21_X1 _39125_ (.A(_14967_),
    .B1(_14963_),
    .B2(_12895_),
    .ZN(_02395_));
 MUX2_X1 _39126_ (.A(\core.keymem.key_mem[7][120] ),
    .B(_12123_),
    .S(_14966_),
    .Z(_02396_));
 MUX2_X1 _39127_ (.A(\core.keymem.key_mem[7][121] ),
    .B(_12159_),
    .S(_14966_),
    .Z(_02397_));
 MUX2_X1 _39128_ (.A(\core.keymem.key_mem[7][122] ),
    .B(_12902_),
    .S(_14966_),
    .Z(_02398_));
 NAND2_X1 _39129_ (.A1(\core.keymem.key_mem[7][123] ),
    .A2(_14960_),
    .ZN(_14968_));
 OAI21_X1 _39130_ (.A(_14968_),
    .B1(_14963_),
    .B2(_12181_),
    .ZN(_02399_));
 NAND2_X1 _39131_ (.A1(\core.keymem.key_mem[7][124] ),
    .A2(_14960_),
    .ZN(_14969_));
 OAI21_X1 _39132_ (.A(_14969_),
    .B1(_14963_),
    .B2(_12925_),
    .ZN(_02400_));
 MUX2_X1 _39133_ (.A(\core.keymem.key_mem[7][125] ),
    .B(_12931_),
    .S(_14966_),
    .Z(_02401_));
 NAND2_X1 _39134_ (.A1(\core.keymem.key_mem[7][126] ),
    .A2(_14960_),
    .ZN(_14970_));
 OAI21_X1 _39135_ (.A(_14970_),
    .B1(_14963_),
    .B2(_12206_),
    .ZN(_02402_));
 MUX2_X1 _39136_ (.A(\core.keymem.key_mem[7][127] ),
    .B(_12944_),
    .S(_14966_),
    .Z(_02403_));
 MUX2_X1 _39137_ (.A(\core.keymem.key_mem[7][12] ),
    .B(_12958_),
    .S(_14966_),
    .Z(_02404_));
 BUF_X4 _39138_ (.A(_14955_),
    .Z(_14971_));
 MUX2_X1 _39139_ (.A(\core.keymem.key_mem[7][13] ),
    .B(_12974_),
    .S(_14971_),
    .Z(_02405_));
 NOR2_X1 _39140_ (.A1(\core.keymem.key_mem[7][14] ),
    .A2(_14957_),
    .ZN(_14972_));
 AOI21_X1 _39141_ (.A(_14972_),
    .B1(_14957_),
    .B2(_13007_),
    .ZN(_02406_));
 MUX2_X1 _39142_ (.A(\core.keymem.key_mem[7][15] ),
    .B(_13017_),
    .S(_14971_),
    .Z(_02407_));
 MUX2_X1 _39143_ (.A(\core.keymem.key_mem[7][16] ),
    .B(_13029_),
    .S(_14971_),
    .Z(_02408_));
 NAND2_X1 _39144_ (.A1(\core.keymem.key_mem[7][17] ),
    .A2(_14960_),
    .ZN(_14973_));
 OAI21_X1 _39145_ (.A(_14973_),
    .B1(_14963_),
    .B2(_13042_),
    .ZN(_02409_));
 MUX2_X1 _39146_ (.A(\core.keymem.key_mem[7][18] ),
    .B(_13094_),
    .S(_14971_),
    .Z(_02410_));
 BUF_X4 _39147_ (.A(_14959_),
    .Z(_14974_));
 NAND2_X1 _39148_ (.A1(\core.keymem.key_mem[7][19] ),
    .A2(_14974_),
    .ZN(_14975_));
 OAI21_X1 _39149_ (.A(_14975_),
    .B1(_14963_),
    .B2(_13109_),
    .ZN(_02411_));
 MUX2_X1 _39150_ (.A(\core.keymem.key_mem[7][1] ),
    .B(_13134_),
    .S(_14971_),
    .Z(_02412_));
 MUX2_X1 _39151_ (.A(\core.keymem.key_mem[7][20] ),
    .B(_13146_),
    .S(_14971_),
    .Z(_02413_));
 MUX2_X1 _39152_ (.A(\core.keymem.key_mem[7][21] ),
    .B(_13155_),
    .S(_14971_),
    .Z(_02414_));
 NOR2_X1 _39153_ (.A1(\core.keymem.key_mem[7][22] ),
    .A2(_14957_),
    .ZN(_14976_));
 AOI21_X1 _39154_ (.A(_14976_),
    .B1(_14957_),
    .B2(_13191_),
    .ZN(_02415_));
 MUX2_X1 _39155_ (.A(\core.keymem.key_mem[7][23] ),
    .B(_13196_),
    .S(_14971_),
    .Z(_02416_));
 NAND2_X1 _39156_ (.A1(\core.keymem.key_mem[7][24] ),
    .A2(_14974_),
    .ZN(_14977_));
 OAI21_X1 _39157_ (.A(_14977_),
    .B1(_14963_),
    .B2(_13211_),
    .ZN(_02417_));
 MUX2_X1 _39158_ (.A(\core.keymem.key_mem[7][25] ),
    .B(_13233_),
    .S(_14971_),
    .Z(_02418_));
 MUX2_X1 _39159_ (.A(\core.keymem.key_mem[7][26] ),
    .B(_13240_),
    .S(_14971_),
    .Z(_02419_));
 BUF_X4 _39160_ (.A(_14955_),
    .Z(_14978_));
 MUX2_X1 _39161_ (.A(\core.keymem.key_mem[7][27] ),
    .B(_13283_),
    .S(_14978_),
    .Z(_02420_));
 MUX2_X1 _39162_ (.A(\core.keymem.key_mem[7][28] ),
    .B(_13324_),
    .S(_14978_),
    .Z(_02421_));
 MUX2_X1 _39163_ (.A(\core.keymem.key_mem[7][29] ),
    .B(_13328_),
    .S(_14978_),
    .Z(_02422_));
 NAND2_X1 _39164_ (.A1(\core.keymem.key_mem[7][2] ),
    .A2(_14974_),
    .ZN(_14979_));
 OAI21_X1 _39165_ (.A(_14979_),
    .B1(_14963_),
    .B2(_13335_),
    .ZN(_02423_));
 MUX2_X1 _39166_ (.A(\core.keymem.key_mem[7][30] ),
    .B(_13378_),
    .S(_14978_),
    .Z(_02424_));
 MUX2_X1 _39167_ (.A(\core.keymem.key_mem[7][31] ),
    .B(_13394_),
    .S(_14978_),
    .Z(_02425_));
 MUX2_X1 _39168_ (.A(\core.keymem.key_mem[7][32] ),
    .B(_12354_),
    .S(_14978_),
    .Z(_02426_));
 MUX2_X1 _39169_ (.A(\core.keymem.key_mem[7][33] ),
    .B(_13401_),
    .S(_14978_),
    .Z(_02427_));
 MUX2_X1 _39170_ (.A(\core.keymem.key_mem[7][34] ),
    .B(_12375_),
    .S(_14978_),
    .Z(_02428_));
 MUX2_X1 _39171_ (.A(\core.keymem.key_mem[7][35] ),
    .B(_13404_),
    .S(_14978_),
    .Z(_02429_));
 NAND2_X1 _39172_ (.A1(\core.keymem.key_mem[7][36] ),
    .A2(_14974_),
    .ZN(_14980_));
 BUF_X4 _39173_ (.A(_14962_),
    .Z(_14981_));
 OAI21_X1 _39174_ (.A(_14980_),
    .B1(_14981_),
    .B2(_12422_),
    .ZN(_02430_));
 NAND2_X1 _39175_ (.A1(\core.keymem.key_mem[7][37] ),
    .A2(_14974_),
    .ZN(_14982_));
 OAI21_X1 _39176_ (.A(_14982_),
    .B1(_14981_),
    .B2(_12438_),
    .ZN(_02431_));
 MUX2_X1 _39177_ (.A(\core.keymem.key_mem[7][38] ),
    .B(_13409_),
    .S(_14978_),
    .Z(_02432_));
 NAND2_X1 _39178_ (.A1(\core.keymem.key_mem[7][39] ),
    .A2(_14974_),
    .ZN(_14983_));
 OAI21_X1 _39179_ (.A(_14983_),
    .B1(_14981_),
    .B2(_13434_),
    .ZN(_02433_));
 NAND2_X1 _39180_ (.A1(\core.keymem.key_mem[7][3] ),
    .A2(_14974_),
    .ZN(_14984_));
 OAI21_X1 _39181_ (.A(_14984_),
    .B1(_14981_),
    .B2(_13448_),
    .ZN(_02434_));
 NAND2_X1 _39182_ (.A1(\core.keymem.key_mem[7][40] ),
    .A2(_14974_),
    .ZN(_14985_));
 OAI21_X1 _39183_ (.A(_14985_),
    .B1(_14981_),
    .B2(_13456_),
    .ZN(_02435_));
 BUF_X4 _39184_ (.A(_14955_),
    .Z(_14986_));
 MUX2_X1 _39185_ (.A(\core.keymem.key_mem[7][41] ),
    .B(_13466_),
    .S(_14986_),
    .Z(_02436_));
 MUX2_X1 _39186_ (.A(\core.keymem.key_mem[7][42] ),
    .B(_13490_),
    .S(_14986_),
    .Z(_02437_));
 NAND2_X1 _39187_ (.A1(\core.keymem.key_mem[7][43] ),
    .A2(_14974_),
    .ZN(_14987_));
 OAI21_X1 _39188_ (.A(_14987_),
    .B1(_14981_),
    .B2(_13496_),
    .ZN(_02438_));
 MUX2_X1 _39189_ (.A(\core.keymem.key_mem[7][44] ),
    .B(_12505_),
    .S(_14986_),
    .Z(_02439_));
 NAND2_X1 _39190_ (.A1(\core.keymem.key_mem[7][45] ),
    .A2(_14974_),
    .ZN(_14988_));
 OAI21_X1 _39191_ (.A(_14988_),
    .B1(_14981_),
    .B2(_13510_),
    .ZN(_02440_));
 BUF_X4 _39192_ (.A(_14959_),
    .Z(_14989_));
 NAND2_X1 _39193_ (.A1(\core.keymem.key_mem[7][46] ),
    .A2(_14989_),
    .ZN(_14990_));
 OAI21_X1 _39194_ (.A(_14990_),
    .B1(_14981_),
    .B2(_13517_),
    .ZN(_02441_));
 NAND2_X1 _39195_ (.A1(\core.keymem.key_mem[7][47] ),
    .A2(_14989_),
    .ZN(_14991_));
 OAI21_X1 _39196_ (.A(_14991_),
    .B1(_14981_),
    .B2(_12519_),
    .ZN(_02442_));
 NAND2_X1 _39197_ (.A1(\core.keymem.key_mem[7][48] ),
    .A2(_14989_),
    .ZN(_14992_));
 OAI21_X1 _39198_ (.A(_14992_),
    .B1(_14981_),
    .B2(_12531_),
    .ZN(_02443_));
 NAND2_X1 _39199_ (.A1(\core.keymem.key_mem[7][49] ),
    .A2(_14989_),
    .ZN(_14993_));
 BUF_X4 _39200_ (.A(_14962_),
    .Z(_14994_));
 OAI21_X1 _39201_ (.A(_14993_),
    .B1(_14994_),
    .B2(_13528_),
    .ZN(_02444_));
 MUX2_X1 _39202_ (.A(\core.keymem.key_mem[7][4] ),
    .B(_13538_),
    .S(_14986_),
    .Z(_02445_));
 MUX2_X1 _39203_ (.A(\core.keymem.key_mem[7][50] ),
    .B(_13557_),
    .S(_14986_),
    .Z(_02446_));
 MUX2_X1 _39204_ (.A(\core.keymem.key_mem[7][51] ),
    .B(_13563_),
    .S(_14986_),
    .Z(_02447_));
 NAND2_X1 _39205_ (.A1(\core.keymem.key_mem[7][52] ),
    .A2(_14989_),
    .ZN(_14995_));
 OAI21_X1 _39206_ (.A(_14995_),
    .B1(_14994_),
    .B2(_12567_),
    .ZN(_02448_));
 NAND2_X1 _39207_ (.A1(\core.keymem.key_mem[7][53] ),
    .A2(_14989_),
    .ZN(_14996_));
 OAI21_X1 _39208_ (.A(_14996_),
    .B1(_14994_),
    .B2(_12583_),
    .ZN(_02449_));
 NAND2_X1 _39209_ (.A1(\core.keymem.key_mem[7][54] ),
    .A2(_14989_),
    .ZN(_14997_));
 OAI21_X1 _39210_ (.A(_14997_),
    .B1(_14994_),
    .B2(_13574_),
    .ZN(_02450_));
 MUX2_X1 _39211_ (.A(\core.keymem.key_mem[7][55] ),
    .B(_13581_),
    .S(_14986_),
    .Z(_02451_));
 MUX2_X1 _39212_ (.A(\core.keymem.key_mem[7][56] ),
    .B(_13589_),
    .S(_14986_),
    .Z(_02452_));
 MUX2_X1 _39213_ (.A(\core.keymem.key_mem[7][57] ),
    .B(_13604_),
    .S(_14986_),
    .Z(_02453_));
 MUX2_X1 _39214_ (.A(\core.keymem.key_mem[7][58] ),
    .B(_13611_),
    .S(_14986_),
    .Z(_02454_));
 BUF_X4 _39215_ (.A(_14955_),
    .Z(_14998_));
 MUX2_X1 _39216_ (.A(\core.keymem.key_mem[7][59] ),
    .B(_13616_),
    .S(_14998_),
    .Z(_02455_));
 MUX2_X1 _39217_ (.A(\core.keymem.key_mem[7][5] ),
    .B(_12605_),
    .S(_14998_),
    .Z(_02456_));
 MUX2_X1 _39218_ (.A(\core.keymem.key_mem[7][60] ),
    .B(_13622_),
    .S(_14998_),
    .Z(_02457_));
 MUX2_X1 _39219_ (.A(\core.keymem.key_mem[7][61] ),
    .B(_13632_),
    .S(_14998_),
    .Z(_02458_));
 MUX2_X1 _39220_ (.A(\core.keymem.key_mem[7][62] ),
    .B(_13636_),
    .S(_14998_),
    .Z(_02459_));
 MUX2_X1 _39221_ (.A(\core.keymem.key_mem[7][63] ),
    .B(_13659_),
    .S(_14998_),
    .Z(_02460_));
 MUX2_X1 _39222_ (.A(\core.keymem.key_mem[7][64] ),
    .B(_12621_),
    .S(_14998_),
    .Z(_02461_));
 NAND2_X1 _39223_ (.A1(\core.keymem.key_mem[7][65] ),
    .A2(_14989_),
    .ZN(_14999_));
 OAI21_X1 _39224_ (.A(_14999_),
    .B1(_14994_),
    .B2(_13672_),
    .ZN(_02462_));
 MUX2_X1 _39225_ (.A(\core.keymem.key_mem[7][66] ),
    .B(_13680_),
    .S(_14998_),
    .Z(_02463_));
 NAND2_X1 _39226_ (.A1(\core.keymem.key_mem[7][67] ),
    .A2(_14989_),
    .ZN(_15000_));
 OAI21_X1 _39227_ (.A(_15000_),
    .B1(_14994_),
    .B2(_13689_),
    .ZN(_02464_));
 NAND2_X1 _39228_ (.A1(\core.keymem.key_mem[7][68] ),
    .A2(_14989_),
    .ZN(_15001_));
 OAI21_X1 _39229_ (.A(_15001_),
    .B1(_14994_),
    .B2(_12634_),
    .ZN(_02465_));
 BUF_X4 _39230_ (.A(_14959_),
    .Z(_15002_));
 NAND2_X1 _39231_ (.A1(\core.keymem.key_mem[7][69] ),
    .A2(_15002_),
    .ZN(_15003_));
 OAI21_X1 _39232_ (.A(_15003_),
    .B1(_14994_),
    .B2(_13699_),
    .ZN(_02466_));
 MUX2_X1 _39233_ (.A(\core.keymem.key_mem[7][6] ),
    .B(_13710_),
    .S(_14998_),
    .Z(_02467_));
 MUX2_X1 _39234_ (.A(\core.keymem.key_mem[7][70] ),
    .B(_13712_),
    .S(_14998_),
    .Z(_02468_));
 NAND2_X1 _39235_ (.A1(\core.keymem.key_mem[7][71] ),
    .A2(_15002_),
    .ZN(_15004_));
 OAI21_X1 _39236_ (.A(_15004_),
    .B1(_14994_),
    .B2(_12658_),
    .ZN(_02469_));
 NAND2_X1 _39237_ (.A1(\core.keymem.key_mem[7][72] ),
    .A2(_15002_),
    .ZN(_15005_));
 OAI21_X1 _39238_ (.A(_15005_),
    .B1(_14994_),
    .B2(_12673_),
    .ZN(_02470_));
 NAND2_X1 _39239_ (.A1(\core.keymem.key_mem[7][73] ),
    .A2(_15002_),
    .ZN(_15006_));
 BUF_X4 _39240_ (.A(_14962_),
    .Z(_15007_));
 OAI21_X1 _39241_ (.A(_15006_),
    .B1(_15007_),
    .B2(_12687_),
    .ZN(_02471_));
 NAND2_X1 _39242_ (.A1(\core.keymem.key_mem[7][74] ),
    .A2(_15002_),
    .ZN(_15008_));
 OAI21_X1 _39243_ (.A(_15008_),
    .B1(_15007_),
    .B2(_13726_),
    .ZN(_02472_));
 NAND2_X1 _39244_ (.A1(\core.keymem.key_mem[7][75] ),
    .A2(_15002_),
    .ZN(_15009_));
 OAI21_X1 _39245_ (.A(_15009_),
    .B1(_15007_),
    .B2(_13732_),
    .ZN(_02473_));
 BUF_X4 _39246_ (.A(_14955_),
    .Z(_15010_));
 MUX2_X1 _39247_ (.A(\core.keymem.key_mem[7][76] ),
    .B(_13740_),
    .S(_15010_),
    .Z(_02474_));
 MUX2_X1 _39248_ (.A(\core.keymem.key_mem[7][77] ),
    .B(_13751_),
    .S(_15010_),
    .Z(_02475_));
 NAND2_X1 _39249_ (.A1(\core.keymem.key_mem[7][78] ),
    .A2(_15002_),
    .ZN(_15011_));
 OAI21_X1 _39250_ (.A(_15011_),
    .B1(_15007_),
    .B2(_12707_),
    .ZN(_02476_));
 MUX2_X1 _39251_ (.A(\core.keymem.key_mem[7][79] ),
    .B(_13758_),
    .S(_15010_),
    .Z(_02477_));
 NAND2_X1 _39252_ (.A1(\core.keymem.key_mem[7][7] ),
    .A2(_15002_),
    .ZN(_15012_));
 OAI21_X1 _39253_ (.A(_15012_),
    .B1(_15007_),
    .B2(_13766_),
    .ZN(_02478_));
 MUX2_X1 _39254_ (.A(\core.keymem.key_mem[7][80] ),
    .B(_13768_),
    .S(_15010_),
    .Z(_02479_));
 NAND2_X1 _39255_ (.A1(\core.keymem.key_mem[7][81] ),
    .A2(_15002_),
    .ZN(_15013_));
 OAI21_X1 _39256_ (.A(_15013_),
    .B1(_15007_),
    .B2(_13774_),
    .ZN(_02480_));
 NAND2_X1 _39257_ (.A1(\core.keymem.key_mem[7][82] ),
    .A2(_15002_),
    .ZN(_15014_));
 OAI21_X1 _39258_ (.A(_15014_),
    .B1(_15007_),
    .B2(_13782_),
    .ZN(_02481_));
 NAND2_X1 _39259_ (.A1(\core.keymem.key_mem[7][83] ),
    .A2(_14962_),
    .ZN(_15015_));
 OAI21_X1 _39260_ (.A(_15015_),
    .B1(_15007_),
    .B2(_13790_),
    .ZN(_02482_));
 NAND2_X1 _39261_ (.A1(\core.keymem.key_mem[7][84] ),
    .A2(_14962_),
    .ZN(_15016_));
 OAI21_X1 _39262_ (.A(_15016_),
    .B1(_15007_),
    .B2(_12724_),
    .ZN(_02483_));
 MUX2_X1 _39263_ (.A(\core.keymem.key_mem[7][85] ),
    .B(_13798_),
    .S(_15010_),
    .Z(_02484_));
 MUX2_X1 _39264_ (.A(\core.keymem.key_mem[7][86] ),
    .B(_12740_),
    .S(_15010_),
    .Z(_02485_));
 MUX2_X1 _39265_ (.A(\core.keymem.key_mem[7][87] ),
    .B(_13804_),
    .S(_15010_),
    .Z(_02486_));
 MUX2_X1 _39266_ (.A(\core.keymem.key_mem[7][88] ),
    .B(_13810_),
    .S(_15010_),
    .Z(_02487_));
 MUX2_X1 _39267_ (.A(\core.keymem.key_mem[7][89] ),
    .B(_13818_),
    .S(_15010_),
    .Z(_02488_));
 MUX2_X1 _39268_ (.A(\core.keymem.key_mem[7][8] ),
    .B(_13854_),
    .S(_15010_),
    .Z(_02489_));
 MUX2_X1 _39269_ (.A(\core.keymem.key_mem[7][90] ),
    .B(_13860_),
    .S(_14956_),
    .Z(_02490_));
 NAND2_X1 _39270_ (.A1(\core.keymem.key_mem[7][91] ),
    .A2(_14962_),
    .ZN(_15017_));
 OAI21_X1 _39271_ (.A(_15017_),
    .B1(_15007_),
    .B2(_13870_),
    .ZN(_02491_));
 NAND2_X1 _39272_ (.A1(\core.keymem.key_mem[7][92] ),
    .A2(_14962_),
    .ZN(_15018_));
 OAI21_X1 _39273_ (.A(_15018_),
    .B1(_14960_),
    .B2(_13880_),
    .ZN(_02492_));
 MUX2_X1 _39274_ (.A(\core.keymem.key_mem[7][93] ),
    .B(_13889_),
    .S(_14956_),
    .Z(_02493_));
 MUX2_X1 _39275_ (.A(\core.keymem.key_mem[7][94] ),
    .B(_13896_),
    .S(_14956_),
    .Z(_02494_));
 MUX2_X1 _39276_ (.A(\core.keymem.key_mem[7][95] ),
    .B(_13903_),
    .S(_14956_),
    .Z(_02495_));
 MUX2_X1 _39277_ (.A(\core.keymem.key_mem[7][96] ),
    .B(_13907_),
    .S(_14956_),
    .Z(_02496_));
 NAND2_X1 _39278_ (.A1(\core.keymem.key_mem[7][97] ),
    .A2(_14962_),
    .ZN(_15019_));
 OAI21_X1 _39279_ (.A(_15019_),
    .B1(_14960_),
    .B2(_12776_),
    .ZN(_02497_));
 NAND2_X1 _39280_ (.A1(\core.keymem.key_mem[7][98] ),
    .A2(_14962_),
    .ZN(_15020_));
 OAI21_X1 _39281_ (.A(_15020_),
    .B1(_14960_),
    .B2(_12787_),
    .ZN(_02498_));
 MUX2_X1 _39282_ (.A(\core.keymem.key_mem[7][99] ),
    .B(_12799_),
    .S(_14956_),
    .Z(_02499_));
 MUX2_X1 _39283_ (.A(\core.keymem.key_mem[7][9] ),
    .B(_13919_),
    .S(_14956_),
    .Z(_02500_));
 NOR2_X4 _39284_ (.A1(_12803_),
    .A2(_13989_),
    .ZN(_15021_));
 BUF_X4 _39285_ (.A(_15021_),
    .Z(_15022_));
 BUF_X4 _39286_ (.A(_15022_),
    .Z(_15023_));
 MUX2_X1 _39287_ (.A(\core.keymem.key_mem[8][0] ),
    .B(_11843_),
    .S(_15023_),
    .Z(_02501_));
 MUX2_X1 _39288_ (.A(\core.keymem.key_mem[8][100] ),
    .B(_11872_),
    .S(_15023_),
    .Z(_02502_));
 MUX2_X1 _39289_ (.A(\core.keymem.key_mem[8][101] ),
    .B(_12813_),
    .S(_15023_),
    .Z(_02503_));
 MUX2_X1 _39290_ (.A(\core.keymem.key_mem[8][102] ),
    .B(_11905_),
    .S(_15023_),
    .Z(_02504_));
 MUX2_X1 _39291_ (.A(\core.keymem.key_mem[8][103] ),
    .B(_11928_),
    .S(_15023_),
    .Z(_02505_));
 OR2_X1 _39292_ (.A1(_12803_),
    .A2(_13989_),
    .ZN(_15024_));
 CLKBUF_X3 _39293_ (.A(_15024_),
    .Z(_15025_));
 BUF_X4 _39294_ (.A(_15025_),
    .Z(_15026_));
 NAND2_X1 _39295_ (.A1(\core.keymem.key_mem[8][104] ),
    .A2(_15026_),
    .ZN(_15027_));
 BUF_X4 _39296_ (.A(_15025_),
    .Z(_15028_));
 BUF_X4 _39297_ (.A(_15028_),
    .Z(_15029_));
 OAI21_X1 _39298_ (.A(_15027_),
    .B1(_15029_),
    .B2(_12822_),
    .ZN(_02506_));
 MUX2_X1 _39299_ (.A(\core.keymem.key_mem[8][105] ),
    .B(_12829_),
    .S(_15023_),
    .Z(_02507_));
 BUF_X4 _39300_ (.A(_15022_),
    .Z(_15030_));
 MUX2_X1 _39301_ (.A(\core.keymem.key_mem[8][106] ),
    .B(_12831_),
    .S(_15030_),
    .Z(_02508_));
 MUX2_X1 _39302_ (.A(\core.keymem.key_mem[8][107] ),
    .B(_11966_),
    .S(_15030_),
    .Z(_02509_));
 MUX2_X1 _39303_ (.A(\core.keymem.key_mem[8][108] ),
    .B(_11980_),
    .S(_15030_),
    .Z(_02510_));
 MUX2_X1 _39304_ (.A(\core.keymem.key_mem[8][109] ),
    .B(_12841_),
    .S(_15030_),
    .Z(_02511_));
 NAND2_X1 _39305_ (.A1(\core.keymem.key_mem[8][10] ),
    .A2(_15026_),
    .ZN(_15031_));
 OAI21_X1 _39306_ (.A(_15031_),
    .B1(_15029_),
    .B2(_12858_),
    .ZN(_02512_));
 MUX2_X1 _39307_ (.A(\core.keymem.key_mem[8][110] ),
    .B(_12003_),
    .S(_15030_),
    .Z(_02513_));
 MUX2_X1 _39308_ (.A(\core.keymem.key_mem[8][111] ),
    .B(_12016_),
    .S(_15030_),
    .Z(_02514_));
 MUX2_X1 _39309_ (.A(\core.keymem.key_mem[8][112] ),
    .B(_12030_),
    .S(_15030_),
    .Z(_02515_));
 MUX2_X1 _39310_ (.A(\core.keymem.key_mem[8][113] ),
    .B(_12868_),
    .S(_15030_),
    .Z(_02516_));
 MUX2_X1 _39311_ (.A(\core.keymem.key_mem[8][114] ),
    .B(_12048_),
    .S(_15030_),
    .Z(_02517_));
 MUX2_X1 _39312_ (.A(\core.keymem.key_mem[8][115] ),
    .B(_12058_),
    .S(_15030_),
    .Z(_02518_));
 BUF_X4 _39313_ (.A(_15022_),
    .Z(_15032_));
 MUX2_X1 _39314_ (.A(\core.keymem.key_mem[8][116] ),
    .B(_12076_),
    .S(_15032_),
    .Z(_02519_));
 MUX2_X1 _39315_ (.A(\core.keymem.key_mem[8][117] ),
    .B(_12877_),
    .S(_15032_),
    .Z(_02520_));
 MUX2_X1 _39316_ (.A(\core.keymem.key_mem[8][118] ),
    .B(_12882_),
    .S(_15032_),
    .Z(_02521_));
 MUX2_X1 _39317_ (.A(\core.keymem.key_mem[8][119] ),
    .B(_12095_),
    .S(_15032_),
    .Z(_02522_));
 NAND2_X1 _39318_ (.A1(\core.keymem.key_mem[8][11] ),
    .A2(_15026_),
    .ZN(_15033_));
 OAI21_X1 _39319_ (.A(_15033_),
    .B1(_15029_),
    .B2(_12895_),
    .ZN(_02523_));
 MUX2_X1 _39320_ (.A(\core.keymem.key_mem[8][120] ),
    .B(_12123_),
    .S(_15032_),
    .Z(_02524_));
 MUX2_X1 _39321_ (.A(\core.keymem.key_mem[8][121] ),
    .B(_12159_),
    .S(_15032_),
    .Z(_02525_));
 MUX2_X1 _39322_ (.A(\core.keymem.key_mem[8][122] ),
    .B(_12902_),
    .S(_15032_),
    .Z(_02526_));
 NAND2_X1 _39323_ (.A1(\core.keymem.key_mem[8][123] ),
    .A2(_15026_),
    .ZN(_15034_));
 OAI21_X1 _39324_ (.A(_15034_),
    .B1(_15029_),
    .B2(_12181_),
    .ZN(_02527_));
 NAND2_X1 _39325_ (.A1(\core.keymem.key_mem[8][124] ),
    .A2(_15026_),
    .ZN(_15035_));
 OAI21_X1 _39326_ (.A(_15035_),
    .B1(_15029_),
    .B2(_12925_),
    .ZN(_02528_));
 MUX2_X1 _39327_ (.A(\core.keymem.key_mem[8][125] ),
    .B(_12931_),
    .S(_15032_),
    .Z(_02529_));
 NAND2_X1 _39328_ (.A1(\core.keymem.key_mem[8][126] ),
    .A2(_15026_),
    .ZN(_15036_));
 OAI21_X1 _39329_ (.A(_15036_),
    .B1(_15029_),
    .B2(_12206_),
    .ZN(_02530_));
 MUX2_X1 _39330_ (.A(\core.keymem.key_mem[8][127] ),
    .B(_12944_),
    .S(_15032_),
    .Z(_02531_));
 MUX2_X1 _39331_ (.A(\core.keymem.key_mem[8][12] ),
    .B(_12958_),
    .S(_15032_),
    .Z(_02532_));
 BUF_X4 _39332_ (.A(_15021_),
    .Z(_15037_));
 MUX2_X1 _39333_ (.A(\core.keymem.key_mem[8][13] ),
    .B(_12974_),
    .S(_15037_),
    .Z(_02533_));
 NOR2_X1 _39334_ (.A1(\core.keymem.key_mem[8][14] ),
    .A2(_15023_),
    .ZN(_15038_));
 AOI21_X1 _39335_ (.A(_15038_),
    .B1(_15023_),
    .B2(_13007_),
    .ZN(_02534_));
 MUX2_X1 _39336_ (.A(\core.keymem.key_mem[8][15] ),
    .B(_13017_),
    .S(_15037_),
    .Z(_02535_));
 MUX2_X1 _39337_ (.A(\core.keymem.key_mem[8][16] ),
    .B(_13028_),
    .S(_15037_),
    .Z(_02536_));
 NAND2_X1 _39338_ (.A1(\core.keymem.key_mem[8][17] ),
    .A2(_15026_),
    .ZN(_15039_));
 OAI21_X1 _39339_ (.A(_15039_),
    .B1(_15029_),
    .B2(_13042_),
    .ZN(_02537_));
 MUX2_X1 _39340_ (.A(\core.keymem.key_mem[8][18] ),
    .B(_13093_),
    .S(_15037_),
    .Z(_02538_));
 BUF_X4 _39341_ (.A(_15025_),
    .Z(_15040_));
 NAND2_X1 _39342_ (.A1(\core.keymem.key_mem[8][19] ),
    .A2(_15040_),
    .ZN(_15041_));
 OAI21_X1 _39343_ (.A(_15041_),
    .B1(_15029_),
    .B2(_13109_),
    .ZN(_02539_));
 MUX2_X1 _39344_ (.A(\core.keymem.key_mem[8][1] ),
    .B(_13134_),
    .S(_15037_),
    .Z(_02540_));
 MUX2_X1 _39345_ (.A(\core.keymem.key_mem[8][20] ),
    .B(_13146_),
    .S(_15037_),
    .Z(_02541_));
 MUX2_X1 _39346_ (.A(\core.keymem.key_mem[8][21] ),
    .B(_13155_),
    .S(_15037_),
    .Z(_02542_));
 NOR2_X1 _39347_ (.A1(\core.keymem.key_mem[8][22] ),
    .A2(_15023_),
    .ZN(_15042_));
 AOI21_X1 _39348_ (.A(_15042_),
    .B1(_15023_),
    .B2(_13191_),
    .ZN(_02543_));
 MUX2_X1 _39349_ (.A(\core.keymem.key_mem[8][23] ),
    .B(_13196_),
    .S(_15037_),
    .Z(_02544_));
 NAND2_X1 _39350_ (.A1(\core.keymem.key_mem[8][24] ),
    .A2(_15040_),
    .ZN(_15043_));
 OAI21_X1 _39351_ (.A(_15043_),
    .B1(_15029_),
    .B2(_13211_),
    .ZN(_02545_));
 MUX2_X1 _39352_ (.A(\core.keymem.key_mem[8][25] ),
    .B(_13232_),
    .S(_15037_),
    .Z(_02546_));
 MUX2_X1 _39353_ (.A(\core.keymem.key_mem[8][26] ),
    .B(_13240_),
    .S(_15037_),
    .Z(_02547_));
 BUF_X4 _39354_ (.A(_15021_),
    .Z(_15044_));
 MUX2_X1 _39355_ (.A(\core.keymem.key_mem[8][27] ),
    .B(_13283_),
    .S(_15044_),
    .Z(_02548_));
 MUX2_X1 _39356_ (.A(\core.keymem.key_mem[8][28] ),
    .B(_13324_),
    .S(_15044_),
    .Z(_02549_));
 MUX2_X1 _39357_ (.A(\core.keymem.key_mem[8][29] ),
    .B(_13328_),
    .S(_15044_),
    .Z(_02550_));
 NAND2_X1 _39358_ (.A1(\core.keymem.key_mem[8][2] ),
    .A2(_15040_),
    .ZN(_15045_));
 OAI21_X1 _39359_ (.A(_15045_),
    .B1(_15029_),
    .B2(_13335_),
    .ZN(_02551_));
 MUX2_X1 _39360_ (.A(\core.keymem.key_mem[8][30] ),
    .B(_13378_),
    .S(_15044_),
    .Z(_02552_));
 MUX2_X1 _39361_ (.A(\core.keymem.key_mem[8][31] ),
    .B(_13394_),
    .S(_15044_),
    .Z(_02553_));
 MUX2_X1 _39362_ (.A(\core.keymem.key_mem[8][32] ),
    .B(_12354_),
    .S(_15044_),
    .Z(_02554_));
 MUX2_X1 _39363_ (.A(\core.keymem.key_mem[8][33] ),
    .B(_13401_),
    .S(_15044_),
    .Z(_02555_));
 MUX2_X1 _39364_ (.A(\core.keymem.key_mem[8][34] ),
    .B(_12375_),
    .S(_15044_),
    .Z(_02556_));
 MUX2_X1 _39365_ (.A(\core.keymem.key_mem[8][35] ),
    .B(_13404_),
    .S(_15044_),
    .Z(_02557_));
 NAND2_X1 _39366_ (.A1(\core.keymem.key_mem[8][36] ),
    .A2(_15040_),
    .ZN(_15046_));
 BUF_X4 _39367_ (.A(_15028_),
    .Z(_15047_));
 OAI21_X1 _39368_ (.A(_15046_),
    .B1(_15047_),
    .B2(_12422_),
    .ZN(_02558_));
 NAND2_X1 _39369_ (.A1(\core.keymem.key_mem[8][37] ),
    .A2(_15040_),
    .ZN(_15048_));
 OAI21_X1 _39370_ (.A(_15048_),
    .B1(_15047_),
    .B2(_12438_),
    .ZN(_02559_));
 MUX2_X1 _39371_ (.A(\core.keymem.key_mem[8][38] ),
    .B(_13409_),
    .S(_15044_),
    .Z(_02560_));
 NAND2_X1 _39372_ (.A1(\core.keymem.key_mem[8][39] ),
    .A2(_15040_),
    .ZN(_15049_));
 OAI21_X1 _39373_ (.A(_15049_),
    .B1(_15047_),
    .B2(_13434_),
    .ZN(_02561_));
 NAND2_X1 _39374_ (.A1(\core.keymem.key_mem[8][3] ),
    .A2(_15040_),
    .ZN(_15050_));
 OAI21_X1 _39375_ (.A(_15050_),
    .B1(_15047_),
    .B2(_13448_),
    .ZN(_02562_));
 NAND2_X1 _39376_ (.A1(\core.keymem.key_mem[8][40] ),
    .A2(_15040_),
    .ZN(_15051_));
 OAI21_X1 _39377_ (.A(_15051_),
    .B1(_15047_),
    .B2(_13456_),
    .ZN(_02563_));
 BUF_X4 _39378_ (.A(_15021_),
    .Z(_15052_));
 MUX2_X1 _39379_ (.A(\core.keymem.key_mem[8][41] ),
    .B(_13466_),
    .S(_15052_),
    .Z(_02564_));
 MUX2_X1 _39380_ (.A(\core.keymem.key_mem[8][42] ),
    .B(_13490_),
    .S(_15052_),
    .Z(_02565_));
 NAND2_X1 _39381_ (.A1(\core.keymem.key_mem[8][43] ),
    .A2(_15040_),
    .ZN(_15053_));
 OAI21_X1 _39382_ (.A(_15053_),
    .B1(_15047_),
    .B2(_13495_),
    .ZN(_02566_));
 MUX2_X1 _39383_ (.A(\core.keymem.key_mem[8][44] ),
    .B(_12505_),
    .S(_15052_),
    .Z(_02567_));
 NAND2_X1 _39384_ (.A1(\core.keymem.key_mem[8][45] ),
    .A2(_15040_),
    .ZN(_15054_));
 OAI21_X1 _39385_ (.A(_15054_),
    .B1(_15047_),
    .B2(_13510_),
    .ZN(_02568_));
 BUF_X4 _39386_ (.A(_15025_),
    .Z(_15055_));
 NAND2_X1 _39387_ (.A1(\core.keymem.key_mem[8][46] ),
    .A2(_15055_),
    .ZN(_15056_));
 OAI21_X1 _39388_ (.A(_15056_),
    .B1(_15047_),
    .B2(_13516_),
    .ZN(_02569_));
 NAND2_X1 _39389_ (.A1(\core.keymem.key_mem[8][47] ),
    .A2(_15055_),
    .ZN(_15057_));
 OAI21_X1 _39390_ (.A(_15057_),
    .B1(_15047_),
    .B2(_12519_),
    .ZN(_02570_));
 NAND2_X1 _39391_ (.A1(\core.keymem.key_mem[8][48] ),
    .A2(_15055_),
    .ZN(_15058_));
 OAI21_X1 _39392_ (.A(_15058_),
    .B1(_15047_),
    .B2(_12531_),
    .ZN(_02571_));
 NAND2_X1 _39393_ (.A1(\core.keymem.key_mem[8][49] ),
    .A2(_15055_),
    .ZN(_15059_));
 BUF_X4 _39394_ (.A(_15028_),
    .Z(_15060_));
 OAI21_X1 _39395_ (.A(_15059_),
    .B1(_15060_),
    .B2(_13528_),
    .ZN(_02572_));
 MUX2_X1 _39396_ (.A(\core.keymem.key_mem[8][4] ),
    .B(_13538_),
    .S(_15052_),
    .Z(_02573_));
 MUX2_X1 _39397_ (.A(\core.keymem.key_mem[8][50] ),
    .B(_13557_),
    .S(_15052_),
    .Z(_02574_));
 MUX2_X1 _39398_ (.A(\core.keymem.key_mem[8][51] ),
    .B(_13563_),
    .S(_15052_),
    .Z(_02575_));
 NAND2_X1 _39399_ (.A1(\core.keymem.key_mem[8][52] ),
    .A2(_15055_),
    .ZN(_15061_));
 OAI21_X1 _39400_ (.A(_15061_),
    .B1(_15060_),
    .B2(_12567_),
    .ZN(_02576_));
 NAND2_X1 _39401_ (.A1(\core.keymem.key_mem[8][53] ),
    .A2(_15055_),
    .ZN(_15062_));
 OAI21_X1 _39402_ (.A(_15062_),
    .B1(_15060_),
    .B2(_12583_),
    .ZN(_02577_));
 NAND2_X1 _39403_ (.A1(\core.keymem.key_mem[8][54] ),
    .A2(_15055_),
    .ZN(_15063_));
 OAI21_X1 _39404_ (.A(_15063_),
    .B1(_15060_),
    .B2(_13574_),
    .ZN(_02578_));
 MUX2_X1 _39405_ (.A(\core.keymem.key_mem[8][55] ),
    .B(_13580_),
    .S(_15052_),
    .Z(_02579_));
 MUX2_X1 _39406_ (.A(\core.keymem.key_mem[8][56] ),
    .B(_13589_),
    .S(_15052_),
    .Z(_02580_));
 MUX2_X1 _39407_ (.A(\core.keymem.key_mem[8][57] ),
    .B(_13603_),
    .S(_15052_),
    .Z(_02581_));
 MUX2_X1 _39408_ (.A(\core.keymem.key_mem[8][58] ),
    .B(_13610_),
    .S(_15052_),
    .Z(_02582_));
 BUF_X4 _39409_ (.A(_15021_),
    .Z(_15064_));
 MUX2_X1 _39410_ (.A(\core.keymem.key_mem[8][59] ),
    .B(_13616_),
    .S(_15064_),
    .Z(_02583_));
 MUX2_X1 _39411_ (.A(\core.keymem.key_mem[8][5] ),
    .B(_12605_),
    .S(_15064_),
    .Z(_02584_));
 MUX2_X1 _39412_ (.A(\core.keymem.key_mem[8][60] ),
    .B(_13622_),
    .S(_15064_),
    .Z(_02585_));
 MUX2_X1 _39413_ (.A(\core.keymem.key_mem[8][61] ),
    .B(_13632_),
    .S(_15064_),
    .Z(_02586_));
 MUX2_X1 _39414_ (.A(\core.keymem.key_mem[8][62] ),
    .B(_13636_),
    .S(_15064_),
    .Z(_02587_));
 MUX2_X1 _39415_ (.A(\core.keymem.key_mem[8][63] ),
    .B(_13658_),
    .S(_15064_),
    .Z(_02588_));
 MUX2_X1 _39416_ (.A(\core.keymem.key_mem[8][64] ),
    .B(_12621_),
    .S(_15064_),
    .Z(_02589_));
 NAND2_X1 _39417_ (.A1(\core.keymem.key_mem[8][65] ),
    .A2(_15055_),
    .ZN(_15065_));
 OAI21_X1 _39418_ (.A(_15065_),
    .B1(_15060_),
    .B2(_13672_),
    .ZN(_02590_));
 MUX2_X1 _39419_ (.A(\core.keymem.key_mem[8][66] ),
    .B(_13680_),
    .S(_15064_),
    .Z(_02591_));
 NAND2_X1 _39420_ (.A1(\core.keymem.key_mem[8][67] ),
    .A2(_15055_),
    .ZN(_15066_));
 OAI21_X1 _39421_ (.A(_15066_),
    .B1(_15060_),
    .B2(_13689_),
    .ZN(_02592_));
 NAND2_X1 _39422_ (.A1(\core.keymem.key_mem[8][68] ),
    .A2(_15055_),
    .ZN(_15067_));
 OAI21_X1 _39423_ (.A(_15067_),
    .B1(_15060_),
    .B2(_12634_),
    .ZN(_02593_));
 BUF_X4 _39424_ (.A(_15025_),
    .Z(_15068_));
 NAND2_X1 _39425_ (.A1(\core.keymem.key_mem[8][69] ),
    .A2(_15068_),
    .ZN(_15069_));
 OAI21_X1 _39426_ (.A(_15069_),
    .B1(_15060_),
    .B2(_13699_),
    .ZN(_02594_));
 MUX2_X1 _39427_ (.A(\core.keymem.key_mem[8][6] ),
    .B(_13710_),
    .S(_15064_),
    .Z(_02595_));
 MUX2_X1 _39428_ (.A(\core.keymem.key_mem[8][70] ),
    .B(_13712_),
    .S(_15064_),
    .Z(_02596_));
 NAND2_X1 _39429_ (.A1(\core.keymem.key_mem[8][71] ),
    .A2(_15068_),
    .ZN(_15070_));
 OAI21_X1 _39430_ (.A(_15070_),
    .B1(_15060_),
    .B2(_12658_),
    .ZN(_02597_));
 NAND2_X1 _39431_ (.A1(\core.keymem.key_mem[8][72] ),
    .A2(_15068_),
    .ZN(_15071_));
 OAI21_X1 _39432_ (.A(_15071_),
    .B1(_15060_),
    .B2(_12673_),
    .ZN(_02598_));
 NAND2_X1 _39433_ (.A1(\core.keymem.key_mem[8][73] ),
    .A2(_15068_),
    .ZN(_15072_));
 BUF_X4 _39434_ (.A(_15028_),
    .Z(_15073_));
 OAI21_X1 _39435_ (.A(_15072_),
    .B1(_15073_),
    .B2(_12687_),
    .ZN(_02599_));
 NAND2_X1 _39436_ (.A1(\core.keymem.key_mem[8][74] ),
    .A2(_15068_),
    .ZN(_15074_));
 OAI21_X1 _39437_ (.A(_15074_),
    .B1(_15073_),
    .B2(_13726_),
    .ZN(_02600_));
 NAND2_X1 _39438_ (.A1(\core.keymem.key_mem[8][75] ),
    .A2(_15068_),
    .ZN(_15075_));
 OAI21_X1 _39439_ (.A(_15075_),
    .B1(_15073_),
    .B2(_13732_),
    .ZN(_02601_));
 BUF_X4 _39440_ (.A(_15021_),
    .Z(_15076_));
 MUX2_X1 _39441_ (.A(\core.keymem.key_mem[8][76] ),
    .B(_13740_),
    .S(_15076_),
    .Z(_02602_));
 MUX2_X1 _39442_ (.A(\core.keymem.key_mem[8][77] ),
    .B(_13751_),
    .S(_15076_),
    .Z(_02603_));
 NAND2_X1 _39443_ (.A1(\core.keymem.key_mem[8][78] ),
    .A2(_15068_),
    .ZN(_15077_));
 OAI21_X1 _39444_ (.A(_15077_),
    .B1(_15073_),
    .B2(_12707_),
    .ZN(_02604_));
 MUX2_X1 _39445_ (.A(\core.keymem.key_mem[8][79] ),
    .B(_13758_),
    .S(_15076_),
    .Z(_02605_));
 NAND2_X1 _39446_ (.A1(\core.keymem.key_mem[8][7] ),
    .A2(_15068_),
    .ZN(_15078_));
 OAI21_X1 _39447_ (.A(_15078_),
    .B1(_15073_),
    .B2(_13766_),
    .ZN(_02606_));
 MUX2_X1 _39448_ (.A(\core.keymem.key_mem[8][80] ),
    .B(_13768_),
    .S(_15076_),
    .Z(_02607_));
 NAND2_X1 _39449_ (.A1(\core.keymem.key_mem[8][81] ),
    .A2(_15068_),
    .ZN(_15079_));
 OAI21_X1 _39450_ (.A(_15079_),
    .B1(_15073_),
    .B2(_13774_),
    .ZN(_02608_));
 NAND2_X1 _39451_ (.A1(\core.keymem.key_mem[8][82] ),
    .A2(_15068_),
    .ZN(_15080_));
 OAI21_X1 _39452_ (.A(_15080_),
    .B1(_15073_),
    .B2(_13782_),
    .ZN(_02609_));
 NAND2_X1 _39453_ (.A1(\core.keymem.key_mem[8][83] ),
    .A2(_15028_),
    .ZN(_15081_));
 OAI21_X1 _39454_ (.A(_15081_),
    .B1(_15073_),
    .B2(_13790_),
    .ZN(_02610_));
 NAND2_X1 _39455_ (.A1(\core.keymem.key_mem[8][84] ),
    .A2(_15028_),
    .ZN(_15082_));
 OAI21_X1 _39456_ (.A(_15082_),
    .B1(_15073_),
    .B2(_12724_),
    .ZN(_02611_));
 MUX2_X1 _39457_ (.A(\core.keymem.key_mem[8][85] ),
    .B(_13798_),
    .S(_15076_),
    .Z(_02612_));
 MUX2_X1 _39458_ (.A(\core.keymem.key_mem[8][86] ),
    .B(_12740_),
    .S(_15076_),
    .Z(_02613_));
 MUX2_X1 _39459_ (.A(\core.keymem.key_mem[8][87] ),
    .B(_13804_),
    .S(_15076_),
    .Z(_02614_));
 MUX2_X1 _39460_ (.A(\core.keymem.key_mem[8][88] ),
    .B(_13809_),
    .S(_15076_),
    .Z(_02615_));
 MUX2_X1 _39461_ (.A(\core.keymem.key_mem[8][89] ),
    .B(_13817_),
    .S(_15076_),
    .Z(_02616_));
 MUX2_X1 _39462_ (.A(\core.keymem.key_mem[8][8] ),
    .B(_13854_),
    .S(_15076_),
    .Z(_02617_));
 MUX2_X1 _39463_ (.A(\core.keymem.key_mem[8][90] ),
    .B(_13859_),
    .S(_15022_),
    .Z(_02618_));
 NAND2_X1 _39464_ (.A1(\core.keymem.key_mem[8][91] ),
    .A2(_15028_),
    .ZN(_15083_));
 OAI21_X1 _39465_ (.A(_15083_),
    .B1(_15073_),
    .B2(_13870_),
    .ZN(_02619_));
 NAND2_X1 _39466_ (.A1(\core.keymem.key_mem[8][92] ),
    .A2(_15028_),
    .ZN(_15084_));
 OAI21_X1 _39467_ (.A(_15084_),
    .B1(_15026_),
    .B2(_13880_),
    .ZN(_02620_));
 MUX2_X1 _39468_ (.A(\core.keymem.key_mem[8][93] ),
    .B(_13889_),
    .S(_15022_),
    .Z(_02621_));
 MUX2_X1 _39469_ (.A(\core.keymem.key_mem[8][94] ),
    .B(_13895_),
    .S(_15022_),
    .Z(_02622_));
 MUX2_X1 _39470_ (.A(\core.keymem.key_mem[8][95] ),
    .B(_13902_),
    .S(_15022_),
    .Z(_02623_));
 MUX2_X1 _39471_ (.A(\core.keymem.key_mem[8][96] ),
    .B(_13907_),
    .S(_15022_),
    .Z(_02624_));
 NAND2_X1 _39472_ (.A1(\core.keymem.key_mem[8][97] ),
    .A2(_15028_),
    .ZN(_15085_));
 OAI21_X1 _39473_ (.A(_15085_),
    .B1(_15026_),
    .B2(_12776_),
    .ZN(_02625_));
 NAND2_X1 _39474_ (.A1(\core.keymem.key_mem[8][98] ),
    .A2(_15028_),
    .ZN(_15086_));
 OAI21_X1 _39475_ (.A(_15086_),
    .B1(_15026_),
    .B2(_12787_),
    .ZN(_02626_));
 MUX2_X1 _39476_ (.A(\core.keymem.key_mem[8][99] ),
    .B(_12799_),
    .S(_15022_),
    .Z(_02627_));
 MUX2_X1 _39477_ (.A(\core.keymem.key_mem[8][9] ),
    .B(_13918_),
    .S(_15022_),
    .Z(_02628_));
 NOR2_X4 _39478_ (.A1(_12803_),
    .A2(_14056_),
    .ZN(_15087_));
 BUF_X4 _39479_ (.A(_15087_),
    .Z(_15088_));
 BUF_X4 _39480_ (.A(_15088_),
    .Z(_15089_));
 MUX2_X1 _39481_ (.A(\core.keymem.key_mem[9][0] ),
    .B(_11843_),
    .S(_15089_),
    .Z(_02629_));
 MUX2_X1 _39482_ (.A(\core.keymem.key_mem[9][100] ),
    .B(_11872_),
    .S(_15089_),
    .Z(_02630_));
 MUX2_X1 _39483_ (.A(\core.keymem.key_mem[9][101] ),
    .B(_12812_),
    .S(_15089_),
    .Z(_02631_));
 MUX2_X1 _39484_ (.A(\core.keymem.key_mem[9][102] ),
    .B(_11905_),
    .S(_15089_),
    .Z(_02632_));
 MUX2_X1 _39485_ (.A(\core.keymem.key_mem[9][103] ),
    .B(_11928_),
    .S(_15089_),
    .Z(_02633_));
 OR2_X1 _39486_ (.A1(_12803_),
    .A2(_14056_),
    .ZN(_15090_));
 CLKBUF_X3 _39487_ (.A(_15090_),
    .Z(_15091_));
 BUF_X4 _39488_ (.A(_15091_),
    .Z(_15092_));
 NAND2_X1 _39489_ (.A1(\core.keymem.key_mem[9][104] ),
    .A2(_15092_),
    .ZN(_15093_));
 BUF_X4 _39490_ (.A(_15091_),
    .Z(_15094_));
 BUF_X4 _39491_ (.A(_15094_),
    .Z(_15095_));
 OAI21_X1 _39492_ (.A(_15093_),
    .B1(_15095_),
    .B2(_12821_),
    .ZN(_02634_));
 MUX2_X1 _39493_ (.A(\core.keymem.key_mem[9][105] ),
    .B(_12829_),
    .S(_15089_),
    .Z(_02635_));
 BUF_X4 _39494_ (.A(_15088_),
    .Z(_15096_));
 MUX2_X1 _39495_ (.A(\core.keymem.key_mem[9][106] ),
    .B(_12831_),
    .S(_15096_),
    .Z(_02636_));
 MUX2_X1 _39496_ (.A(\core.keymem.key_mem[9][107] ),
    .B(_11966_),
    .S(_15096_),
    .Z(_02637_));
 MUX2_X1 _39497_ (.A(\core.keymem.key_mem[9][108] ),
    .B(_11980_),
    .S(_15096_),
    .Z(_02638_));
 MUX2_X1 _39498_ (.A(\core.keymem.key_mem[9][109] ),
    .B(_12841_),
    .S(_15096_),
    .Z(_02639_));
 NAND2_X1 _39499_ (.A1(\core.keymem.key_mem[9][10] ),
    .A2(_15092_),
    .ZN(_15097_));
 OAI21_X1 _39500_ (.A(_15097_),
    .B1(_15095_),
    .B2(_12857_),
    .ZN(_02640_));
 MUX2_X1 _39501_ (.A(\core.keymem.key_mem[9][110] ),
    .B(_12003_),
    .S(_15096_),
    .Z(_02641_));
 MUX2_X1 _39502_ (.A(\core.keymem.key_mem[9][111] ),
    .B(_12016_),
    .S(_15096_),
    .Z(_02642_));
 MUX2_X1 _39503_ (.A(\core.keymem.key_mem[9][112] ),
    .B(_12030_),
    .S(_15096_),
    .Z(_02643_));
 MUX2_X1 _39504_ (.A(\core.keymem.key_mem[9][113] ),
    .B(_12867_),
    .S(_15096_),
    .Z(_02644_));
 MUX2_X1 _39505_ (.A(\core.keymem.key_mem[9][114] ),
    .B(_12048_),
    .S(_15096_),
    .Z(_02645_));
 MUX2_X1 _39506_ (.A(\core.keymem.key_mem[9][115] ),
    .B(_12058_),
    .S(_15096_),
    .Z(_02646_));
 BUF_X4 _39507_ (.A(_15088_),
    .Z(_15098_));
 MUX2_X1 _39508_ (.A(\core.keymem.key_mem[9][116] ),
    .B(_12076_),
    .S(_15098_),
    .Z(_02647_));
 MUX2_X1 _39509_ (.A(\core.keymem.key_mem[9][117] ),
    .B(_12876_),
    .S(_15098_),
    .Z(_02648_));
 MUX2_X1 _39510_ (.A(\core.keymem.key_mem[9][118] ),
    .B(_12881_),
    .S(_15098_),
    .Z(_02649_));
 MUX2_X1 _39511_ (.A(\core.keymem.key_mem[9][119] ),
    .B(_12095_),
    .S(_15098_),
    .Z(_02650_));
 NAND2_X1 _39512_ (.A1(\core.keymem.key_mem[9][11] ),
    .A2(_15092_),
    .ZN(_15099_));
 OAI21_X1 _39513_ (.A(_15099_),
    .B1(_15095_),
    .B2(_12894_),
    .ZN(_02651_));
 MUX2_X1 _39514_ (.A(\core.keymem.key_mem[9][120] ),
    .B(_12123_),
    .S(_15098_),
    .Z(_02652_));
 MUX2_X1 _39515_ (.A(\core.keymem.key_mem[9][121] ),
    .B(_12159_),
    .S(_15098_),
    .Z(_02653_));
 MUX2_X1 _39516_ (.A(\core.keymem.key_mem[9][122] ),
    .B(_12902_),
    .S(_15098_),
    .Z(_02654_));
 NAND2_X1 _39517_ (.A1(\core.keymem.key_mem[9][123] ),
    .A2(_15092_),
    .ZN(_15100_));
 OAI21_X1 _39518_ (.A(_15100_),
    .B1(_15095_),
    .B2(_12181_),
    .ZN(_02655_));
 NAND2_X1 _39519_ (.A1(\core.keymem.key_mem[9][124] ),
    .A2(_15092_),
    .ZN(_15101_));
 OAI21_X1 _39520_ (.A(_15101_),
    .B1(_15095_),
    .B2(_12925_),
    .ZN(_02656_));
 MUX2_X1 _39521_ (.A(\core.keymem.key_mem[9][125] ),
    .B(_12931_),
    .S(_15098_),
    .Z(_02657_));
 NAND2_X1 _39522_ (.A1(\core.keymem.key_mem[9][126] ),
    .A2(_15092_),
    .ZN(_15102_));
 OAI21_X1 _39523_ (.A(_15102_),
    .B1(_15095_),
    .B2(_12206_),
    .ZN(_02658_));
 MUX2_X1 _39524_ (.A(\core.keymem.key_mem[9][127] ),
    .B(_12944_),
    .S(_15098_),
    .Z(_02659_));
 MUX2_X1 _39525_ (.A(\core.keymem.key_mem[9][12] ),
    .B(_12957_),
    .S(_15098_),
    .Z(_02660_));
 BUF_X4 _39526_ (.A(_15087_),
    .Z(_15103_));
 MUX2_X1 _39527_ (.A(\core.keymem.key_mem[9][13] ),
    .B(_12973_),
    .S(_15103_),
    .Z(_02661_));
 NOR2_X1 _39528_ (.A1(\core.keymem.key_mem[9][14] ),
    .A2(_15089_),
    .ZN(_15104_));
 AOI21_X1 _39529_ (.A(_15104_),
    .B1(_15089_),
    .B2(_13006_),
    .ZN(_02662_));
 MUX2_X1 _39530_ (.A(\core.keymem.key_mem[9][15] ),
    .B(_13016_),
    .S(_15103_),
    .Z(_02663_));
 MUX2_X1 _39531_ (.A(\core.keymem.key_mem[9][16] ),
    .B(_13028_),
    .S(_15103_),
    .Z(_02664_));
 NAND2_X1 _39532_ (.A1(\core.keymem.key_mem[9][17] ),
    .A2(_15092_),
    .ZN(_15105_));
 OAI21_X1 _39533_ (.A(_15105_),
    .B1(_15095_),
    .B2(_13041_),
    .ZN(_02665_));
 MUX2_X1 _39534_ (.A(\core.keymem.key_mem[9][18] ),
    .B(_13093_),
    .S(_15103_),
    .Z(_02666_));
 BUF_X4 _39535_ (.A(_15091_),
    .Z(_15106_));
 NAND2_X1 _39536_ (.A1(\core.keymem.key_mem[9][19] ),
    .A2(_15106_),
    .ZN(_15107_));
 OAI21_X1 _39537_ (.A(_15107_),
    .B1(_15095_),
    .B2(_13108_),
    .ZN(_02667_));
 MUX2_X1 _39538_ (.A(\core.keymem.key_mem[9][1] ),
    .B(_13133_),
    .S(_15103_),
    .Z(_02668_));
 MUX2_X1 _39539_ (.A(\core.keymem.key_mem[9][20] ),
    .B(_13145_),
    .S(_15103_),
    .Z(_02669_));
 MUX2_X1 _39540_ (.A(\core.keymem.key_mem[9][21] ),
    .B(_13154_),
    .S(_15103_),
    .Z(_02670_));
 NOR2_X1 _39541_ (.A1(\core.keymem.key_mem[9][22] ),
    .A2(_15089_),
    .ZN(_15108_));
 AOI21_X1 _39542_ (.A(_15108_),
    .B1(_15089_),
    .B2(_13190_),
    .ZN(_02671_));
 MUX2_X1 _39543_ (.A(\core.keymem.key_mem[9][23] ),
    .B(_13195_),
    .S(_15103_),
    .Z(_02672_));
 NAND2_X1 _39544_ (.A1(\core.keymem.key_mem[9][24] ),
    .A2(_15106_),
    .ZN(_15109_));
 OAI21_X1 _39545_ (.A(_15109_),
    .B1(_15095_),
    .B2(_13211_),
    .ZN(_02673_));
 MUX2_X1 _39546_ (.A(\core.keymem.key_mem[9][25] ),
    .B(_13232_),
    .S(_15103_),
    .Z(_02674_));
 MUX2_X1 _39547_ (.A(\core.keymem.key_mem[9][26] ),
    .B(_13240_),
    .S(_15103_),
    .Z(_02675_));
 BUF_X4 _39548_ (.A(_15087_),
    .Z(_15110_));
 MUX2_X1 _39549_ (.A(\core.keymem.key_mem[9][27] ),
    .B(_13283_),
    .S(_15110_),
    .Z(_02676_));
 MUX2_X1 _39550_ (.A(\core.keymem.key_mem[9][28] ),
    .B(_13324_),
    .S(_15110_),
    .Z(_02677_));
 MUX2_X1 _39551_ (.A(\core.keymem.key_mem[9][29] ),
    .B(_13328_),
    .S(_15110_),
    .Z(_02678_));
 NAND2_X1 _39552_ (.A1(\core.keymem.key_mem[9][2] ),
    .A2(_15106_),
    .ZN(_15111_));
 OAI21_X1 _39553_ (.A(_15111_),
    .B1(_15095_),
    .B2(_13334_),
    .ZN(_02679_));
 MUX2_X1 _39554_ (.A(\core.keymem.key_mem[9][30] ),
    .B(_13378_),
    .S(_15110_),
    .Z(_02680_));
 MUX2_X1 _39555_ (.A(\core.keymem.key_mem[9][31] ),
    .B(_13394_),
    .S(_15110_),
    .Z(_02681_));
 MUX2_X1 _39556_ (.A(\core.keymem.key_mem[9][32] ),
    .B(_12354_),
    .S(_15110_),
    .Z(_02682_));
 MUX2_X1 _39557_ (.A(\core.keymem.key_mem[9][33] ),
    .B(_13401_),
    .S(_15110_),
    .Z(_02683_));
 MUX2_X1 _39558_ (.A(\core.keymem.key_mem[9][34] ),
    .B(_12375_),
    .S(_15110_),
    .Z(_02684_));
 MUX2_X1 _39559_ (.A(\core.keymem.key_mem[9][35] ),
    .B(_13404_),
    .S(_15110_),
    .Z(_02685_));
 NAND2_X1 _39560_ (.A1(\core.keymem.key_mem[9][36] ),
    .A2(_15106_),
    .ZN(_15112_));
 BUF_X4 _39561_ (.A(_15094_),
    .Z(_15113_));
 OAI21_X1 _39562_ (.A(_15112_),
    .B1(_15113_),
    .B2(_12422_),
    .ZN(_02686_));
 NAND2_X1 _39563_ (.A1(\core.keymem.key_mem[9][37] ),
    .A2(_15106_),
    .ZN(_15114_));
 OAI21_X1 _39564_ (.A(_15114_),
    .B1(_15113_),
    .B2(_12438_),
    .ZN(_02687_));
 MUX2_X1 _39565_ (.A(\core.keymem.key_mem[9][38] ),
    .B(_13409_),
    .S(_15110_),
    .Z(_02688_));
 NAND2_X1 _39566_ (.A1(\core.keymem.key_mem[9][39] ),
    .A2(_15106_),
    .ZN(_15115_));
 OAI21_X1 _39567_ (.A(_15115_),
    .B1(_15113_),
    .B2(_13434_),
    .ZN(_02689_));
 NAND2_X1 _39568_ (.A1(\core.keymem.key_mem[9][3] ),
    .A2(_15106_),
    .ZN(_15116_));
 OAI21_X1 _39569_ (.A(_15116_),
    .B1(_15113_),
    .B2(_13447_),
    .ZN(_02690_));
 NAND2_X1 _39570_ (.A1(\core.keymem.key_mem[9][40] ),
    .A2(_15106_),
    .ZN(_15117_));
 OAI21_X1 _39571_ (.A(_15117_),
    .B1(_15113_),
    .B2(_13456_),
    .ZN(_02691_));
 BUF_X4 _39572_ (.A(_15087_),
    .Z(_15118_));
 MUX2_X1 _39573_ (.A(\core.keymem.key_mem[9][41] ),
    .B(_13466_),
    .S(_15118_),
    .Z(_02692_));
 MUX2_X1 _39574_ (.A(\core.keymem.key_mem[9][42] ),
    .B(_13489_),
    .S(_15118_),
    .Z(_02693_));
 NAND2_X1 _39575_ (.A1(\core.keymem.key_mem[9][43] ),
    .A2(_15106_),
    .ZN(_15119_));
 OAI21_X1 _39576_ (.A(_15119_),
    .B1(_15113_),
    .B2(_13495_),
    .ZN(_02694_));
 MUX2_X1 _39577_ (.A(\core.keymem.key_mem[9][44] ),
    .B(_12505_),
    .S(_15118_),
    .Z(_02695_));
 NAND2_X1 _39578_ (.A1(\core.keymem.key_mem[9][45] ),
    .A2(_15106_),
    .ZN(_15120_));
 OAI21_X1 _39579_ (.A(_15120_),
    .B1(_15113_),
    .B2(_13509_),
    .ZN(_02696_));
 BUF_X4 _39580_ (.A(_15091_),
    .Z(_15121_));
 NAND2_X1 _39581_ (.A1(\core.keymem.key_mem[9][46] ),
    .A2(_15121_),
    .ZN(_15122_));
 OAI21_X1 _39582_ (.A(_15122_),
    .B1(_15113_),
    .B2(_13516_),
    .ZN(_02697_));
 NAND2_X1 _39583_ (.A1(\core.keymem.key_mem[9][47] ),
    .A2(_15121_),
    .ZN(_15123_));
 OAI21_X1 _39584_ (.A(_15123_),
    .B1(_15113_),
    .B2(_12519_),
    .ZN(_02698_));
 NAND2_X1 _39585_ (.A1(\core.keymem.key_mem[9][48] ),
    .A2(_15121_),
    .ZN(_15124_));
 OAI21_X1 _39586_ (.A(_15124_),
    .B1(_15113_),
    .B2(_12531_),
    .ZN(_02699_));
 NAND2_X1 _39587_ (.A1(\core.keymem.key_mem[9][49] ),
    .A2(_15121_),
    .ZN(_15125_));
 BUF_X4 _39588_ (.A(_15094_),
    .Z(_15126_));
 OAI21_X1 _39589_ (.A(_15125_),
    .B1(_15126_),
    .B2(_13528_),
    .ZN(_02700_));
 MUX2_X1 _39590_ (.A(\core.keymem.key_mem[9][4] ),
    .B(_13537_),
    .S(_15118_),
    .Z(_02701_));
 MUX2_X1 _39591_ (.A(\core.keymem.key_mem[9][50] ),
    .B(_13556_),
    .S(_15118_),
    .Z(_02702_));
 MUX2_X1 _39592_ (.A(\core.keymem.key_mem[9][51] ),
    .B(_13563_),
    .S(_15118_),
    .Z(_02703_));
 NAND2_X1 _39593_ (.A1(\core.keymem.key_mem[9][52] ),
    .A2(_15121_),
    .ZN(_15127_));
 OAI21_X1 _39594_ (.A(_15127_),
    .B1(_15126_),
    .B2(_12567_),
    .ZN(_02704_));
 NAND2_X1 _39595_ (.A1(\core.keymem.key_mem[9][53] ),
    .A2(_15121_),
    .ZN(_15128_));
 OAI21_X1 _39596_ (.A(_15128_),
    .B1(_15126_),
    .B2(_12583_),
    .ZN(_02705_));
 NAND2_X1 _39597_ (.A1(\core.keymem.key_mem[9][54] ),
    .A2(_15121_),
    .ZN(_15129_));
 OAI21_X1 _39598_ (.A(_15129_),
    .B1(_15126_),
    .B2(_13574_),
    .ZN(_02706_));
 MUX2_X1 _39599_ (.A(\core.keymem.key_mem[9][55] ),
    .B(_13580_),
    .S(_15118_),
    .Z(_02707_));
 MUX2_X1 _39600_ (.A(\core.keymem.key_mem[9][56] ),
    .B(_13588_),
    .S(_15118_),
    .Z(_02708_));
 MUX2_X1 _39601_ (.A(\core.keymem.key_mem[9][57] ),
    .B(_13603_),
    .S(_15118_),
    .Z(_02709_));
 MUX2_X1 _39602_ (.A(\core.keymem.key_mem[9][58] ),
    .B(_13610_),
    .S(_15118_),
    .Z(_02710_));
 BUF_X4 _39603_ (.A(_15087_),
    .Z(_15130_));
 MUX2_X1 _39604_ (.A(\core.keymem.key_mem[9][59] ),
    .B(_13615_),
    .S(_15130_),
    .Z(_02711_));
 MUX2_X1 _39605_ (.A(\core.keymem.key_mem[9][5] ),
    .B(_12605_),
    .S(_15130_),
    .Z(_02712_));
 MUX2_X1 _39606_ (.A(\core.keymem.key_mem[9][60] ),
    .B(_13621_),
    .S(_15130_),
    .Z(_02713_));
 MUX2_X1 _39607_ (.A(\core.keymem.key_mem[9][61] ),
    .B(_13631_),
    .S(_15130_),
    .Z(_02714_));
 MUX2_X1 _39608_ (.A(\core.keymem.key_mem[9][62] ),
    .B(_13636_),
    .S(_15130_),
    .Z(_02715_));
 MUX2_X1 _39609_ (.A(\core.keymem.key_mem[9][63] ),
    .B(_13658_),
    .S(_15130_),
    .Z(_02716_));
 MUX2_X1 _39610_ (.A(\core.keymem.key_mem[9][64] ),
    .B(_12621_),
    .S(_15130_),
    .Z(_02717_));
 NAND2_X1 _39611_ (.A1(\core.keymem.key_mem[9][65] ),
    .A2(_15121_),
    .ZN(_15131_));
 OAI21_X1 _39612_ (.A(_15131_),
    .B1(_15126_),
    .B2(_13672_),
    .ZN(_02718_));
 MUX2_X1 _39613_ (.A(\core.keymem.key_mem[9][66] ),
    .B(_13680_),
    .S(_15130_),
    .Z(_02719_));
 NAND2_X1 _39614_ (.A1(\core.keymem.key_mem[9][67] ),
    .A2(_15121_),
    .ZN(_15132_));
 OAI21_X1 _39615_ (.A(_15132_),
    .B1(_15126_),
    .B2(_13689_),
    .ZN(_02720_));
 NAND2_X1 _39616_ (.A1(\core.keymem.key_mem[9][68] ),
    .A2(_15121_),
    .ZN(_15133_));
 OAI21_X1 _39617_ (.A(_15133_),
    .B1(_15126_),
    .B2(_12634_),
    .ZN(_02721_));
 BUF_X4 _39618_ (.A(_15091_),
    .Z(_15134_));
 NAND2_X1 _39619_ (.A1(\core.keymem.key_mem[9][69] ),
    .A2(_15134_),
    .ZN(_15135_));
 OAI21_X1 _39620_ (.A(_15135_),
    .B1(_15126_),
    .B2(_13699_),
    .ZN(_02722_));
 MUX2_X1 _39621_ (.A(\core.keymem.key_mem[9][6] ),
    .B(_13710_),
    .S(_15130_),
    .Z(_02723_));
 MUX2_X1 _39622_ (.A(\core.keymem.key_mem[9][70] ),
    .B(_13712_),
    .S(_15130_),
    .Z(_02724_));
 NAND2_X1 _39623_ (.A1(\core.keymem.key_mem[9][71] ),
    .A2(_15134_),
    .ZN(_15136_));
 OAI21_X1 _39624_ (.A(_15136_),
    .B1(_15126_),
    .B2(_12658_),
    .ZN(_02725_));
 NAND2_X1 _39625_ (.A1(\core.keymem.key_mem[9][72] ),
    .A2(_15134_),
    .ZN(_15137_));
 OAI21_X1 _39626_ (.A(_15137_),
    .B1(_15126_),
    .B2(_12673_),
    .ZN(_02726_));
 NAND2_X1 _39627_ (.A1(\core.keymem.key_mem[9][73] ),
    .A2(_15134_),
    .ZN(_15138_));
 BUF_X4 _39628_ (.A(_15094_),
    .Z(_15139_));
 OAI21_X1 _39629_ (.A(_15138_),
    .B1(_15139_),
    .B2(_12687_),
    .ZN(_02727_));
 NAND2_X1 _39630_ (.A1(\core.keymem.key_mem[9][74] ),
    .A2(_15134_),
    .ZN(_15140_));
 OAI21_X1 _39631_ (.A(_15140_),
    .B1(_15139_),
    .B2(_13725_),
    .ZN(_02728_));
 NAND2_X1 _39632_ (.A1(\core.keymem.key_mem[9][75] ),
    .A2(_15134_),
    .ZN(_15141_));
 OAI21_X1 _39633_ (.A(_15141_),
    .B1(_15139_),
    .B2(_13732_),
    .ZN(_02729_));
 BUF_X4 _39634_ (.A(_15087_),
    .Z(_15142_));
 MUX2_X1 _39635_ (.A(\core.keymem.key_mem[9][76] ),
    .B(_13740_),
    .S(_15142_),
    .Z(_02730_));
 MUX2_X1 _39636_ (.A(\core.keymem.key_mem[9][77] ),
    .B(_13750_),
    .S(_15142_),
    .Z(_02731_));
 NAND2_X1 _39637_ (.A1(\core.keymem.key_mem[9][78] ),
    .A2(_15134_),
    .ZN(_15143_));
 OAI21_X1 _39638_ (.A(_15143_),
    .B1(_15139_),
    .B2(_12707_),
    .ZN(_02732_));
 MUX2_X1 _39639_ (.A(\core.keymem.key_mem[9][79] ),
    .B(_13757_),
    .S(_15142_),
    .Z(_02733_));
 NAND2_X1 _39640_ (.A1(\core.keymem.key_mem[9][7] ),
    .A2(_15134_),
    .ZN(_15144_));
 OAI21_X1 _39641_ (.A(_15144_),
    .B1(_15139_),
    .B2(_13766_),
    .ZN(_02734_));
 MUX2_X1 _39642_ (.A(\core.keymem.key_mem[9][80] ),
    .B(_13768_),
    .S(_15142_),
    .Z(_02735_));
 NAND2_X1 _39643_ (.A1(\core.keymem.key_mem[9][81] ),
    .A2(_15134_),
    .ZN(_15145_));
 OAI21_X1 _39644_ (.A(_15145_),
    .B1(_15139_),
    .B2(_13774_),
    .ZN(_02736_));
 NAND2_X1 _39645_ (.A1(\core.keymem.key_mem[9][82] ),
    .A2(_15134_),
    .ZN(_15146_));
 OAI21_X1 _39646_ (.A(_15146_),
    .B1(_15139_),
    .B2(_13782_),
    .ZN(_02737_));
 NAND2_X1 _39647_ (.A1(\core.keymem.key_mem[9][83] ),
    .A2(_15094_),
    .ZN(_15147_));
 OAI21_X1 _39648_ (.A(_15147_),
    .B1(_15139_),
    .B2(_13790_),
    .ZN(_02738_));
 NAND2_X1 _39649_ (.A1(\core.keymem.key_mem[9][84] ),
    .A2(_15094_),
    .ZN(_15148_));
 OAI21_X1 _39650_ (.A(_15148_),
    .B1(_15139_),
    .B2(_12724_),
    .ZN(_02739_));
 MUX2_X1 _39651_ (.A(\core.keymem.key_mem[9][85] ),
    .B(_13797_),
    .S(_15142_),
    .Z(_02740_));
 MUX2_X1 _39652_ (.A(\core.keymem.key_mem[9][86] ),
    .B(_12740_),
    .S(_15142_),
    .Z(_02741_));
 MUX2_X1 _39653_ (.A(\core.keymem.key_mem[9][87] ),
    .B(_13803_),
    .S(_15142_),
    .Z(_02742_));
 MUX2_X1 _39654_ (.A(\core.keymem.key_mem[9][88] ),
    .B(_13809_),
    .S(_15142_),
    .Z(_02743_));
 MUX2_X1 _39655_ (.A(\core.keymem.key_mem[9][89] ),
    .B(_13817_),
    .S(_15142_),
    .Z(_02744_));
 MUX2_X1 _39656_ (.A(\core.keymem.key_mem[9][8] ),
    .B(_13853_),
    .S(_15142_),
    .Z(_02745_));
 MUX2_X1 _39657_ (.A(\core.keymem.key_mem[9][90] ),
    .B(_13859_),
    .S(_15088_),
    .Z(_02746_));
 NAND2_X1 _39658_ (.A1(\core.keymem.key_mem[9][91] ),
    .A2(_15094_),
    .ZN(_15149_));
 OAI21_X1 _39659_ (.A(_15149_),
    .B1(_15139_),
    .B2(_13869_),
    .ZN(_02747_));
 NAND2_X1 _39660_ (.A1(\core.keymem.key_mem[9][92] ),
    .A2(_15094_),
    .ZN(_15150_));
 OAI21_X1 _39661_ (.A(_15150_),
    .B1(_15092_),
    .B2(_13879_),
    .ZN(_02748_));
 MUX2_X1 _39662_ (.A(\core.keymem.key_mem[9][93] ),
    .B(_13888_),
    .S(_15088_),
    .Z(_02749_));
 MUX2_X1 _39663_ (.A(\core.keymem.key_mem[9][94] ),
    .B(_13895_),
    .S(_15088_),
    .Z(_02750_));
 MUX2_X1 _39664_ (.A(\core.keymem.key_mem[9][95] ),
    .B(_13902_),
    .S(_15088_),
    .Z(_02751_));
 MUX2_X1 _39665_ (.A(\core.keymem.key_mem[9][96] ),
    .B(_13906_),
    .S(_15088_),
    .Z(_02752_));
 NAND2_X1 _39666_ (.A1(\core.keymem.key_mem[9][97] ),
    .A2(_15094_),
    .ZN(_15151_));
 OAI21_X1 _39667_ (.A(_15151_),
    .B1(_15092_),
    .B2(_12776_),
    .ZN(_02753_));
 NAND2_X1 _39668_ (.A1(\core.keymem.key_mem[9][98] ),
    .A2(_15094_),
    .ZN(_15152_));
 OAI21_X1 _39669_ (.A(_15152_),
    .B1(_15092_),
    .B2(_12787_),
    .ZN(_02754_));
 MUX2_X1 _39670_ (.A(\core.keymem.key_mem[9][99] ),
    .B(_12799_),
    .S(_15088_),
    .Z(_02755_));
 MUX2_X1 _39671_ (.A(\core.keymem.key_mem[9][9] ),
    .B(_13918_),
    .S(_15088_),
    .Z(_02756_));
 CLKBUF_X3 _39672_ (.A(_22091_),
    .Z(_15153_));
 NOR3_X4 _39673_ (.A1(_11804_),
    .A2(_15153_),
    .A3(_12946_),
    .ZN(_15154_));
 BUF_X4 _39674_ (.A(_15154_),
    .Z(_15155_));
 BUF_X4 _39675_ (.A(_15155_),
    .Z(_15156_));
 NOR2_X1 _39676_ (.A1(\core.keymem.prev_key0_reg[0] ),
    .A2(_15156_),
    .ZN(_15157_));
 NOR2_X1 _39677_ (.A1(_00327_),
    .A2(_12834_),
    .ZN(_15158_));
 BUF_X4 _39678_ (.A(_13011_),
    .Z(_15159_));
 BUF_X4 _39679_ (.A(_15159_),
    .Z(_15160_));
 AOI21_X1 _39680_ (.A(_15158_),
    .B1(_15160_),
    .B2(_06858_),
    .ZN(_15161_));
 BUF_X4 _39681_ (.A(_15154_),
    .Z(_15162_));
 BUF_X4 _39682_ (.A(_15162_),
    .Z(_15163_));
 AOI21_X1 _39683_ (.A(_15157_),
    .B1(_15161_),
    .B2(_15163_),
    .ZN(_02757_));
 BUF_X4 _39684_ (.A(_13136_),
    .Z(_15164_));
 OAI22_X1 _39685_ (.A1(_00127_),
    .A2(_14201_),
    .B1(_15164_),
    .B2(_00128_),
    .ZN(_15165_));
 BUF_X4 _39686_ (.A(_15155_),
    .Z(_15166_));
 MUX2_X1 _39687_ (.A(\core.keymem.prev_key0_reg[100] ),
    .B(_15165_),
    .S(_15166_),
    .Z(_02758_));
 OAI22_X1 _39688_ (.A1(_00129_),
    .A2(_14201_),
    .B1(_15164_),
    .B2(_00377_),
    .ZN(_15167_));
 MUX2_X1 _39689_ (.A(\core.keymem.prev_key0_reg[101] ),
    .B(_15167_),
    .S(_15166_),
    .Z(_02759_));
 OAI22_X1 _39690_ (.A1(_00130_),
    .A2(_14201_),
    .B1(_15164_),
    .B2(_00379_),
    .ZN(_15168_));
 MUX2_X1 _39691_ (.A(_11894_),
    .B(_15168_),
    .S(_15166_),
    .Z(_02760_));
 BUF_X4 _39692_ (.A(_13136_),
    .Z(_15169_));
 OAI21_X1 _39693_ (.A(_11915_),
    .B1(_15169_),
    .B2(_00132_),
    .ZN(_15170_));
 MUX2_X1 _39694_ (.A(_11918_),
    .B(_15170_),
    .S(_15166_),
    .Z(_02761_));
 NOR2_X1 _39695_ (.A1(_12667_),
    .A2(_15156_),
    .ZN(_15171_));
 NOR2_X1 _39696_ (.A1(_00133_),
    .A2(_13720_),
    .ZN(_15172_));
 AOI21_X1 _39697_ (.A(_15172_),
    .B1(_15160_),
    .B2(\core.keymem.prev_key1_reg[104] ),
    .ZN(_15173_));
 AOI21_X1 _39698_ (.A(_15171_),
    .B1(_15173_),
    .B2(_15163_),
    .ZN(_02762_));
 NOR2_X1 _39699_ (.A1(\core.keymem.prev_key0_reg[105] ),
    .A2(_15156_),
    .ZN(_15174_));
 NOR2_X1 _39700_ (.A1(_00134_),
    .A2(_14447_),
    .ZN(_15175_));
 AOI21_X1 _39701_ (.A(_15175_),
    .B1(_15160_),
    .B2(\core.keymem.prev_key1_reg[105] ),
    .ZN(_15176_));
 AOI21_X1 _39702_ (.A(_15174_),
    .B1(_15176_),
    .B2(_15163_),
    .ZN(_02763_));
 OAI21_X1 _39703_ (.A(_11935_),
    .B1(_15169_),
    .B2(_00136_),
    .ZN(_15177_));
 MUX2_X1 _39704_ (.A(_11937_),
    .B(_15177_),
    .S(_15166_),
    .Z(_02764_));
 BUF_X4 _39705_ (.A(_13136_),
    .Z(_15178_));
 OAI22_X2 _39706_ (.A1(_00137_),
    .A2(_14201_),
    .B1(_15178_),
    .B2(_00138_),
    .ZN(_15179_));
 MUX2_X1 _39707_ (.A(\core.keymem.prev_key0_reg[107] ),
    .B(_15179_),
    .S(_15166_),
    .Z(_02765_));
 OAI21_X1 _39708_ (.A(_11977_),
    .B1(_15169_),
    .B2(_00140_),
    .ZN(_15180_));
 BUF_X4 _39709_ (.A(_15155_),
    .Z(_15181_));
 MUX2_X1 _39710_ (.A(_11969_),
    .B(_15180_),
    .S(_15181_),
    .Z(_02766_));
 BUF_X4 _39711_ (.A(_15155_),
    .Z(_15182_));
 NOR2_X1 _39712_ (.A1(_12835_),
    .A2(_15182_),
    .ZN(_15183_));
 NOR2_X1 _39713_ (.A1(_00141_),
    .A2(_13875_),
    .ZN(_15184_));
 AOI21_X1 _39714_ (.A(_15184_),
    .B1(_15160_),
    .B2(\core.keymem.prev_key1_reg[109] ),
    .ZN(_15185_));
 AOI21_X1 _39715_ (.A(_15183_),
    .B1(_15185_),
    .B2(_15163_),
    .ZN(_02767_));
 OAI22_X1 _39716_ (.A1(_11983_),
    .A2(_14201_),
    .B1(_15178_),
    .B2(_07272_),
    .ZN(_15186_));
 MUX2_X1 _39717_ (.A(\core.keymem.prev_key0_reg[10] ),
    .B(_15186_),
    .S(_15181_),
    .Z(_02768_));
 NOR2_X1 _39718_ (.A1(_11992_),
    .A2(_15182_),
    .ZN(_15187_));
 NOR2_X1 _39719_ (.A1(_00142_),
    .A2(_12834_),
    .ZN(_15188_));
 AOI21_X1 _39720_ (.A(_15188_),
    .B1(_15160_),
    .B2(_11999_),
    .ZN(_15189_));
 AOI21_X1 _39721_ (.A(_15187_),
    .B1(_15189_),
    .B2(_15163_),
    .ZN(_02769_));
 OAI21_X1 _39722_ (.A(_12011_),
    .B1(_15169_),
    .B2(_00144_),
    .ZN(_15190_));
 MUX2_X1 _39723_ (.A(\core.keymem.prev_key0_reg[111] ),
    .B(_15190_),
    .S(_15181_),
    .Z(_02770_));
 NOR2_X1 _39724_ (.A1(\core.keymem.prev_key0_reg[112] ),
    .A2(_15182_),
    .ZN(_15191_));
 AOI21_X1 _39725_ (.A(_12024_),
    .B1(_15160_),
    .B2(_12025_),
    .ZN(_15192_));
 AOI21_X1 _39726_ (.A(_15191_),
    .B1(_15192_),
    .B2(_15163_),
    .ZN(_02771_));
 NOR2_X1 _39727_ (.A1(\core.keymem.prev_key0_reg[113] ),
    .A2(_15182_),
    .ZN(_15193_));
 NOR2_X1 _39728_ (.A1(_00146_),
    .A2(_13720_),
    .ZN(_15194_));
 AOI21_X1 _39729_ (.A(_15194_),
    .B1(_15160_),
    .B2(\core.keymem.prev_key1_reg[113] ),
    .ZN(_15195_));
 AOI21_X1 _39730_ (.A(_15193_),
    .B1(_15195_),
    .B2(_15163_),
    .ZN(_02772_));
 OAI22_X1 _39731_ (.A1(_00147_),
    .A2(_14201_),
    .B1(_15178_),
    .B2(_00148_),
    .ZN(_15196_));
 MUX2_X1 _39732_ (.A(_12037_),
    .B(_15196_),
    .S(_15181_),
    .Z(_02773_));
 OAI21_X1 _39733_ (.A(_12055_),
    .B1(_15169_),
    .B2(_00150_),
    .ZN(_15197_));
 MUX2_X1 _39734_ (.A(\core.keymem.prev_key0_reg[115] ),
    .B(_15197_),
    .S(_15181_),
    .Z(_02774_));
 OAI21_X1 _39735_ (.A(_12072_),
    .B1(_15169_),
    .B2(_00152_),
    .ZN(_15198_));
 MUX2_X1 _39736_ (.A(_12061_),
    .B(_15198_),
    .S(_15181_),
    .Z(_02775_));
 NOR2_X1 _39737_ (.A1(\core.keymem.prev_key0_reg[117] ),
    .A2(_15182_),
    .ZN(_15199_));
 NOR2_X1 _39738_ (.A1(_00153_),
    .A2(_13720_),
    .ZN(_15200_));
 AOI21_X1 _39739_ (.A(_15200_),
    .B1(_15160_),
    .B2(\core.keymem.prev_key1_reg[117] ),
    .ZN(_15201_));
 AOI21_X1 _39740_ (.A(_15199_),
    .B1(_15201_),
    .B2(_15163_),
    .ZN(_02776_));
 NOR2_X1 _39741_ (.A1(\core.keymem.prev_key0_reg[118] ),
    .A2(_15182_),
    .ZN(_15202_));
 NOR2_X2 _39742_ (.A1(_00154_),
    .A2(_14447_),
    .ZN(_15203_));
 AOI21_X1 _39743_ (.A(_15203_),
    .B1(_15160_),
    .B2(\core.keymem.prev_key1_reg[118] ),
    .ZN(_15204_));
 AOI21_X1 _39744_ (.A(_15202_),
    .B1(_15204_),
    .B2(_15163_),
    .ZN(_02777_));
 OAI21_X1 _39745_ (.A(_12087_),
    .B1(_15169_),
    .B2(_00156_),
    .ZN(_15205_));
 MUX2_X1 _39746_ (.A(_12089_),
    .B(_15205_),
    .S(_15181_),
    .Z(_02778_));
 NOR2_X1 _39747_ (.A1(\core.keymem.prev_key0_reg[11] ),
    .A2(_15182_),
    .ZN(_15206_));
 AOI21_X1 _39748_ (.A(_14253_),
    .B1(_15160_),
    .B2(_07382_),
    .ZN(_15207_));
 AOI21_X1 _39749_ (.A(_15206_),
    .B1(_15207_),
    .B2(_15163_),
    .ZN(_02779_));
 OAI22_X1 _39750_ (.A1(_00157_),
    .A2(_14201_),
    .B1(_15178_),
    .B2(_00018_),
    .ZN(_15208_));
 MUX2_X1 _39751_ (.A(\core.keymem.prev_key0_reg[120] ),
    .B(_15208_),
    .S(_15181_),
    .Z(_02780_));
 BUF_X4 _39752_ (.A(_12871_),
    .Z(_15209_));
 OAI22_X1 _39753_ (.A1(_00159_),
    .A2(_15209_),
    .B1(_15178_),
    .B2(_00021_),
    .ZN(_15210_));
 MUX2_X1 _39754_ (.A(_12126_),
    .B(_15210_),
    .S(_15181_),
    .Z(_02781_));
 OAI21_X1 _39755_ (.A(_12897_),
    .B1(_15169_),
    .B2(_00024_),
    .ZN(_15211_));
 MUX2_X1 _39756_ (.A(\core.keymem.prev_key0_reg[122] ),
    .B(_15211_),
    .S(_15181_),
    .Z(_02782_));
 OAI22_X1 _39757_ (.A1(_00163_),
    .A2(_15209_),
    .B1(_15178_),
    .B2(_00027_),
    .ZN(_15212_));
 BUF_X4 _39758_ (.A(_15154_),
    .Z(_15213_));
 MUX2_X1 _39759_ (.A(_12173_),
    .B(_15212_),
    .S(_15213_),
    .Z(_02783_));
 OAI22_X2 _39760_ (.A1(_00165_),
    .A2(_15209_),
    .B1(_15178_),
    .B2(_00030_),
    .ZN(_15214_));
 MUX2_X1 _39761_ (.A(_12919_),
    .B(_15214_),
    .S(_15213_),
    .Z(_02784_));
 OAI22_X1 _39762_ (.A1(_12189_),
    .A2(_15209_),
    .B1(_15178_),
    .B2(_00033_),
    .ZN(_15215_));
 MUX2_X1 _39763_ (.A(\core.keymem.prev_key0_reg[125] ),
    .B(_15215_),
    .S(_15213_),
    .Z(_02785_));
 OAI22_X1 _39764_ (.A1(_00169_),
    .A2(_15209_),
    .B1(_15178_),
    .B2(_00036_),
    .ZN(_15216_));
 MUX2_X1 _39765_ (.A(_12200_),
    .B(_15216_),
    .S(_15213_),
    .Z(_02786_));
 OAI21_X1 _39766_ (.A(_12934_),
    .B1(_15169_),
    .B2(_00039_),
    .ZN(_15217_));
 MUX2_X1 _39767_ (.A(_12936_),
    .B(_15217_),
    .S(_15213_),
    .Z(_02787_));
 NOR2_X1 _39768_ (.A1(\core.keymem.prev_key0_reg[12] ),
    .A2(_15182_),
    .ZN(_15218_));
 BUF_X4 _39769_ (.A(_15159_),
    .Z(_15219_));
 AOI21_X1 _39770_ (.A(_12948_),
    .B1(_15219_),
    .B2(_07313_),
    .ZN(_15220_));
 BUF_X4 _39771_ (.A(_15162_),
    .Z(_15221_));
 AOI21_X1 _39772_ (.A(_15218_),
    .B1(_15220_),
    .B2(_15221_),
    .ZN(_02788_));
 OAI21_X1 _39773_ (.A(_14283_),
    .B1(_15169_),
    .B2(_00384_),
    .ZN(_15222_));
 MUX2_X1 _39774_ (.A(\core.keymem.prev_key0_reg[13] ),
    .B(_15222_),
    .S(_15213_),
    .Z(_02789_));
 OAI22_X1 _39775_ (.A1(_00409_),
    .A2(_15209_),
    .B1(_15178_),
    .B2(_00387_),
    .ZN(_15223_));
 MUX2_X1 _39776_ (.A(_12978_),
    .B(_15223_),
    .S(_15213_),
    .Z(_02790_));
 OAI21_X1 _39777_ (.A(_14305_),
    .B1(_15164_),
    .B2(_00390_),
    .ZN(_15224_));
 MUX2_X1 _39778_ (.A(\core.keymem.prev_key0_reg[15] ),
    .B(_15224_),
    .S(_15213_),
    .Z(_02791_));
 BUF_X4 _39779_ (.A(_13136_),
    .Z(_15225_));
 OAI22_X1 _39780_ (.A1(_00411_),
    .A2(_15209_),
    .B1(_15225_),
    .B2(_08253_),
    .ZN(_15226_));
 MUX2_X1 _39781_ (.A(\core.keymem.prev_key0_reg[16] ),
    .B(_15226_),
    .S(_15213_),
    .Z(_02792_));
 OAI22_X1 _39782_ (.A1(_00434_),
    .A2(_15209_),
    .B1(_15225_),
    .B2(_08192_),
    .ZN(_15227_));
 MUX2_X1 _39783_ (.A(\core.keymem.prev_key0_reg[17] ),
    .B(_15227_),
    .S(_15213_),
    .Z(_02793_));
 OAI22_X1 _39784_ (.A1(_00435_),
    .A2(_15209_),
    .B1(_15225_),
    .B2(_08214_),
    .ZN(_15228_));
 BUF_X4 _39785_ (.A(_15154_),
    .Z(_15229_));
 MUX2_X1 _39786_ (.A(_13044_),
    .B(_15228_),
    .S(_15229_),
    .Z(_02794_));
 OAI22_X1 _39787_ (.A1(_00436_),
    .A2(_15209_),
    .B1(_15225_),
    .B2(_08205_),
    .ZN(_15230_));
 MUX2_X1 _39788_ (.A(\core.keymem.prev_key0_reg[19] ),
    .B(_15230_),
    .S(_15229_),
    .Z(_02795_));
 BUF_X4 _39789_ (.A(_12871_),
    .Z(_15231_));
 OAI22_X1 _39790_ (.A1(_00371_),
    .A2(_15231_),
    .B1(_15225_),
    .B2(_06796_),
    .ZN(_15232_));
 MUX2_X1 _39791_ (.A(\core.keymem.prev_key0_reg[1] ),
    .B(_15232_),
    .S(_15229_),
    .Z(_02796_));
 OAI21_X1 _39792_ (.A(_14325_),
    .B1(_15164_),
    .B2(_08318_),
    .ZN(_15233_));
 MUX2_X1 _39793_ (.A(\core.keymem.prev_key0_reg[20] ),
    .B(_15233_),
    .S(_15229_),
    .Z(_02797_));
 NOR2_X1 _39794_ (.A1(\core.keymem.prev_key0_reg[21] ),
    .A2(_15182_),
    .ZN(_15234_));
 AOI21_X1 _39795_ (.A(_14329_),
    .B1(_15219_),
    .B2(_08231_),
    .ZN(_15235_));
 AOI21_X1 _39796_ (.A(_15234_),
    .B1(_15235_),
    .B2(_15221_),
    .ZN(_02798_));
 OAI21_X1 _39797_ (.A(_14332_),
    .B1(_15164_),
    .B2(_00417_),
    .ZN(_15236_));
 MUX2_X1 _39798_ (.A(\core.keymem.prev_key0_reg[22] ),
    .B(_15236_),
    .S(_15229_),
    .Z(_02799_));
 OAI22_X1 _39799_ (.A1(_00016_),
    .A2(_15231_),
    .B1(_15225_),
    .B2(_00420_),
    .ZN(_15237_));
 MUX2_X1 _39800_ (.A(\core.keymem.prev_key0_reg[23] ),
    .B(_15237_),
    .S(_15229_),
    .Z(_02800_));
 NOR2_X1 _39801_ (.A1(\core.keymem.prev_key0_reg[24] ),
    .A2(_15182_),
    .ZN(_15238_));
 AOI21_X1 _39802_ (.A(_13210_),
    .B1(_15219_),
    .B2(_09318_),
    .ZN(_15239_));
 AOI21_X1 _39803_ (.A(_15238_),
    .B1(_15239_),
    .B2(_15221_),
    .ZN(_02801_));
 OAI22_X1 _39804_ (.A1(_00020_),
    .A2(_15231_),
    .B1(_15225_),
    .B2(_09308_),
    .ZN(_15240_));
 MUX2_X1 _39805_ (.A(\core.keymem.prev_key0_reg[25] ),
    .B(_15240_),
    .S(_15229_),
    .Z(_02802_));
 OAI22_X1 _39806_ (.A1(_00023_),
    .A2(_15231_),
    .B1(_15225_),
    .B2(_09238_),
    .ZN(_15241_));
 MUX2_X1 _39807_ (.A(\core.keymem.prev_key0_reg[26] ),
    .B(_15241_),
    .S(_15229_),
    .Z(_02803_));
 OAI22_X1 _39808_ (.A1(_00026_),
    .A2(_15231_),
    .B1(_15225_),
    .B2(_09229_),
    .ZN(_15242_));
 MUX2_X1 _39809_ (.A(\core.keymem.prev_key0_reg[27] ),
    .B(_15242_),
    .S(_15229_),
    .Z(_02804_));
 BUF_X4 _39810_ (.A(_15155_),
    .Z(_15243_));
 NOR2_X1 _39811_ (.A1(\core.keymem.prev_key0_reg[28] ),
    .A2(_15243_),
    .ZN(_15244_));
 AOI21_X1 _39812_ (.A(_13316_),
    .B1(_15219_),
    .B2(_09282_),
    .ZN(_15245_));
 AOI21_X1 _39813_ (.A(_15244_),
    .B1(_15245_),
    .B2(_15221_),
    .ZN(_02805_));
 NOR2_X1 _39814_ (.A1(\core.keymem.prev_key0_reg[29] ),
    .A2(_15243_),
    .ZN(_15246_));
 AOI21_X1 _39815_ (.A(_12291_),
    .B1(_15219_),
    .B2(_09273_),
    .ZN(_15247_));
 AOI21_X1 _39816_ (.A(_15246_),
    .B1(_15247_),
    .B2(_15221_),
    .ZN(_02806_));
 OAI22_X1 _39817_ (.A1(_00373_),
    .A2(_15231_),
    .B1(_15225_),
    .B2(_06783_),
    .ZN(_15248_));
 MUX2_X1 _39818_ (.A(\core.keymem.prev_key0_reg[2] ),
    .B(_15248_),
    .S(_15229_),
    .Z(_02807_));
 BUF_X4 _39819_ (.A(_13136_),
    .Z(_15249_));
 OAI22_X1 _39820_ (.A1(_00035_),
    .A2(_15231_),
    .B1(_15249_),
    .B2(_00335_),
    .ZN(_15250_));
 BUF_X4 _39821_ (.A(_15154_),
    .Z(_15251_));
 MUX2_X1 _39822_ (.A(\core.keymem.prev_key0_reg[30] ),
    .B(_15250_),
    .S(_15251_),
    .Z(_02808_));
 OAI22_X1 _39823_ (.A1(_00038_),
    .A2(_15231_),
    .B1(_15249_),
    .B2(_00338_),
    .ZN(_15252_));
 MUX2_X1 _39824_ (.A(\core.keymem.prev_key0_reg[31] ),
    .B(_15252_),
    .S(_15251_),
    .Z(_02809_));
 NOR2_X1 _39825_ (.A1(\core.keymem.prev_key0_reg[32] ),
    .A2(_15243_),
    .ZN(_15253_));
 NOR2_X1 _39826_ (.A1(_00041_),
    .A2(_12262_),
    .ZN(_15254_));
 AOI21_X1 _39827_ (.A(_15254_),
    .B1(_15219_),
    .B2(\core.keymem.prev_key1_reg[32] ),
    .ZN(_15255_));
 AOI21_X1 _39828_ (.A(_15253_),
    .B1(_15255_),
    .B2(_15221_),
    .ZN(_02810_));
 NOR2_X1 _39829_ (.A1(_13117_),
    .A2(_15243_),
    .ZN(_15256_));
 AOI21_X1 _39830_ (.A(_12357_),
    .B1(_15219_),
    .B2(\core.keymem.prev_key1_reg[33] ),
    .ZN(_15257_));
 AOI21_X1 _39831_ (.A(_15256_),
    .B1(_15257_),
    .B2(_15221_),
    .ZN(_02811_));
 NOR2_X1 _39832_ (.A1(\core.keymem.prev_key0_reg[34] ),
    .A2(_15243_),
    .ZN(_15258_));
 AOI21_X1 _39833_ (.A(_12363_),
    .B1(_15219_),
    .B2(\core.keymem.prev_key1_reg[34] ),
    .ZN(_15259_));
 AOI21_X1 _39834_ (.A(_15258_),
    .B1(_15259_),
    .B2(_15221_),
    .ZN(_02812_));
 NOR2_X1 _39835_ (.A1(_12383_),
    .A2(_15243_),
    .ZN(_15260_));
 AOI21_X1 _39836_ (.A(_12408_),
    .B1(_15219_),
    .B2(\core.keymem.prev_key1_reg[35] ),
    .ZN(_15261_));
 AOI21_X1 _39837_ (.A(_15260_),
    .B1(_15261_),
    .B2(_15221_),
    .ZN(_02813_));
 NOR2_X1 _39838_ (.A1(\core.keymem.prev_key0_reg[36] ),
    .A2(_15243_),
    .ZN(_15262_));
 AOI21_X1 _39839_ (.A(_12414_),
    .B1(_15219_),
    .B2(\core.keymem.prev_key1_reg[36] ),
    .ZN(_15263_));
 AOI21_X1 _39840_ (.A(_15262_),
    .B1(_15263_),
    .B2(_15221_),
    .ZN(_02814_));
 NOR2_X1 _39841_ (.A1(\core.keymem.prev_key0_reg[37] ),
    .A2(_15243_),
    .ZN(_15264_));
 BUF_X4 _39842_ (.A(_15159_),
    .Z(_15265_));
 AOI21_X1 _39843_ (.A(_12432_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[37] ),
    .ZN(_15266_));
 BUF_X4 _39844_ (.A(_15162_),
    .Z(_15267_));
 AOI21_X1 _39845_ (.A(_15264_),
    .B1(_15266_),
    .B2(_15267_),
    .ZN(_02815_));
 NOR2_X1 _39846_ (.A1(_12442_),
    .A2(_15243_),
    .ZN(_15268_));
 AOI21_X1 _39847_ (.A(_12463_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[38] ),
    .ZN(_15269_));
 AOI21_X1 _39848_ (.A(_15268_),
    .B1(_15269_),
    .B2(_15267_),
    .ZN(_02816_));
 INV_X1 _39849_ (.A(\core.keymem.prev_key1_reg[39] ),
    .ZN(_15270_));
 OAI22_X1 _39850_ (.A1(_00048_),
    .A2(_15231_),
    .B1(_15249_),
    .B2(_15270_),
    .ZN(_15271_));
 MUX2_X1 _39851_ (.A(_13417_),
    .B(_15271_),
    .S(_15251_),
    .Z(_02817_));
 OAI22_X1 _39852_ (.A1(_00374_),
    .A2(_15231_),
    .B1(_15249_),
    .B2(_06708_),
    .ZN(_15272_));
 MUX2_X1 _39853_ (.A(\core.keymem.prev_key0_reg[3] ),
    .B(_15272_),
    .S(_15251_),
    .Z(_02818_));
 NOR2_X1 _39854_ (.A1(_13451_),
    .A2(_15243_),
    .ZN(_15273_));
 NOR2_X1 _39855_ (.A1(_00049_),
    .A2(_12158_),
    .ZN(_15274_));
 AOI21_X1 _39856_ (.A(_15274_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[40] ),
    .ZN(_15275_));
 AOI21_X1 _39857_ (.A(_15273_),
    .B1(_15275_),
    .B2(_15267_),
    .ZN(_02819_));
 BUF_X4 _39858_ (.A(_15155_),
    .Z(_15276_));
 NOR2_X1 _39859_ (.A1(\core.keymem.prev_key0_reg[41] ),
    .A2(_15276_),
    .ZN(_15277_));
 AOI21_X1 _39860_ (.A(_13458_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[41] ),
    .ZN(_15278_));
 AOI21_X1 _39861_ (.A(_15277_),
    .B1(_15278_),
    .B2(_15267_),
    .ZN(_02820_));
 NOR2_X1 _39862_ (.A1(_12845_),
    .A2(_15276_),
    .ZN(_15279_));
 NOR2_X2 _39863_ (.A1(_00051_),
    .A2(_13875_),
    .ZN(_15280_));
 AOI21_X2 _39864_ (.A(_15280_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[42] ),
    .ZN(_15281_));
 AOI21_X1 _39865_ (.A(_15279_),
    .B1(_15281_),
    .B2(_15267_),
    .ZN(_02821_));
 NOR2_X1 _39866_ (.A1(\core.keymem.prev_key0_reg[43] ),
    .A2(_15276_),
    .ZN(_15282_));
 NOR2_X1 _39867_ (.A1(_00052_),
    .A2(_12185_),
    .ZN(_15283_));
 AOI21_X1 _39868_ (.A(_15283_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[43] ),
    .ZN(_15284_));
 AOI21_X1 _39869_ (.A(_15282_),
    .B1(_15284_),
    .B2(_15267_),
    .ZN(_02822_));
 NOR2_X1 _39870_ (.A1(_12481_),
    .A2(_15276_),
    .ZN(_15285_));
 AOI21_X2 _39871_ (.A(_12500_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[44] ),
    .ZN(_15286_));
 AOI21_X1 _39872_ (.A(_15285_),
    .B1(_15286_),
    .B2(_15267_),
    .ZN(_02823_));
 NOR2_X1 _39873_ (.A1(_12962_),
    .A2(_15276_),
    .ZN(_15287_));
 NOR2_X1 _39874_ (.A1(_00054_),
    .A2(_14447_),
    .ZN(_15288_));
 AOI21_X1 _39875_ (.A(_15288_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[45] ),
    .ZN(_15289_));
 AOI21_X1 _39876_ (.A(_15287_),
    .B1(_15289_),
    .B2(_15267_),
    .ZN(_02824_));
 NOR2_X1 _39877_ (.A1(_12979_),
    .A2(_15276_),
    .ZN(_15290_));
 NOR2_X1 _39878_ (.A1(_00055_),
    .A2(_12186_),
    .ZN(_15291_));
 AOI21_X1 _39879_ (.A(_15291_),
    .B1(_15265_),
    .B2(_12987_),
    .ZN(_15292_));
 AOI21_X1 _39880_ (.A(_15290_),
    .B1(_15292_),
    .B2(_15267_),
    .ZN(_02825_));
 NOR2_X1 _39881_ (.A1(\core.keymem.prev_key0_reg[47] ),
    .A2(_15276_),
    .ZN(_15293_));
 NOR2_X1 _39882_ (.A1(_00056_),
    .A2(_12262_),
    .ZN(_15294_));
 AOI21_X1 _39883_ (.A(_15294_),
    .B1(_15265_),
    .B2(\core.keymem.prev_key1_reg[47] ),
    .ZN(_15295_));
 AOI21_X1 _39884_ (.A(_15293_),
    .B1(_15295_),
    .B2(_15267_),
    .ZN(_02826_));
 NOR2_X1 _39885_ (.A1(\core.keymem.prev_key0_reg[48] ),
    .A2(_15276_),
    .ZN(_15296_));
 BUF_X4 _39886_ (.A(_13011_),
    .Z(_15297_));
 AOI21_X1 _39887_ (.A(_12525_),
    .B1(_15297_),
    .B2(_12526_),
    .ZN(_15298_));
 BUF_X4 _39888_ (.A(_15162_),
    .Z(_15299_));
 AOI21_X1 _39889_ (.A(_15296_),
    .B1(_15298_),
    .B2(_15299_),
    .ZN(_02827_));
 BUF_X4 _39890_ (.A(_12871_),
    .Z(_15300_));
 OAI22_X1 _39891_ (.A1(_00058_),
    .A2(_15300_),
    .B1(_15249_),
    .B2(_13525_),
    .ZN(_15301_));
 MUX2_X1 _39892_ (.A(\core.keymem.prev_key0_reg[49] ),
    .B(_15301_),
    .S(_15251_),
    .Z(_02828_));
 NOR2_X1 _39893_ (.A1(\core.keymem.prev_key0_reg[4] ),
    .A2(_15276_),
    .ZN(_15302_));
 AOI21_X1 _39894_ (.A(_14395_),
    .B1(_15297_),
    .B2(_06775_),
    .ZN(_15303_));
 AOI21_X1 _39895_ (.A(_15302_),
    .B1(_15303_),
    .B2(_15299_),
    .ZN(_02829_));
 OAI22_X2 _39896_ (.A1(_00059_),
    .A2(_15300_),
    .B1(_15249_),
    .B2(_13088_),
    .ZN(_15304_));
 MUX2_X1 _39897_ (.A(_13046_),
    .B(_15304_),
    .S(_15251_),
    .Z(_02830_));
 NOR2_X1 _39898_ (.A1(\core.keymem.prev_key0_reg[51] ),
    .A2(_15276_),
    .ZN(_15305_));
 AOI21_X1 _39899_ (.A(_13558_),
    .B1(_15297_),
    .B2(\core.keymem.prev_key1_reg[51] ),
    .ZN(_15306_));
 AOI21_X1 _39900_ (.A(_15305_),
    .B1(_15306_),
    .B2(_15299_),
    .ZN(_02831_));
 BUF_X4 _39901_ (.A(_15155_),
    .Z(_15307_));
 NOR2_X1 _39902_ (.A1(_12548_),
    .A2(_15307_),
    .ZN(_15308_));
 AOI21_X1 _39903_ (.A(_12542_),
    .B1(_15297_),
    .B2(\core.keymem.prev_key1_reg[52] ),
    .ZN(_15309_));
 AOI21_X1 _39904_ (.A(_15308_),
    .B1(_15309_),
    .B2(_15299_),
    .ZN(_02832_));
 NOR2_X1 _39905_ (.A1(\core.keymem.prev_key0_reg[53] ),
    .A2(_15307_),
    .ZN(_15310_));
 AOI21_X1 _39906_ (.A(_12576_),
    .B1(_15297_),
    .B2(\core.keymem.prev_key1_reg[53] ),
    .ZN(_15311_));
 AOI21_X1 _39907_ (.A(_15310_),
    .B1(_15311_),
    .B2(_15299_),
    .ZN(_02833_));
 NOR2_X1 _39908_ (.A1(_13172_),
    .A2(_15307_),
    .ZN(_15312_));
 AOI21_X1 _39909_ (.A(_13571_),
    .B1(_15297_),
    .B2(_13158_),
    .ZN(_15313_));
 AOI21_X1 _39910_ (.A(_15312_),
    .B1(_15313_),
    .B2(_15299_),
    .ZN(_02834_));
 INV_X1 _39911_ (.A(\core.keymem.prev_key1_reg[55] ),
    .ZN(_15314_));
 OAI22_X2 _39912_ (.A1(_00064_),
    .A2(_15300_),
    .B1(_15249_),
    .B2(_15314_),
    .ZN(_15315_));
 MUX2_X1 _39913_ (.A(_12242_),
    .B(_15315_),
    .S(_15251_),
    .Z(_02835_));
 INV_X1 _39914_ (.A(\core.keymem.prev_key1_reg[56] ),
    .ZN(_15316_));
 OAI22_X1 _39915_ (.A1(_00065_),
    .A2(_15300_),
    .B1(_15249_),
    .B2(_15316_),
    .ZN(_15317_));
 MUX2_X1 _39916_ (.A(\core.keymem.prev_key0_reg[56] ),
    .B(_15317_),
    .S(_15251_),
    .Z(_02836_));
 INV_X1 _39917_ (.A(\core.keymem.prev_key1_reg[57] ),
    .ZN(_15318_));
 OAI22_X1 _39918_ (.A1(_00067_),
    .A2(_15300_),
    .B1(_15249_),
    .B2(_15318_),
    .ZN(_15319_));
 MUX2_X1 _39919_ (.A(_13221_),
    .B(_15319_),
    .S(_15251_),
    .Z(_02837_));
 NOR2_X1 _39920_ (.A1(\core.keymem.prev_key0_reg[58] ),
    .A2(_15307_),
    .ZN(_15320_));
 AOI21_X1 _39921_ (.A(_14419_),
    .B1(_15297_),
    .B2(\core.keymem.prev_key1_reg[58] ),
    .ZN(_15321_));
 AOI21_X1 _39922_ (.A(_15320_),
    .B1(_15321_),
    .B2(_15299_),
    .ZN(_02838_));
 NOR2_X1 _39923_ (.A1(_13242_),
    .A2(_15307_),
    .ZN(_15322_));
 AOI21_X1 _39924_ (.A(_14423_),
    .B1(_15297_),
    .B2(\core.keymem.prev_key1_reg[59] ),
    .ZN(_15323_));
 AOI21_X1 _39925_ (.A(_15322_),
    .B1(_15323_),
    .B2(_15299_),
    .ZN(_02839_));
 OR2_X1 _39926_ (.A1(_00376_),
    .A2(_11863_),
    .ZN(_15324_));
 OAI21_X1 _39927_ (.A(_15324_),
    .B1(_15164_),
    .B2(_06778_),
    .ZN(_15325_));
 MUX2_X1 _39928_ (.A(\core.keymem.prev_key0_reg[5] ),
    .B(_15325_),
    .S(_15251_),
    .Z(_02840_));
 NOR2_X1 _39929_ (.A1(\core.keymem.prev_key0_reg[60] ),
    .A2(_15307_),
    .ZN(_15326_));
 AOI21_X1 _39930_ (.A(_14427_),
    .B1(_15297_),
    .B2(\core.keymem.prev_key1_reg[60] ),
    .ZN(_15327_));
 AOI21_X1 _39931_ (.A(_15326_),
    .B1(_15327_),
    .B2(_15299_),
    .ZN(_02841_));
 NOR2_X1 _39932_ (.A1(\core.keymem.prev_key0_reg[61] ),
    .A2(_15307_),
    .ZN(_15328_));
 NOR2_X1 _39933_ (.A1(_00075_),
    .A2(_11875_),
    .ZN(_15329_));
 AOI21_X1 _39934_ (.A(_15329_),
    .B1(_15297_),
    .B2(\core.keymem.prev_key1_reg[61] ),
    .ZN(_15330_));
 AOI21_X1 _39935_ (.A(_15328_),
    .B1(_15330_),
    .B2(_15299_),
    .ZN(_02842_));
 NOR2_X1 _39936_ (.A1(_13342_),
    .A2(_15307_),
    .ZN(_15331_));
 AOI22_X1 _39937_ (.A1(_12610_),
    .A2(_14238_),
    .B1(_15159_),
    .B2(\core.keymem.prev_key1_reg[62] ),
    .ZN(_15332_));
 BUF_X4 _39938_ (.A(_15162_),
    .Z(_15333_));
 AOI21_X1 _39939_ (.A(_15331_),
    .B1(_15332_),
    .B2(_15333_),
    .ZN(_02843_));
 NOR2_X1 _39940_ (.A1(\core.keymem.prev_key0_reg[63] ),
    .A2(_15307_),
    .ZN(_15334_));
 BUF_X4 _39941_ (.A(_13011_),
    .Z(_15335_));
 AOI21_X1 _39942_ (.A(_14441_),
    .B1(_15335_),
    .B2(\core.keymem.prev_key1_reg[63] ),
    .ZN(_15336_));
 AOI21_X1 _39943_ (.A(_15334_),
    .B1(_15336_),
    .B2(_15333_),
    .ZN(_02844_));
 OAI22_X1 _39944_ (.A1(_00081_),
    .A2(_15300_),
    .B1(_15249_),
    .B2(_12615_),
    .ZN(_15337_));
 BUF_X4 _39945_ (.A(_15154_),
    .Z(_15338_));
 MUX2_X1 _39946_ (.A(\core.keymem.prev_key0_reg[64] ),
    .B(_15337_),
    .S(_15338_),
    .Z(_02845_));
 BUF_X4 _39947_ (.A(_13136_),
    .Z(_15339_));
 OAI22_X1 _39948_ (.A1(_00082_),
    .A2(_15300_),
    .B1(_15339_),
    .B2(_13662_),
    .ZN(_15340_));
 MUX2_X1 _39949_ (.A(_13118_),
    .B(_15340_),
    .S(_15338_),
    .Z(_02846_));
 NOR2_X1 _39950_ (.A1(_12325_),
    .A2(_15307_),
    .ZN(_15341_));
 AOI21_X1 _39951_ (.A(_14448_),
    .B1(_15335_),
    .B2(\core.keymem.prev_key1_reg[66] ),
    .ZN(_15342_));
 AOI21_X1 _39952_ (.A(_15341_),
    .B1(_15342_),
    .B2(_15333_),
    .ZN(_02847_));
 BUF_X4 _39953_ (.A(_15155_),
    .Z(_15343_));
 NOR2_X1 _39954_ (.A1(_12384_),
    .A2(_15343_),
    .ZN(_15344_));
 NOR2_X1 _39955_ (.A1(_00084_),
    .A2(_12262_),
    .ZN(_15345_));
 AOI21_X1 _39956_ (.A(_15345_),
    .B1(_15335_),
    .B2(\core.keymem.prev_key1_reg[67] ),
    .ZN(_15346_));
 AOI21_X1 _39957_ (.A(_15344_),
    .B1(_15346_),
    .B2(_15333_),
    .ZN(_02848_));
 NOR2_X1 _39958_ (.A1(\core.keymem.prev_key0_reg[68] ),
    .A2(_15343_),
    .ZN(_15347_));
 NOR2_X1 _39959_ (.A1(_00085_),
    .A2(_11885_),
    .ZN(_15348_));
 AOI21_X1 _39960_ (.A(_15348_),
    .B1(_15335_),
    .B2(\core.keymem.prev_key1_reg[68] ),
    .ZN(_15349_));
 AOI21_X1 _39961_ (.A(_15347_),
    .B1(_15349_),
    .B2(_15333_),
    .ZN(_02849_));
 NOR2_X1 _39962_ (.A1(\core.keymem.prev_key0_reg[69] ),
    .A2(_15343_),
    .ZN(_15350_));
 NOR2_X1 _39963_ (.A1(_00086_),
    .A2(_14447_),
    .ZN(_15351_));
 AOI21_X1 _39964_ (.A(_15351_),
    .B1(_15335_),
    .B2(_12434_),
    .ZN(_15352_));
 AOI21_X1 _39965_ (.A(_15350_),
    .B1(_15352_),
    .B2(_15333_),
    .ZN(_02850_));
 OAI21_X1 _39966_ (.A(_13709_),
    .B1(_15164_),
    .B2(_00354_),
    .ZN(_15353_));
 MUX2_X1 _39967_ (.A(\core.keymem.prev_key0_reg[6] ),
    .B(_15353_),
    .S(_15338_),
    .Z(_02851_));
 NOR2_X1 _39968_ (.A1(_12443_),
    .A2(_15343_),
    .ZN(_15354_));
 AOI21_X1 _39969_ (.A(_12642_),
    .B1(_15335_),
    .B2(_12464_),
    .ZN(_15355_));
 AOI21_X1 _39970_ (.A(_15354_),
    .B1(_15355_),
    .B2(_15333_),
    .ZN(_02852_));
 NOR2_X1 _39971_ (.A1(_12653_),
    .A2(_15343_),
    .ZN(_15356_));
 NOR2_X1 _39972_ (.A1(_00088_),
    .A2(_12002_),
    .ZN(_15357_));
 AOI21_X1 _39973_ (.A(_15357_),
    .B1(_15335_),
    .B2(\core.keymem.prev_key1_reg[71] ),
    .ZN(_15358_));
 AOI21_X1 _39974_ (.A(_15356_),
    .B1(_15358_),
    .B2(_15333_),
    .ZN(_02853_));
 NOR2_X1 _39975_ (.A1(_12666_),
    .A2(_15343_),
    .ZN(_15359_));
 AOI21_X1 _39976_ (.A(_12661_),
    .B1(_15335_),
    .B2(\core.keymem.prev_key1_reg[72] ),
    .ZN(_15360_));
 AOI21_X1 _39977_ (.A(_15359_),
    .B1(_15360_),
    .B2(_15333_),
    .ZN(_02854_));
 INV_X1 _39978_ (.A(_12683_),
    .ZN(_15361_));
 OAI22_X1 _39979_ (.A1(_00090_),
    .A2(_15300_),
    .B1(_15339_),
    .B2(_15361_),
    .ZN(_15362_));
 MUX2_X1 _39980_ (.A(\core.keymem.prev_key0_reg[73] ),
    .B(_15362_),
    .S(_15338_),
    .Z(_02855_));
 NOR2_X1 _39981_ (.A1(_12846_),
    .A2(_15343_),
    .ZN(_15363_));
 AOI21_X2 _39982_ (.A(_14463_),
    .B1(_15335_),
    .B2(\core.keymem.prev_key1_reg[74] ),
    .ZN(_15364_));
 AOI21_X1 _39983_ (.A(_15363_),
    .B1(_15364_),
    .B2(_15333_),
    .ZN(_02856_));
 NOR2_X1 _39984_ (.A1(\core.keymem.prev_key0_reg[75] ),
    .A2(_15343_),
    .ZN(_15365_));
 NOR2_X1 _39985_ (.A1(_00092_),
    .A2(_11885_),
    .ZN(_15366_));
 AOI21_X1 _39986_ (.A(_15366_),
    .B1(_15335_),
    .B2(\core.keymem.prev_key1_reg[75] ),
    .ZN(_15367_));
 BUF_X4 _39987_ (.A(_15155_),
    .Z(_15368_));
 AOI21_X1 _39988_ (.A(_15365_),
    .B1(_15367_),
    .B2(_15368_),
    .ZN(_02857_));
 INV_X1 _39989_ (.A(\core.keymem.prev_key1_reg[76] ),
    .ZN(_15369_));
 OAI22_X2 _39990_ (.A1(_00093_),
    .A2(_15300_),
    .B1(_15339_),
    .B2(_15369_),
    .ZN(_15370_));
 MUX2_X1 _39991_ (.A(_12482_),
    .B(_15370_),
    .S(_15338_),
    .Z(_02858_));
 NOR2_X1 _39992_ (.A1(_12960_),
    .A2(_15343_),
    .ZN(_15371_));
 BUF_X4 _39993_ (.A(_13011_),
    .Z(_15372_));
 AOI21_X1 _39994_ (.A(_13743_),
    .B1(_15372_),
    .B2(\core.keymem.prev_key1_reg[77] ),
    .ZN(_15373_));
 AOI21_X1 _39995_ (.A(_15371_),
    .B1(_15373_),
    .B2(_15368_),
    .ZN(_02859_));
 NOR2_X1 _39996_ (.A1(_12698_),
    .A2(_15343_),
    .ZN(_15374_));
 NOR2_X1 _39997_ (.A1(_00095_),
    .A2(_13720_),
    .ZN(_15375_));
 AOI21_X1 _39998_ (.A(_15375_),
    .B1(_15372_),
    .B2(_12701_),
    .ZN(_15376_));
 AOI21_X1 _39999_ (.A(_15374_),
    .B1(_15376_),
    .B2(_15368_),
    .ZN(_02860_));
 BUF_X4 _40000_ (.A(_15155_),
    .Z(_15377_));
 NOR2_X1 _40001_ (.A1(\core.keymem.prev_key0_reg[79] ),
    .A2(_15377_),
    .ZN(_15378_));
 AOI21_X1 _40002_ (.A(_14475_),
    .B1(_15372_),
    .B2(\core.keymem.prev_key1_reg[79] ),
    .ZN(_15379_));
 AOI21_X1 _40003_ (.A(_15378_),
    .B1(_15379_),
    .B2(_15368_),
    .ZN(_02861_));
 OAI22_X2 _40004_ (.A1(_00380_),
    .A2(_15300_),
    .B1(_15339_),
    .B2(_00357_),
    .ZN(_15380_));
 MUX2_X1 _40005_ (.A(\core.keymem.prev_key0_reg[7] ),
    .B(_15380_),
    .S(_15338_),
    .Z(_02862_));
 INV_X1 _40006_ (.A(_12527_),
    .ZN(_15381_));
 OAI22_X1 _40007_ (.A1(_00097_),
    .A2(_14488_),
    .B1(_15339_),
    .B2(_15381_),
    .ZN(_15382_));
 MUX2_X1 _40008_ (.A(\core.keymem.prev_key0_reg[80] ),
    .B(_15382_),
    .S(_15338_),
    .Z(_02863_));
 NOR2_X1 _40009_ (.A1(\core.keymem.prev_key0_reg[81] ),
    .A2(_15377_),
    .ZN(_15383_));
 NOR2_X1 _40010_ (.A1(_00098_),
    .A2(_12834_),
    .ZN(_15384_));
 AOI21_X1 _40011_ (.A(_15384_),
    .B1(_15372_),
    .B2(\core.keymem.prev_key1_reg[81] ),
    .ZN(_15385_));
 AOI21_X1 _40012_ (.A(_15383_),
    .B1(_15385_),
    .B2(_15368_),
    .ZN(_02864_));
 NOR2_X1 _40013_ (.A1(_13048_),
    .A2(_15377_),
    .ZN(_15386_));
 NOR2_X1 _40014_ (.A1(_00099_),
    .A2(_13331_),
    .ZN(_15387_));
 AOI21_X1 _40015_ (.A(_15387_),
    .B1(_15372_),
    .B2(\core.keymem.prev_key1_reg[82] ),
    .ZN(_15388_));
 AOI21_X1 _40016_ (.A(_15386_),
    .B1(_15388_),
    .B2(_15368_),
    .ZN(_02865_));
 NOR2_X1 _40017_ (.A1(\core.keymem.prev_key0_reg[83] ),
    .A2(_15377_),
    .ZN(_15389_));
 AOI21_X1 _40018_ (.A(_13785_),
    .B1(_15372_),
    .B2(\core.keymem.prev_key1_reg[83] ),
    .ZN(_15390_));
 AOI21_X1 _40019_ (.A(_15389_),
    .B1(_15390_),
    .B2(_15368_),
    .ZN(_02866_));
 NOR2_X1 _40020_ (.A1(_12549_),
    .A2(_15377_),
    .ZN(_15391_));
 AOI21_X1 _40021_ (.A(_12721_),
    .B1(_15372_),
    .B2(\core.keymem.prev_key1_reg[84] ),
    .ZN(_15392_));
 AOI21_X1 _40022_ (.A(_15391_),
    .B1(_15392_),
    .B2(_15368_),
    .ZN(_02867_));
 NOR2_X1 _40023_ (.A1(\core.keymem.prev_key0_reg[85] ),
    .A2(_15377_),
    .ZN(_15393_));
 AOI21_X1 _40024_ (.A(_13793_),
    .B1(_15372_),
    .B2(_12579_),
    .ZN(_15394_));
 AOI21_X1 _40025_ (.A(_15393_),
    .B1(_15394_),
    .B2(_15368_),
    .ZN(_02868_));
 NOR2_X1 _40026_ (.A1(_12732_),
    .A2(_15377_),
    .ZN(_15395_));
 NOR2_X1 _40027_ (.A1(_00103_),
    .A2(_14447_),
    .ZN(_15396_));
 AOI21_X1 _40028_ (.A(_15396_),
    .B1(_15372_),
    .B2(_12727_),
    .ZN(_15397_));
 AOI21_X1 _40029_ (.A(_15395_),
    .B1(_15397_),
    .B2(_15368_),
    .ZN(_02869_));
 NOR2_X1 _40030_ (.A1(_12244_),
    .A2(_15377_),
    .ZN(_15398_));
 AOI21_X1 _40031_ (.A(_14487_),
    .B1(_15372_),
    .B2(\core.keymem.prev_key1_reg[87] ),
    .ZN(_15399_));
 AOI21_X1 _40032_ (.A(_15398_),
    .B1(_15399_),
    .B2(_15156_),
    .ZN(_02870_));
 NOR2_X1 _40033_ (.A1(\core.keymem.prev_key0_reg[88] ),
    .A2(_15377_),
    .ZN(_15400_));
 NOR2_X2 _40034_ (.A1(_00105_),
    .A2(_12186_),
    .ZN(_15401_));
 AOI21_X1 _40035_ (.A(_15401_),
    .B1(_15159_),
    .B2(_13204_),
    .ZN(_15402_));
 AOI21_X1 _40036_ (.A(_15400_),
    .B1(_15402_),
    .B2(_15156_),
    .ZN(_02871_));
 INV_X1 _40037_ (.A(_13213_),
    .ZN(_15403_));
 OAI22_X2 _40038_ (.A1(_00107_),
    .A2(_14488_),
    .B1(_15339_),
    .B2(_15403_),
    .ZN(_15404_));
 MUX2_X1 _40039_ (.A(_13223_),
    .B(_15404_),
    .S(_15338_),
    .Z(_02872_));
 NAND2_X1 _40040_ (.A1(_12746_),
    .A2(_12779_),
    .ZN(_15405_));
 OAI21_X1 _40041_ (.A(_15405_),
    .B1(_15164_),
    .B2(_07262_),
    .ZN(_15406_));
 MUX2_X1 _40042_ (.A(_13822_),
    .B(_15406_),
    .S(_15338_),
    .Z(_02873_));
 NOR2_X1 _40043_ (.A1(\core.keymem.prev_key0_reg[90] ),
    .A2(_15377_),
    .ZN(_15407_));
 NOR2_X1 _40044_ (.A1(_00109_),
    .A2(_12834_),
    .ZN(_15408_));
 AOI21_X1 _40045_ (.A(_15408_),
    .B1(_15159_),
    .B2(_12279_),
    .ZN(_15409_));
 AOI21_X1 _40046_ (.A(_15407_),
    .B1(_15409_),
    .B2(_15156_),
    .ZN(_02874_));
 NOR2_X1 _40047_ (.A1(_13244_),
    .A2(_15166_),
    .ZN(_15410_));
 NOR2_X1 _40048_ (.A1(_00111_),
    .A2(_13875_),
    .ZN(_15411_));
 AOI21_X2 _40049_ (.A(_15411_),
    .B1(_15159_),
    .B2(_13277_),
    .ZN(_15412_));
 AOI21_X1 _40050_ (.A(_15410_),
    .B1(_15412_),
    .B2(_15156_),
    .ZN(_02875_));
 OAI22_X4 _40051_ (.A1(_00113_),
    .A2(_14488_),
    .B1(_15339_),
    .B2(_13876_),
    .ZN(_15413_));
 MUX2_X1 _40052_ (.A(_13287_),
    .B(_15413_),
    .S(_15338_),
    .Z(_02876_));
 INV_X1 _40053_ (.A(_12294_),
    .ZN(_15414_));
 OAI22_X1 _40054_ (.A1(_00115_),
    .A2(_14488_),
    .B1(_15339_),
    .B2(_15414_),
    .ZN(_15415_));
 MUX2_X1 _40055_ (.A(_12307_),
    .B(_15415_),
    .S(_15162_),
    .Z(_02877_));
 NOR2_X1 _40056_ (.A1(_13344_),
    .A2(_15166_),
    .ZN(_15416_));
 NOR2_X1 _40057_ (.A1(_00117_),
    .A2(_12185_),
    .ZN(_15417_));
 AOI21_X2 _40058_ (.A(_15417_),
    .B1(_15159_),
    .B2(_13336_),
    .ZN(_15418_));
 AOI21_X1 _40059_ (.A(_15416_),
    .B1(_15418_),
    .B2(_15156_),
    .ZN(_02878_));
 NOR2_X1 _40060_ (.A1(_13382_),
    .A2(_15166_),
    .ZN(_15419_));
 NOR2_X1 _40061_ (.A1(_00119_),
    .A2(_12158_),
    .ZN(_15420_));
 AOI21_X1 _40062_ (.A(_15420_),
    .B1(_15159_),
    .B2(_13387_),
    .ZN(_15421_));
 AOI21_X1 _40063_ (.A(_15419_),
    .B1(_15421_),
    .B2(_15156_),
    .ZN(_02879_));
 OAI22_X1 _40064_ (.A1(_00121_),
    .A2(_14488_),
    .B1(_15339_),
    .B2(_00328_),
    .ZN(_15422_));
 MUX2_X1 _40065_ (.A(\core.keymem.prev_key0_reg[96] ),
    .B(_15422_),
    .S(_15162_),
    .Z(_02880_));
 OAI22_X1 _40066_ (.A1(_00122_),
    .A2(_14488_),
    .B1(_15339_),
    .B2(_00372_),
    .ZN(_15423_));
 MUX2_X1 _40067_ (.A(\core.keymem.prev_key0_reg[97] ),
    .B(_15423_),
    .S(_15162_),
    .Z(_02881_));
 OAI22_X2 _40068_ (.A1(_00123_),
    .A2(_14488_),
    .B1(_13136_),
    .B2(_00124_),
    .ZN(_15424_));
 MUX2_X1 _40069_ (.A(\core.keymem.prev_key0_reg[98] ),
    .B(_15424_),
    .S(_15162_),
    .Z(_02882_));
 OAI21_X1 _40070_ (.A(_12793_),
    .B1(_15164_),
    .B2(_00126_),
    .ZN(_15425_));
 MUX2_X1 _40071_ (.A(_12385_),
    .B(_15425_),
    .S(_15162_),
    .Z(_02883_));
 NOR2_X1 _40072_ (.A1(\core.keymem.prev_key0_reg[9] ),
    .A2(_15166_),
    .ZN(_15426_));
 AOI21_X1 _40073_ (.A(_14532_),
    .B1(_15159_),
    .B2(_07370_),
    .ZN(_15427_));
 AOI21_X1 _40074_ (.A(_15426_),
    .B1(_15427_),
    .B2(_15156_),
    .ZN(_02884_));
 INV_X4 _40075_ (.A(_15153_),
    .ZN(_15428_));
 AOI21_X4 _40076_ (.A(_11803_),
    .B1(_15428_),
    .B2(_11798_),
    .ZN(_15429_));
 BUF_X4 _40077_ (.A(_15429_),
    .Z(_15430_));
 BUF_X4 _40078_ (.A(_15430_),
    .Z(_15431_));
 BUF_X4 _40079_ (.A(_15431_),
    .Z(_15432_));
 BUF_X4 _40080_ (.A(_12786_),
    .Z(_15433_));
 AOI21_X1 _40081_ (.A(_15433_),
    .B1(_11821_),
    .B2(_11839_),
    .ZN(_15434_));
 BUF_X4 _40082_ (.A(_14274_),
    .Z(_15435_));
 AOI21_X1 _40083_ (.A(_15158_),
    .B1(_11810_),
    .B2(_14222_),
    .ZN(_15436_));
 NOR2_X1 _40084_ (.A1(_15435_),
    .A2(_15436_),
    .ZN(_15437_));
 OAI21_X2 _40085_ (.A(_15432_),
    .B1(_15434_),
    .B2(_15437_),
    .ZN(_15438_));
 BUF_X4 _40086_ (.A(_15430_),
    .Z(_15439_));
 BUF_X4 _40087_ (.A(_15439_),
    .Z(_15440_));
 OAI21_X1 _40088_ (.A(_15438_),
    .B1(_15440_),
    .B2(_06859_),
    .ZN(_02885_));
 OAI21_X4 _40089_ (.A(_16228_),
    .B1(_15153_),
    .B2(_11960_),
    .ZN(_15441_));
 BUF_X4 _40090_ (.A(_15441_),
    .Z(_15442_));
 BUF_X4 _40091_ (.A(_15442_),
    .Z(_15443_));
 NAND2_X1 _40092_ (.A1(\core.keymem.prev_key1_reg[100] ),
    .A2(_15443_),
    .ZN(_15444_));
 OAI21_X1 _40093_ (.A(_11870_),
    .B1(_11861_),
    .B2(_14293_),
    .ZN(_15445_));
 BUF_X4 _40094_ (.A(_15441_),
    .Z(_15446_));
 BUF_X4 _40095_ (.A(_15446_),
    .Z(_15447_));
 BUF_X4 _40096_ (.A(_15447_),
    .Z(_15448_));
 OAI21_X1 _40097_ (.A(_15444_),
    .B1(_15445_),
    .B2(_15448_),
    .ZN(_02886_));
 BUF_X4 _40098_ (.A(_12786_),
    .Z(_15449_));
 NOR2_X1 _40099_ (.A1(_00129_),
    .A2(_13331_),
    .ZN(_15450_));
 BUF_X4 _40100_ (.A(_14447_),
    .Z(_15451_));
 AOI21_X1 _40101_ (.A(_15450_),
    .B1(_12433_),
    .B2(_15451_),
    .ZN(_15452_));
 OAI22_X1 _40102_ (.A1(_15449_),
    .A2(_12811_),
    .B1(_15452_),
    .B2(_14362_),
    .ZN(_15453_));
 BUF_X4 _40103_ (.A(_15431_),
    .Z(_15454_));
 MUX2_X1 _40104_ (.A(\core.keymem.prev_key1_reg[101] ),
    .B(_15453_),
    .S(_15454_),
    .Z(_02887_));
 AOI21_X1 _40105_ (.A(_11886_),
    .B1(_11887_),
    .B2(_15451_),
    .ZN(_15455_));
 OAI22_X1 _40106_ (.A1(_15449_),
    .A2(_11902_),
    .B1(_15455_),
    .B2(_14362_),
    .ZN(_15456_));
 BUF_X4 _40107_ (.A(_15431_),
    .Z(_15457_));
 MUX2_X1 _40108_ (.A(\core.keymem.prev_key1_reg[102] ),
    .B(_15456_),
    .S(_15457_),
    .Z(_02888_));
 NAND2_X1 _40109_ (.A1(\core.keymem.prev_key1_reg[103] ),
    .A2(_15443_),
    .ZN(_15458_));
 OAI21_X1 _40110_ (.A(_15454_),
    .B1(_11913_),
    .B2(_06680_),
    .ZN(_15459_));
 OAI21_X1 _40111_ (.A(_15458_),
    .B1(_15459_),
    .B2(_11927_),
    .ZN(_02889_));
 NAND2_X1 _40112_ (.A1(\core.keymem.prev_key1_reg[104] ),
    .A2(_15443_),
    .ZN(_15460_));
 AOI21_X1 _40113_ (.A(_15172_),
    .B1(_12663_),
    .B2(_15451_),
    .ZN(_15461_));
 NOR2_X1 _40114_ (.A1(_14289_),
    .A2(_15461_),
    .ZN(_15462_));
 AOI21_X1 _40115_ (.A(_15462_),
    .B1(_12820_),
    .B2(_14439_),
    .ZN(_15463_));
 OAI21_X1 _40116_ (.A(_15460_),
    .B1(_15463_),
    .B2(_15448_),
    .ZN(_02890_));
 AOI21_X1 _40117_ (.A(_15175_),
    .B1(_12684_),
    .B2(_15451_),
    .ZN(_15464_));
 OAI22_X1 _40118_ (.A1(_15449_),
    .A2(_12828_),
    .B1(_15464_),
    .B2(_14362_),
    .ZN(_15465_));
 MUX2_X1 _40119_ (.A(\core.keymem.prev_key1_reg[105] ),
    .B(_15465_),
    .S(_15457_),
    .Z(_02891_));
 NAND2_X1 _40120_ (.A1(\core.keymem.prev_key1_reg[106] ),
    .A2(_15443_),
    .ZN(_15466_));
 OAI21_X1 _40121_ (.A(_15466_),
    .B1(_15448_),
    .B2(_11950_),
    .ZN(_02892_));
 NOR2_X1 _40122_ (.A1(_11965_),
    .A2(_11958_),
    .ZN(_15467_));
 MUX2_X1 _40123_ (.A(\core.keymem.prev_key1_reg[107] ),
    .B(_15467_),
    .S(_15457_),
    .Z(_02893_));
 NAND2_X1 _40124_ (.A1(\core.keymem.prev_key1_reg[108] ),
    .A2(_15443_),
    .ZN(_15468_));
 NAND2_X1 _40125_ (.A1(_14293_),
    .A2(_11979_),
    .ZN(_15469_));
 BUF_X4 _40126_ (.A(_15431_),
    .Z(_15470_));
 NAND2_X1 _40127_ (.A1(_15469_),
    .A2(_15470_),
    .ZN(_15471_));
 OAI21_X1 _40128_ (.A(_15468_),
    .B1(_15471_),
    .B2(_11976_),
    .ZN(_02894_));
 NOR2_X1 _40129_ (.A1(_14282_),
    .A2(_12840_),
    .ZN(_15472_));
 NOR2_X1 _40130_ (.A1(_15184_),
    .A2(_15472_),
    .ZN(_15473_));
 OAI21_X1 _40131_ (.A(_14404_),
    .B1(_14367_),
    .B2(\core.key[109] ),
    .ZN(_15474_));
 OAI22_X1 _40132_ (.A1(_14289_),
    .A2(_15473_),
    .B1(_15474_),
    .B2(_12838_),
    .ZN(_15475_));
 MUX2_X1 _40133_ (.A(\core.keymem.prev_key1_reg[109] ),
    .B(_15475_),
    .S(_15457_),
    .Z(_02895_));
 NAND2_X2 _40134_ (.A1(_12808_),
    .A2(_15430_),
    .ZN(_15476_));
 BUF_X4 _40135_ (.A(_15476_),
    .Z(_15477_));
 NOR2_X1 _40136_ (.A1(_14282_),
    .A2(_12855_),
    .ZN(_15478_));
 AOI22_X1 _40137_ (.A1(_11983_),
    .A2(_14242_),
    .B1(_15478_),
    .B2(\core.keymem.prev_key1_reg[10] ),
    .ZN(_15479_));
 AOI21_X1 _40138_ (.A(_15446_),
    .B1(_12855_),
    .B2(_14265_),
    .ZN(_15480_));
 OAI22_X1 _40139_ (.A1(_15477_),
    .A2(_15479_),
    .B1(_15480_),
    .B2(\core.keymem.prev_key1_reg[10] ),
    .ZN(_15481_));
 NOR2_X4 _40140_ (.A1(_12292_),
    .A2(_15441_),
    .ZN(_15482_));
 INV_X1 _40141_ (.A(_12851_),
    .ZN(_15483_));
 OAI21_X1 _40142_ (.A(_14226_),
    .B1(_12850_),
    .B2(_15483_),
    .ZN(_15484_));
 AOI21_X1 _40143_ (.A(_15481_),
    .B1(_15482_),
    .B2(_15484_),
    .ZN(_02896_));
 AOI21_X1 _40144_ (.A(_15188_),
    .B1(_12703_),
    .B2(_14313_),
    .ZN(_15485_));
 OAI21_X1 _40145_ (.A(_11998_),
    .B1(_15485_),
    .B2(_14289_),
    .ZN(_15486_));
 MUX2_X1 _40146_ (.A(_11999_),
    .B(_15486_),
    .S(_15457_),
    .Z(_02897_));
 NOR3_X1 _40147_ (.A1(_12015_),
    .A2(_12009_),
    .A3(_15442_),
    .ZN(_15487_));
 AOI21_X1 _40148_ (.A(_15487_),
    .B1(_15443_),
    .B2(\core.keymem.prev_key1_reg[111] ),
    .ZN(_15488_));
 INV_X1 _40149_ (.A(_15488_),
    .ZN(_02898_));
 AOI21_X1 _40150_ (.A(_12024_),
    .B1(_12026_),
    .B2(_14313_),
    .ZN(_15489_));
 BUF_X4 _40151_ (.A(_14274_),
    .Z(_15490_));
 OAI21_X1 _40152_ (.A(_12023_),
    .B1(_15489_),
    .B2(_15490_),
    .ZN(_15491_));
 MUX2_X1 _40153_ (.A(_12025_),
    .B(_15491_),
    .S(_15457_),
    .Z(_02899_));
 NAND2_X1 _40154_ (.A1(\core.keymem.prev_key1_reg[113] ),
    .A2(_15443_),
    .ZN(_15492_));
 AOI21_X1 _40155_ (.A(_15194_),
    .B1(_12865_),
    .B2(_15451_),
    .ZN(_15493_));
 NOR2_X1 _40156_ (.A1(_14289_),
    .A2(_15493_),
    .ZN(_15494_));
 AOI21_X1 _40157_ (.A(_15494_),
    .B1(_12864_),
    .B2(_14439_),
    .ZN(_15495_));
 OAI21_X1 _40158_ (.A(_15492_),
    .B1(_15495_),
    .B2(_15448_),
    .ZN(_02900_));
 MUX2_X1 _40159_ (.A(_00147_),
    .B(_12047_),
    .S(_12158_),
    .Z(_15496_));
 OAI22_X1 _40160_ (.A1(_15449_),
    .A2(_12045_),
    .B1(_15496_),
    .B2(_14362_),
    .ZN(_15497_));
 MUX2_X1 _40161_ (.A(\core.keymem.prev_key1_reg[114] ),
    .B(_15497_),
    .S(_15457_),
    .Z(_02901_));
 BUF_X4 _40162_ (.A(_15442_),
    .Z(_15498_));
 NAND2_X1 _40163_ (.A1(\core.keymem.prev_key1_reg[115] ),
    .A2(_15498_),
    .ZN(_15499_));
 NAND2_X1 _40164_ (.A1(_14293_),
    .A2(_12057_),
    .ZN(_15500_));
 NAND2_X1 _40165_ (.A1(_15500_),
    .A2(_15470_),
    .ZN(_15501_));
 OAI21_X1 _40166_ (.A(_15499_),
    .B1(_15501_),
    .B2(_12054_),
    .ZN(_02902_));
 NAND2_X1 _40167_ (.A1(\core.keymem.prev_key1_reg[116] ),
    .A2(_15498_),
    .ZN(_15502_));
 NAND2_X1 _40168_ (.A1(_14293_),
    .A2(_12075_),
    .ZN(_15503_));
 NAND2_X1 _40169_ (.A1(_15503_),
    .A2(_15470_),
    .ZN(_15504_));
 OAI21_X1 _40170_ (.A(_15502_),
    .B1(_15504_),
    .B2(_12071_),
    .ZN(_02903_));
 NAND2_X1 _40171_ (.A1(\core.keymem.prev_key1_reg[117] ),
    .A2(_15498_),
    .ZN(_15505_));
 AOI21_X1 _40172_ (.A(_15200_),
    .B1(_12578_),
    .B2(_15451_),
    .ZN(_15506_));
 NOR2_X1 _40173_ (.A1(_14289_),
    .A2(_15506_),
    .ZN(_15507_));
 AOI21_X1 _40174_ (.A(_15507_),
    .B1(_12873_),
    .B2(_14439_),
    .ZN(_15508_));
 BUF_X4 _40175_ (.A(_15447_),
    .Z(_15509_));
 OAI21_X1 _40176_ (.A(_15505_),
    .B1(_15508_),
    .B2(_15509_),
    .ZN(_02904_));
 AOI21_X1 _40177_ (.A(_15203_),
    .B1(_12728_),
    .B2(_15451_),
    .ZN(_15510_));
 OAI22_X1 _40178_ (.A1(_15449_),
    .A2(_12880_),
    .B1(_15510_),
    .B2(_14362_),
    .ZN(_15511_));
 MUX2_X1 _40179_ (.A(\core.keymem.prev_key1_reg[118] ),
    .B(_15511_),
    .S(_15457_),
    .Z(_02905_));
 NOR3_X1 _40180_ (.A1(_12094_),
    .A2(_12085_),
    .A3(_15442_),
    .ZN(_15512_));
 AOI21_X1 _40181_ (.A(_15512_),
    .B1(_15443_),
    .B2(\core.keymem.prev_key1_reg[119] ),
    .ZN(_15513_));
 INV_X1 _40182_ (.A(_15513_),
    .ZN(_02906_));
 NAND2_X4 _40183_ (.A1(_12148_),
    .A2(_15429_),
    .ZN(_15514_));
 AOI21_X1 _40184_ (.A(_15514_),
    .B1(_12893_),
    .B2(_14226_),
    .ZN(_15515_));
 NOR2_X1 _40185_ (.A1(_12860_),
    .A2(_12887_),
    .ZN(_15516_));
 AOI22_X1 _40186_ (.A1(_00406_),
    .A2(_14264_),
    .B1(_15516_),
    .B2(\core.keymem.prev_key1_reg[11] ),
    .ZN(_15517_));
 AOI21_X1 _40187_ (.A(_15446_),
    .B1(_12887_),
    .B2(_14265_),
    .ZN(_15518_));
 OAI22_X1 _40188_ (.A1(_15477_),
    .A2(_15517_),
    .B1(_15518_),
    .B2(\core.keymem.prev_key1_reg[11] ),
    .ZN(_15519_));
 NOR2_X1 _40189_ (.A1(_15515_),
    .A2(_15519_),
    .ZN(_02907_));
 MUX2_X1 _40190_ (.A(_00157_),
    .B(_12122_),
    .S(_12834_),
    .Z(_15520_));
 OAI21_X1 _40191_ (.A(_12120_),
    .B1(_15520_),
    .B2(_15490_),
    .ZN(_15521_));
 MUX2_X1 _40192_ (.A(\core.keymem.prev_key1_reg[120] ),
    .B(_15521_),
    .S(_15457_),
    .Z(_02908_));
 INV_X1 _40193_ (.A(_00160_),
    .ZN(_15522_));
 AOI21_X1 _40194_ (.A(_12147_),
    .B1(_14464_),
    .B2(_15522_),
    .ZN(_15523_));
 NOR2_X1 _40195_ (.A1(_00159_),
    .A2(_13331_),
    .ZN(_15524_));
 AOI21_X1 _40196_ (.A(_15524_),
    .B1(_12155_),
    .B2(_15451_),
    .ZN(_15525_));
 OAI22_X1 _40197_ (.A1(_15449_),
    .A2(_15523_),
    .B1(_15525_),
    .B2(_14362_),
    .ZN(_15526_));
 MUX2_X1 _40198_ (.A(\core.keymem.prev_key1_reg[121] ),
    .B(_15526_),
    .S(_15457_),
    .Z(_02909_));
 MUX2_X1 _40199_ (.A(_00161_),
    .B(_12901_),
    .S(_12158_),
    .Z(_15527_));
 BUF_X4 _40200_ (.A(_13132_),
    .Z(_15528_));
 OAI22_X1 _40201_ (.A1(_15449_),
    .A2(_12900_),
    .B1(_15527_),
    .B2(_15528_),
    .ZN(_15529_));
 BUF_X4 _40202_ (.A(_15431_),
    .Z(_15530_));
 MUX2_X1 _40203_ (.A(\core.keymem.prev_key1_reg[122] ),
    .B(_15529_),
    .S(_15530_),
    .Z(_02910_));
 MUX2_X1 _40204_ (.A(_00164_),
    .B(_12179_),
    .S(_12844_),
    .Z(_15531_));
 MUX2_X1 _40205_ (.A(_00163_),
    .B(_12168_),
    .S(_12158_),
    .Z(_15532_));
 OAI22_X1 _40206_ (.A1(_15449_),
    .A2(_15531_),
    .B1(_15532_),
    .B2(_15528_),
    .ZN(_15533_));
 MUX2_X1 _40207_ (.A(\core.keymem.prev_key1_reg[123] ),
    .B(_15533_),
    .S(_15530_),
    .Z(_02911_));
 AOI21_X1 _40208_ (.A(_13441_),
    .B1(_12186_),
    .B2(_12924_),
    .ZN(_15534_));
 AOI21_X1 _40209_ (.A(_14274_),
    .B1(_12907_),
    .B2(_12913_),
    .ZN(_15535_));
 NOR2_X1 _40210_ (.A1(_15534_),
    .A2(_15535_),
    .ZN(_15536_));
 MUX2_X1 _40211_ (.A(\core.keymem.prev_key1_reg[124] ),
    .B(_15536_),
    .S(_15530_),
    .Z(_02912_));
 AOI21_X1 _40212_ (.A(_12927_),
    .B1(_12306_),
    .B2(_14267_),
    .ZN(_15537_));
 MUX2_X1 _40213_ (.A(_12189_),
    .B(_12930_),
    .S(_12158_),
    .Z(_15538_));
 OAI22_X1 _40214_ (.A1(_15449_),
    .A2(_15537_),
    .B1(_15538_),
    .B2(_15528_),
    .ZN(_15539_));
 MUX2_X1 _40215_ (.A(\core.keymem.prev_key1_reg[125] ),
    .B(_15539_),
    .S(_15530_),
    .Z(_02913_));
 NOR2_X1 _40216_ (.A1(\core.keymem.prev_key1_reg[126] ),
    .A2(_15454_),
    .ZN(_15540_));
 BUF_X4 _40217_ (.A(_15446_),
    .Z(_15541_));
 NAND2_X1 _40218_ (.A1(_14248_),
    .A2(_12196_),
    .ZN(_15542_));
 AOI21_X1 _40219_ (.A(_14362_),
    .B1(_00169_),
    .B2(_14264_),
    .ZN(_15543_));
 AOI21_X1 _40220_ (.A(_15541_),
    .B1(_15542_),
    .B2(_15543_),
    .ZN(_15544_));
 OAI21_X1 _40221_ (.A(_14439_),
    .B1(_12205_),
    .B2(_12198_),
    .ZN(_15545_));
 AOI21_X1 _40222_ (.A(_15540_),
    .B1(_15544_),
    .B2(_15545_),
    .ZN(_02914_));
 MUX2_X1 _40223_ (.A(_00171_),
    .B(_12943_),
    .S(_12158_),
    .Z(_15546_));
 OAI22_X1 _40224_ (.A1(_15449_),
    .A2(_12941_),
    .B1(_15546_),
    .B2(_15528_),
    .ZN(_15547_));
 MUX2_X1 _40225_ (.A(\core.keymem.prev_key1_reg[127] ),
    .B(_15547_),
    .S(_15530_),
    .Z(_02915_));
 NOR2_X1 _40226_ (.A1(_14282_),
    .A2(_12503_),
    .ZN(_15548_));
 AOI22_X1 _40227_ (.A1(_00407_),
    .A2(_14242_),
    .B1(_15548_),
    .B2(_07313_),
    .ZN(_15549_));
 AOI21_X1 _40228_ (.A(_15446_),
    .B1(_12503_),
    .B2(_14265_),
    .ZN(_15550_));
 OAI22_X1 _40229_ (.A1(_15477_),
    .A2(_15549_),
    .B1(_15550_),
    .B2(_07313_),
    .ZN(_15551_));
 MUX2_X1 _40230_ (.A(\core.key[12] ),
    .B(_12955_),
    .S(_14267_),
    .Z(_15552_));
 NAND2_X1 _40231_ (.A1(_14226_),
    .A2(_15552_),
    .ZN(_15553_));
 AOI21_X1 _40232_ (.A(_15551_),
    .B1(_15553_),
    .B2(_15482_),
    .ZN(_02916_));
 NOR3_X1 _40233_ (.A1(_14238_),
    .A2(_12969_),
    .A3(_12967_),
    .ZN(_15554_));
 OAI21_X1 _40234_ (.A(\core.keymem.prev_key1_reg[13] ),
    .B1(_15541_),
    .B2(_15554_),
    .ZN(_15555_));
 AOI21_X1 _40235_ (.A(_12884_),
    .B1(_12969_),
    .B2(_14287_),
    .ZN(_15556_));
 OR2_X1 _40236_ (.A1(_12967_),
    .A2(_15556_),
    .ZN(_15557_));
 OAI21_X1 _40237_ (.A(_14238_),
    .B1(_00408_),
    .B2(_15490_),
    .ZN(_15558_));
 NAND2_X1 _40238_ (.A1(_15470_),
    .A2(_15558_),
    .ZN(_15559_));
 OAI21_X1 _40239_ (.A(_15555_),
    .B1(_15557_),
    .B2(_15559_),
    .ZN(_02917_));
 OAI21_X1 _40240_ (.A(_15482_),
    .B1(_12983_),
    .B2(_14264_),
    .ZN(_15560_));
 XNOR2_X1 _40241_ (.A(_12987_),
    .B(_12704_),
    .ZN(_15561_));
 AOI21_X1 _40242_ (.A(_15442_),
    .B1(_15561_),
    .B2(_14265_),
    .ZN(_15562_));
 OAI21_X1 _40243_ (.A(_15560_),
    .B1(_15562_),
    .B2(_07349_),
    .ZN(_15563_));
 NAND2_X1 _40244_ (.A1(_14248_),
    .A2(_12989_),
    .ZN(_15564_));
 OAI21_X1 _40245_ (.A(_14302_),
    .B1(_15564_),
    .B2(_07466_),
    .ZN(_15565_));
 INV_X1 _40246_ (.A(_15476_),
    .ZN(_15566_));
 AOI21_X1 _40247_ (.A(_15563_),
    .B1(_15565_),
    .B2(_15566_),
    .ZN(_02918_));
 NOR2_X1 _40248_ (.A1(_14205_),
    .A2(_12517_),
    .ZN(_15567_));
 AOI22_X1 _40249_ (.A1(_00410_),
    .A2(_14264_),
    .B1(_15567_),
    .B2(_07357_),
    .ZN(_15568_));
 AOI21_X1 _40250_ (.A(_15442_),
    .B1(_12517_),
    .B2(_14265_),
    .ZN(_15569_));
 OAI22_X1 _40251_ (.A1(_15477_),
    .A2(_15568_),
    .B1(_15569_),
    .B2(_07357_),
    .ZN(_15570_));
 AOI221_X1 _40252_ (.A(_15514_),
    .B1(_13010_),
    .B2(_13011_),
    .C1(\core.key[15] ),
    .C2(_12946_),
    .ZN(_15571_));
 NOR2_X1 _40253_ (.A1(_15570_),
    .A2(_15571_),
    .ZN(_02919_));
 AOI21_X1 _40254_ (.A(_06679_),
    .B1(_00411_),
    .B2(_14304_),
    .ZN(_15572_));
 NAND2_X1 _40255_ (.A1(_12526_),
    .A2(_12025_),
    .ZN(_15573_));
 NAND2_X1 _40256_ (.A1(_08253_),
    .A2(_12527_),
    .ZN(_15574_));
 OAI22_X1 _40257_ (.A1(_12025_),
    .A2(_13025_),
    .B1(_15573_),
    .B2(_15574_),
    .ZN(_15575_));
 NAND2_X1 _40258_ (.A1(_12186_),
    .A2(_15575_),
    .ZN(_15576_));
 NOR3_X1 _40259_ (.A1(_08253_),
    .A2(_12527_),
    .A3(_15573_),
    .ZN(_15577_));
 XNOR2_X1 _40260_ (.A(_12526_),
    .B(_12025_),
    .ZN(_15578_));
 NOR2_X1 _40261_ (.A1(_13024_),
    .A2(_15578_),
    .ZN(_15579_));
 MUX2_X1 _40262_ (.A(_15577_),
    .B(_15579_),
    .S(_10613_),
    .Z(_15580_));
 AOI21_X1 _40263_ (.A(_13023_),
    .B1(_12025_),
    .B2(_10613_),
    .ZN(_15581_));
 AOI21_X1 _40264_ (.A(_15581_),
    .B1(_12026_),
    .B2(_13023_),
    .ZN(_15582_));
 AOI21_X1 _40265_ (.A(_15580_),
    .B1(_15582_),
    .B2(_13024_),
    .ZN(_15583_));
 OAI221_X1 _40266_ (.A(_15572_),
    .B1(_15576_),
    .B2(_10613_),
    .C1(_15583_),
    .C2(_14238_),
    .ZN(_15584_));
 MUX2_X1 _40267_ (.A(\core.key[16] ),
    .B(_13021_),
    .S(_14367_),
    .Z(_15585_));
 AOI21_X1 _40268_ (.A(_15447_),
    .B1(_15585_),
    .B2(_12336_),
    .ZN(_15586_));
 AOI22_X1 _40269_ (.A1(_08253_),
    .A2(_15509_),
    .B1(_15584_),
    .B2(_15586_),
    .ZN(_02920_));
 AOI21_X1 _40270_ (.A(_13132_),
    .B1(_00434_),
    .B2(_14282_),
    .ZN(_15587_));
 OAI21_X1 _40271_ (.A(_15587_),
    .B1(_13040_),
    .B2(_14304_),
    .ZN(_15588_));
 AOI21_X1 _40272_ (.A(_15446_),
    .B1(_12269_),
    .B2(\core.key[17] ),
    .ZN(_15589_));
 NAND2_X1 _40273_ (.A1(_12311_),
    .A2(_13034_),
    .ZN(_15590_));
 AND3_X1 _40274_ (.A1(_15588_),
    .A2(_15589_),
    .A3(_15590_),
    .ZN(_15591_));
 BUF_X4 _40275_ (.A(_15447_),
    .Z(_15592_));
 INV_X1 _40276_ (.A(\core.keymem.prev_key1_reg[17] ),
    .ZN(_15593_));
 AOI21_X1 _40277_ (.A(_15591_),
    .B1(_15592_),
    .B2(_15593_),
    .ZN(_02921_));
 NAND2_X1 _40278_ (.A1(_13441_),
    .A2(_14316_),
    .ZN(_15594_));
 AOI21_X1 _40279_ (.A(_15594_),
    .B1(_13092_),
    .B2(_14245_),
    .ZN(_15595_));
 AOI21_X1 _40280_ (.A(_15433_),
    .B1(_13084_),
    .B2(_13085_),
    .ZN(_15596_));
 NOR3_X1 _40281_ (.A1(_15447_),
    .A2(_15595_),
    .A3(_15596_),
    .ZN(_15597_));
 AOI21_X1 _40282_ (.A(_15597_),
    .B1(_15592_),
    .B2(_13087_),
    .ZN(_02922_));
 NAND3_X1 _40283_ (.A1(\core.keymem.prev_key1_reg[19] ),
    .A2(_14447_),
    .A3(_13101_),
    .ZN(_15598_));
 AOI21_X1 _40284_ (.A(_12951_),
    .B1(_00436_),
    .B2(_12193_),
    .ZN(_15599_));
 NAND2_X1 _40285_ (.A1(\core.key[19] ),
    .A2(_13415_),
    .ZN(_15600_));
 OAI21_X1 _40286_ (.A(_15600_),
    .B1(_13106_),
    .B2(_14277_),
    .ZN(_15601_));
 AOI221_X2 _40287_ (.A(_15446_),
    .B1(_15598_),
    .B2(_15599_),
    .C1(_15601_),
    .C2(_14404_),
    .ZN(_15602_));
 OAI21_X1 _40288_ (.A(_15470_),
    .B1(_13101_),
    .B2(_12884_),
    .ZN(_15603_));
 INV_X1 _40289_ (.A(\core.keymem.prev_key1_reg[19] ),
    .ZN(_15604_));
 AOI21_X1 _40290_ (.A(_15602_),
    .B1(_15603_),
    .B2(_15604_),
    .ZN(_02923_));
 NAND2_X1 _40291_ (.A1(_13114_),
    .A2(_15454_),
    .ZN(_15605_));
 NAND2_X1 _40292_ (.A1(\core.keymem.prev_key1_reg[1] ),
    .A2(_15447_),
    .ZN(_15606_));
 AOI22_X1 _40293_ (.A1(_13131_),
    .A2(_15482_),
    .B1(_15605_),
    .B2(_15606_),
    .ZN(_02924_));
 NOR2_X1 _40294_ (.A1(_14205_),
    .A2(_12546_),
    .ZN(_15607_));
 AOI22_X1 _40295_ (.A1(_00437_),
    .A2(_14264_),
    .B1(_15607_),
    .B2(_08233_),
    .ZN(_15608_));
 AOI21_X1 _40296_ (.A(_15442_),
    .B1(_12546_),
    .B2(_14265_),
    .ZN(_15609_));
 OAI22_X1 _40297_ (.A1(_15477_),
    .A2(_15608_),
    .B1(_15609_),
    .B2(_08233_),
    .ZN(_15610_));
 NAND2_X1 _40298_ (.A1(_13139_),
    .A2(_15482_),
    .ZN(_15611_));
 NOR2_X1 _40299_ (.A1(_13138_),
    .A2(_15611_),
    .ZN(_15612_));
 NOR2_X1 _40300_ (.A1(_15610_),
    .A2(_15612_),
    .ZN(_02925_));
 NAND3_X1 _40301_ (.A1(\core.keymem.prev_key1_reg[21] ),
    .A2(_13875_),
    .A3(_12581_),
    .ZN(_15613_));
 NAND2_X1 _40302_ (.A1(_00438_),
    .A2(_14282_),
    .ZN(_15614_));
 AOI21_X1 _40303_ (.A(_15476_),
    .B1(_15613_),
    .B2(_15614_),
    .ZN(_15615_));
 OAI21_X1 _40304_ (.A(_15430_),
    .B1(_12581_),
    .B2(_12884_),
    .ZN(_15616_));
 INV_X1 _40305_ (.A(\core.keymem.prev_key1_reg[21] ),
    .ZN(_15617_));
 OR2_X1 _40306_ (.A1(_14304_),
    .A2(_13152_),
    .ZN(_15618_));
 AOI221_X1 _40307_ (.A(_15615_),
    .B1(_15616_),
    .B2(_15617_),
    .C1(_15618_),
    .C2(_15482_),
    .ZN(_02926_));
 XNOR2_X1 _40308_ (.A(_12738_),
    .B(_13173_),
    .ZN(_15619_));
 AOI221_X2 _40309_ (.A(_15514_),
    .B1(_15619_),
    .B2(_13011_),
    .C1(_12946_),
    .C2(\core.key[22] ),
    .ZN(_15620_));
 NAND2_X1 _40310_ (.A1(_12028_),
    .A2(_13572_),
    .ZN(_15621_));
 NAND2_X1 _40311_ (.A1(_15430_),
    .A2(_15621_),
    .ZN(_15622_));
 NAND2_X1 _40312_ (.A1(_08298_),
    .A2(_13875_),
    .ZN(_15623_));
 OAI22_X2 _40313_ (.A1(_12235_),
    .A2(_14313_),
    .B1(_13572_),
    .B2(_15623_),
    .ZN(_15624_));
 AOI221_X2 _40314_ (.A(_15620_),
    .B1(_15622_),
    .B2(_08299_),
    .C1(_15566_),
    .C2(_15624_),
    .ZN(_02927_));
 MUX2_X1 _40315_ (.A(\core.keymem.prev_key1_reg[23] ),
    .B(_13195_),
    .S(_15530_),
    .Z(_02928_));
 BUF_X4 _40316_ (.A(_15430_),
    .Z(_15625_));
 MUX2_X1 _40317_ (.A(_00017_),
    .B(_13208_),
    .S(_13875_),
    .Z(_15626_));
 OAI21_X1 _40318_ (.A(_15625_),
    .B1(_15626_),
    .B2(_15435_),
    .ZN(_15627_));
 OAI22_X1 _40319_ (.A1(_09318_),
    .A2(_15432_),
    .B1(_15627_),
    .B2(_13203_),
    .ZN(_15628_));
 INV_X1 _40320_ (.A(_15628_),
    .ZN(_02929_));
 NOR2_X1 _40321_ (.A1(\core.keymem.prev_key1_reg[25] ),
    .A2(_15454_),
    .ZN(_15629_));
 MUX2_X1 _40322_ (.A(_12274_),
    .B(_13217_),
    .S(_12871_),
    .Z(_15630_));
 AOI21_X1 _40323_ (.A(_15541_),
    .B1(_15630_),
    .B2(_14293_),
    .ZN(_15631_));
 OR3_X1 _40324_ (.A1(_15433_),
    .A2(_13231_),
    .A3(_13219_),
    .ZN(_15632_));
 AOI21_X1 _40325_ (.A(_15629_),
    .B1(_15631_),
    .B2(_15632_),
    .ZN(_02930_));
 NOR2_X1 _40326_ (.A1(_12277_),
    .A2(_12284_),
    .ZN(_15633_));
 OAI21_X1 _40327_ (.A(_13239_),
    .B1(_15633_),
    .B2(_15490_),
    .ZN(_15634_));
 MUX2_X1 _40328_ (.A(\core.keymem.prev_key1_reg[26] ),
    .B(_15634_),
    .S(_15530_),
    .Z(_02931_));
 MUX2_X1 _40329_ (.A(_00026_),
    .B(_13281_),
    .S(_12185_),
    .Z(_15635_));
 NOR2_X1 _40330_ (.A1(_06680_),
    .A2(_15635_),
    .ZN(_15636_));
 OAI21_X1 _40331_ (.A(_15432_),
    .B1(_15636_),
    .B2(_13276_),
    .ZN(_15637_));
 INV_X1 _40332_ (.A(\core.keymem.prev_key1_reg[27] ),
    .ZN(_15638_));
 OAI21_X1 _40333_ (.A(_15637_),
    .B1(_15440_),
    .B2(_15638_),
    .ZN(_02932_));
 NOR2_X1 _40334_ (.A1(_14205_),
    .A2(_13321_),
    .ZN(_15639_));
 OAI21_X1 _40335_ (.A(_13441_),
    .B1(_13316_),
    .B2(_15639_),
    .ZN(_15640_));
 NAND2_X1 _40336_ (.A1(_13315_),
    .A2(_15640_),
    .ZN(_15641_));
 MUX2_X1 _40337_ (.A(_09282_),
    .B(_15641_),
    .S(_15530_),
    .Z(_02933_));
 OAI21_X1 _40338_ (.A(_13326_),
    .B1(_13327_),
    .B2(_12241_),
    .ZN(_15642_));
 MUX2_X1 _40339_ (.A(\core.keymem.prev_key1_reg[29] ),
    .B(_15642_),
    .S(_15530_),
    .Z(_02934_));
 NAND2_X1 _40340_ (.A1(\core.keymem.prev_key1_reg[2] ),
    .A2(_15498_),
    .ZN(_15643_));
 OAI21_X1 _40341_ (.A(_15643_),
    .B1(_15448_),
    .B2(_13334_),
    .ZN(_02935_));
 MUX2_X1 _40342_ (.A(_00035_),
    .B(_13340_),
    .S(_12185_),
    .Z(_15644_));
 NOR2_X1 _40343_ (.A1(_15435_),
    .A2(_15644_),
    .ZN(_15645_));
 OAI21_X1 _40344_ (.A(_15432_),
    .B1(_15645_),
    .B2(_13377_),
    .ZN(_15646_));
 OAI21_X1 _40345_ (.A(_15646_),
    .B1(_15440_),
    .B2(_09358_),
    .ZN(_02936_));
 NOR2_X1 _40346_ (.A1(_00038_),
    .A2(_12262_),
    .ZN(_15647_));
 AOI21_X1 _40347_ (.A(_15647_),
    .B1(_13391_),
    .B2(_14313_),
    .ZN(_15648_));
 OAI21_X1 _40348_ (.A(_15625_),
    .B1(_15648_),
    .B2(_15435_),
    .ZN(_15649_));
 OAI22_X1 _40349_ (.A1(_09268_),
    .A2(_15432_),
    .B1(_15649_),
    .B2(_13386_),
    .ZN(_15650_));
 INV_X1 _40350_ (.A(_15650_),
    .ZN(_02937_));
 NOR2_X1 _40351_ (.A1(_14205_),
    .A2(_12352_),
    .ZN(_15651_));
 NOR2_X1 _40352_ (.A1(_15254_),
    .A2(_15651_),
    .ZN(_15652_));
 OAI21_X1 _40353_ (.A(_12346_),
    .B1(_15652_),
    .B2(_15490_),
    .ZN(_15653_));
 MUX2_X1 _40354_ (.A(\core.keymem.prev_key1_reg[32] ),
    .B(_15653_),
    .S(_15530_),
    .Z(_02938_));
 AOI21_X1 _40355_ (.A(_12357_),
    .B1(_12360_),
    .B2(_14313_),
    .ZN(_15654_));
 OAI21_X1 _40356_ (.A(_13400_),
    .B1(_15654_),
    .B2(_15490_),
    .ZN(_15655_));
 BUF_X4 _40357_ (.A(_15430_),
    .Z(_15656_));
 MUX2_X1 _40358_ (.A(\core.keymem.prev_key1_reg[33] ),
    .B(_15655_),
    .S(_15656_),
    .Z(_02939_));
 BUF_X4 _40359_ (.A(_14447_),
    .Z(_15657_));
 AOI21_X1 _40360_ (.A(_12363_),
    .B1(_12317_),
    .B2(_15657_),
    .ZN(_15658_));
 OAI22_X1 _40361_ (.A1(_12374_),
    .A2(_12366_),
    .B1(_15658_),
    .B2(_15528_),
    .ZN(_15659_));
 MUX2_X1 _40362_ (.A(\core.keymem.prev_key1_reg[34] ),
    .B(_15659_),
    .S(_15656_),
    .Z(_02940_));
 AOI21_X1 _40363_ (.A(_12408_),
    .B1(_12411_),
    .B2(_14222_),
    .ZN(_15660_));
 OAI21_X1 _40364_ (.A(_12407_),
    .B1(_15660_),
    .B2(_15490_),
    .ZN(_15661_));
 MUX2_X1 _40365_ (.A(\core.keymem.prev_key1_reg[35] ),
    .B(_15661_),
    .S(_15656_),
    .Z(_02941_));
 NAND2_X1 _40366_ (.A1(_12184_),
    .A2(_12417_),
    .ZN(_15662_));
 OAI21_X1 _40367_ (.A(_15662_),
    .B1(_12002_),
    .B2(_00045_),
    .ZN(_15663_));
 AOI221_X2 _40368_ (.A(_15446_),
    .B1(_15663_),
    .B2(_12972_),
    .C1(_14404_),
    .C2(_12421_),
    .ZN(_15664_));
 INV_X1 _40369_ (.A(\core.keymem.prev_key1_reg[36] ),
    .ZN(_15665_));
 AOI21_X1 _40370_ (.A(_15664_),
    .B1(_15592_),
    .B2(_15665_),
    .ZN(_02942_));
 AOI21_X1 _40371_ (.A(_12432_),
    .B1(_12436_),
    .B2(_14313_),
    .ZN(_15666_));
 NOR2_X1 _40372_ (.A1(_15435_),
    .A2(_15666_),
    .ZN(_15667_));
 OAI21_X1 _40373_ (.A(_15470_),
    .B1(_15667_),
    .B2(_12431_),
    .ZN(_15668_));
 INV_X1 _40374_ (.A(\core.keymem.prev_key1_reg[37] ),
    .ZN(_15669_));
 OAI21_X1 _40375_ (.A(_15668_),
    .B1(_15440_),
    .B2(_15669_),
    .ZN(_02943_));
 AOI21_X1 _40376_ (.A(_12463_),
    .B1(_12466_),
    .B2(_14222_),
    .ZN(_15670_));
 OAI21_X1 _40377_ (.A(_12462_),
    .B1(_15670_),
    .B2(_15490_),
    .ZN(_15671_));
 MUX2_X1 _40378_ (.A(\core.keymem.prev_key1_reg[38] ),
    .B(_15671_),
    .S(_15656_),
    .Z(_02944_));
 BUF_X4 _40379_ (.A(_12786_),
    .Z(_15672_));
 OAI21_X1 _40380_ (.A(_13433_),
    .B1(_14267_),
    .B2(\core.key[39] ),
    .ZN(_15673_));
 MUX2_X1 _40381_ (.A(_00048_),
    .B(_13412_),
    .S(_13720_),
    .Z(_15674_));
 OAI22_X1 _40382_ (.A1(_15672_),
    .A2(_15673_),
    .B1(_15674_),
    .B2(_15528_),
    .ZN(_15675_));
 MUX2_X1 _40383_ (.A(\core.keymem.prev_key1_reg[39] ),
    .B(_15675_),
    .S(_15656_),
    .Z(_02945_));
 OAI21_X1 _40384_ (.A(_14364_),
    .B1(_13445_),
    .B2(_14278_),
    .ZN(_15676_));
 AOI21_X1 _40385_ (.A(_15514_),
    .B1(_15676_),
    .B2(_14226_),
    .ZN(_15677_));
 NAND3_X1 _40386_ (.A1(\core.keymem.prev_key1_reg[3] ),
    .A2(_14245_),
    .A3(_12411_),
    .ZN(_15678_));
 AOI21_X1 _40387_ (.A(_15476_),
    .B1(_15678_),
    .B2(_13437_),
    .ZN(_15679_));
 OR2_X1 _40388_ (.A1(_12884_),
    .A2(_12411_),
    .ZN(_15680_));
 AOI21_X1 _40389_ (.A(\core.keymem.prev_key1_reg[3] ),
    .B1(_15625_),
    .B2(_15680_),
    .ZN(_15681_));
 NOR3_X1 _40390_ (.A1(_15677_),
    .A2(_15679_),
    .A3(_15681_),
    .ZN(_02946_));
 AOI21_X1 _40391_ (.A(_15274_),
    .B1(_13455_),
    .B2(_14222_),
    .ZN(_15682_));
 OAI21_X1 _40392_ (.A(_14404_),
    .B1(_14367_),
    .B2(\core.key[40] ),
    .ZN(_15683_));
 AND2_X1 _40393_ (.A1(_14367_),
    .A2(_13453_),
    .ZN(_15684_));
 OAI22_X1 _40394_ (.A1(_14289_),
    .A2(_15682_),
    .B1(_15683_),
    .B2(_15684_),
    .ZN(_15685_));
 MUX2_X1 _40395_ (.A(\core.keymem.prev_key1_reg[40] ),
    .B(_15685_),
    .S(_15656_),
    .Z(_02947_));
 AOI21_X1 _40396_ (.A(_13458_),
    .B1(_13460_),
    .B2(_15657_),
    .ZN(_15686_));
 OAI22_X1 _40397_ (.A1(_13465_),
    .A2(_13462_),
    .B1(_15686_),
    .B2(_15528_),
    .ZN(_15687_));
 MUX2_X1 _40398_ (.A(\core.keymem.prev_key1_reg[41] ),
    .B(_15687_),
    .S(_15656_),
    .Z(_02948_));
 NAND3_X1 _40399_ (.A1(_12336_),
    .A2(_13485_),
    .A3(_13486_),
    .ZN(_15688_));
 OAI21_X1 _40400_ (.A(_13441_),
    .B1(_15280_),
    .B2(_15478_),
    .ZN(_15689_));
 NAND2_X1 _40401_ (.A1(_15688_),
    .A2(_15689_),
    .ZN(_15690_));
 MUX2_X1 _40402_ (.A(\core.keymem.prev_key1_reg[42] ),
    .B(_15690_),
    .S(_15656_),
    .Z(_02949_));
 NOR3_X1 _40403_ (.A1(_06679_),
    .A2(_15283_),
    .A3(_15516_),
    .ZN(_15691_));
 AOI21_X1 _40404_ (.A(_13441_),
    .B1(_14313_),
    .B2(_13494_),
    .ZN(_15692_));
 NOR2_X1 _40405_ (.A1(_15691_),
    .A2(_15692_),
    .ZN(_15693_));
 MUX2_X1 _40406_ (.A(\core.keymem.prev_key1_reg[43] ),
    .B(_15693_),
    .S(_15656_),
    .Z(_02950_));
 NOR2_X1 _40407_ (.A1(_12500_),
    .A2(_15548_),
    .ZN(_15694_));
 NOR2_X1 _40408_ (.A1(_15435_),
    .A2(_15694_),
    .ZN(_15695_));
 OAI21_X1 _40409_ (.A(_15470_),
    .B1(_15695_),
    .B2(_12499_),
    .ZN(_15696_));
 INV_X1 _40410_ (.A(\core.keymem.prev_key1_reg[44] ),
    .ZN(_15697_));
 OAI21_X1 _40411_ (.A(_15696_),
    .B1(_15440_),
    .B2(_15697_),
    .ZN(_02951_));
 NAND2_X1 _40412_ (.A1(_13506_),
    .A2(_13507_),
    .ZN(_15698_));
 AOI21_X1 _40413_ (.A(_15288_),
    .B1(_12969_),
    .B2(_15657_),
    .ZN(_15699_));
 OAI22_X1 _40414_ (.A1(_15672_),
    .A2(_15698_),
    .B1(_15699_),
    .B2(_15528_),
    .ZN(_15700_));
 MUX2_X1 _40415_ (.A(\core.keymem.prev_key1_reg[45] ),
    .B(_15700_),
    .S(_15656_),
    .Z(_02952_));
 NOR2_X1 _40416_ (.A1(_14242_),
    .A2(_15561_),
    .ZN(_15701_));
 OAI21_X1 _40417_ (.A(_14293_),
    .B1(_15291_),
    .B2(_15701_),
    .ZN(_15702_));
 AOI21_X1 _40418_ (.A(_13513_),
    .B1(_13514_),
    .B2(_14267_),
    .ZN(_15703_));
 AOI21_X1 _40419_ (.A(_15447_),
    .B1(_15703_),
    .B2(_12336_),
    .ZN(_15704_));
 AOI22_X1 _40420_ (.A1(_12988_),
    .A2(_15509_),
    .B1(_15702_),
    .B2(_15704_),
    .ZN(_02953_));
 NOR2_X1 _40421_ (.A1(_15294_),
    .A2(_15567_),
    .ZN(_15705_));
 OAI21_X1 _40422_ (.A(_15625_),
    .B1(_15705_),
    .B2(_15435_),
    .ZN(_15706_));
 OAI22_X1 _40423_ (.A1(\core.keymem.prev_key1_reg[47] ),
    .A2(_15432_),
    .B1(_15706_),
    .B2(_12514_),
    .ZN(_15707_));
 INV_X1 _40424_ (.A(_15707_),
    .ZN(_02954_));
 NAND2_X2 _40425_ (.A1(_12336_),
    .A2(_15430_),
    .ZN(_15708_));
 INV_X1 _40426_ (.A(\core.key[48] ),
    .ZN(_15709_));
 MUX2_X1 _40427_ (.A(_15709_),
    .B(_12523_),
    .S(_12844_),
    .Z(_15710_));
 OR2_X1 _40428_ (.A1(_15708_),
    .A2(_15710_),
    .ZN(_15711_));
 NOR3_X1 _40429_ (.A1(_12526_),
    .A2(_14304_),
    .A3(_12528_),
    .ZN(_15712_));
 NOR2_X1 _40430_ (.A1(_12525_),
    .A2(_15712_),
    .ZN(_15713_));
 AOI21_X1 _40431_ (.A(_15447_),
    .B1(_12528_),
    .B2(_14265_),
    .ZN(_15714_));
 OAI221_X1 _40432_ (.A(_15711_),
    .B1(_15713_),
    .B2(_15477_),
    .C1(_15714_),
    .C2(_13023_),
    .ZN(_02955_));
 MUX2_X1 _40433_ (.A(_00058_),
    .B(_13526_),
    .S(_13331_),
    .Z(_15715_));
 OR2_X1 _40434_ (.A1(_14289_),
    .A2(_15715_),
    .ZN(_15716_));
 OAI21_X1 _40435_ (.A(_12335_),
    .B1(_14367_),
    .B2(\core.key[49] ),
    .ZN(_15717_));
 AOI21_X1 _40436_ (.A(_15717_),
    .B1(_13523_),
    .B2(_14267_),
    .ZN(_15718_));
 NOR2_X1 _40437_ (.A1(_15447_),
    .A2(_15718_),
    .ZN(_15719_));
 AOI22_X1 _40438_ (.A1(_13525_),
    .A2(_15509_),
    .B1(_15716_),
    .B2(_15719_),
    .ZN(_02956_));
 AOI21_X1 _40439_ (.A(_12972_),
    .B1(\core.key[4] ),
    .B2(_14277_),
    .ZN(_15720_));
 NOR2_X1 _40440_ (.A1(_14274_),
    .A2(_14395_),
    .ZN(_15721_));
 NOR2_X1 _40441_ (.A1(_15720_),
    .A2(_15721_),
    .ZN(_15722_));
 NOR2_X1 _40442_ (.A1(_15490_),
    .A2(_00375_),
    .ZN(_15723_));
 OAI221_X1 _40443_ (.A(_15454_),
    .B1(_15722_),
    .B2(_13537_),
    .C1(_14226_),
    .C2(_15723_),
    .ZN(_15724_));
 OAI21_X1 _40444_ (.A(_15724_),
    .B1(_15440_),
    .B2(_06776_),
    .ZN(_02957_));
 OAI21_X1 _40445_ (.A(_14404_),
    .B1(_14267_),
    .B2(\core.key[50] ),
    .ZN(_15725_));
 MUX2_X1 _40446_ (.A(_00059_),
    .B(_13091_),
    .S(_13720_),
    .Z(_15726_));
 OAI22_X1 _40447_ (.A1(_13554_),
    .A2(_15725_),
    .B1(_15726_),
    .B2(_15528_),
    .ZN(_15727_));
 BUF_X4 _40448_ (.A(_15430_),
    .Z(_15728_));
 MUX2_X1 _40449_ (.A(\core.keymem.prev_key1_reg[50] ),
    .B(_15727_),
    .S(_15728_),
    .Z(_02958_));
 AOI21_X1 _40450_ (.A(_13558_),
    .B1(_13101_),
    .B2(_15657_),
    .ZN(_15729_));
 OAI22_X1 _40451_ (.A1(_13562_),
    .A2(_13560_),
    .B1(_15729_),
    .B2(_15528_),
    .ZN(_15730_));
 MUX2_X1 _40452_ (.A(\core.keymem.prev_key1_reg[51] ),
    .B(_15730_),
    .S(_15728_),
    .Z(_02959_));
 INV_X1 _40453_ (.A(\core.key[52] ),
    .ZN(_15731_));
 AOI21_X1 _40454_ (.A(_12786_),
    .B1(_14464_),
    .B2(_15731_),
    .ZN(_15732_));
 OAI21_X1 _40455_ (.A(_15732_),
    .B1(_12566_),
    .B2(_14278_),
    .ZN(_15733_));
 OAI21_X1 _40456_ (.A(_14293_),
    .B1(_12542_),
    .B2(_15607_),
    .ZN(_15734_));
 NAND3_X1 _40457_ (.A1(_15454_),
    .A2(_15733_),
    .A3(_15734_),
    .ZN(_15735_));
 OR2_X1 _40458_ (.A1(\core.keymem.prev_key1_reg[52] ),
    .A2(_15625_),
    .ZN(_15736_));
 AND2_X1 _40459_ (.A1(_15735_),
    .A2(_15736_),
    .ZN(_02960_));
 AOI21_X1 _40460_ (.A(_12576_),
    .B1(_12581_),
    .B2(_14313_),
    .ZN(_15737_));
 NOR2_X1 _40461_ (.A1(_15435_),
    .A2(_15737_),
    .ZN(_15738_));
 OAI21_X1 _40462_ (.A(_15470_),
    .B1(_15738_),
    .B2(_12575_),
    .ZN(_15739_));
 INV_X1 _40463_ (.A(\core.keymem.prev_key1_reg[53] ),
    .ZN(_15740_));
 OAI21_X1 _40464_ (.A(_15739_),
    .B1(_15440_),
    .B2(_15740_),
    .ZN(_02961_));
 NAND2_X4 _40465_ (.A1(_12971_),
    .A2(_12680_),
    .ZN(_15741_));
 NOR2_X1 _40466_ (.A1(_00063_),
    .A2(_15741_),
    .ZN(_15742_));
 NOR4_X1 _40467_ (.A1(_13570_),
    .A2(_13573_),
    .A3(_15442_),
    .A4(_15742_),
    .ZN(_15743_));
 AOI21_X1 _40468_ (.A(_15743_),
    .B1(_15592_),
    .B2(_13166_),
    .ZN(_02962_));
 MUX2_X1 _40469_ (.A(_00064_),
    .B(_12266_),
    .S(_13720_),
    .Z(_15744_));
 BUF_X4 _40470_ (.A(_13132_),
    .Z(_15745_));
 OAI22_X1 _40471_ (.A1(_15672_),
    .A2(_13579_),
    .B1(_15744_),
    .B2(_15745_),
    .ZN(_15746_));
 MUX2_X1 _40472_ (.A(\core.keymem.prev_key1_reg[55] ),
    .B(_15746_),
    .S(_15728_),
    .Z(_02963_));
 AOI21_X1 _40473_ (.A(_13584_),
    .B1(_13586_),
    .B2(_14367_),
    .ZN(_15747_));
 OAI222_X2 _40474_ (.A1(_15433_),
    .A2(_15747_),
    .B1(_13582_),
    .B2(_12884_),
    .C1(_15741_),
    .C2(_00065_),
    .ZN(_15748_));
 MUX2_X1 _40475_ (.A(\core.keymem.prev_key1_reg[56] ),
    .B(_15748_),
    .S(_15728_),
    .Z(_02964_));
 MUX2_X1 _40476_ (.A(_00067_),
    .B(_13602_),
    .S(_13720_),
    .Z(_15749_));
 OAI22_X1 _40477_ (.A1(_15672_),
    .A2(_13601_),
    .B1(_15749_),
    .B2(_15745_),
    .ZN(_15750_));
 MUX2_X1 _40478_ (.A(\core.keymem.prev_key1_reg[57] ),
    .B(_15750_),
    .S(_15728_),
    .Z(_02965_));
 NAND2_X1 _40479_ (.A1(\core.keymem.prev_key1_reg[58] ),
    .A2(_15541_),
    .ZN(_15751_));
 MUX2_X1 _40480_ (.A(_00070_),
    .B(_13609_),
    .S(_14267_),
    .Z(_15752_));
 AOI21_X1 _40481_ (.A(_14419_),
    .B1(_13606_),
    .B2(_14248_),
    .ZN(_15753_));
 OAI221_X1 _40482_ (.A(_15751_),
    .B1(_15752_),
    .B2(_15708_),
    .C1(_15477_),
    .C2(_15753_),
    .ZN(_02966_));
 NAND2_X1 _40483_ (.A1(\core.keymem.prev_key1_reg[59] ),
    .A2(_15541_),
    .ZN(_15754_));
 NOR2_X1 _40484_ (.A1(_14242_),
    .A2(_13614_),
    .ZN(_15755_));
 NOR2_X1 _40485_ (.A1(_14423_),
    .A2(_15755_),
    .ZN(_15756_));
 MUX2_X1 _40486_ (.A(_00072_),
    .B(_13613_),
    .S(_14267_),
    .Z(_15757_));
 OAI221_X1 _40487_ (.A(_15754_),
    .B1(_15756_),
    .B2(_15477_),
    .C1(_15708_),
    .C2(_15757_),
    .ZN(_02967_));
 OAI21_X1 _40488_ (.A(_15324_),
    .B1(_12597_),
    .B2(_12193_),
    .ZN(_15758_));
 INV_X1 _40489_ (.A(\core.key[5] ),
    .ZN(_15759_));
 OAI21_X1 _40490_ (.A(_12604_),
    .B1(_12844_),
    .B2(_15759_),
    .ZN(_15760_));
 AOI221_X2 _40491_ (.A(_15446_),
    .B1(_15758_),
    .B2(_12972_),
    .C1(_14404_),
    .C2(_15760_),
    .ZN(_15761_));
 INV_X1 _40492_ (.A(\core.keymem.prev_key1_reg[5] ),
    .ZN(_15762_));
 AOI21_X1 _40493_ (.A(_15761_),
    .B1(_15592_),
    .B2(_15762_),
    .ZN(_02968_));
 OR3_X1 _40494_ (.A1(_00074_),
    .A2(_12844_),
    .A3(_12786_),
    .ZN(_15763_));
 MUX2_X1 _40495_ (.A(_00073_),
    .B(_13620_),
    .S(_14447_),
    .Z(_15764_));
 OAI221_X1 _40496_ (.A(_15763_),
    .B1(_13619_),
    .B2(_12241_),
    .C1(_15490_),
    .C2(_15764_),
    .ZN(_15765_));
 MUX2_X1 _40497_ (.A(\core.keymem.prev_key1_reg[60] ),
    .B(_15765_),
    .S(_15728_),
    .Z(_02969_));
 NOR3_X1 _40498_ (.A1(_11916_),
    .A2(_00076_),
    .A3(_12302_),
    .ZN(_15766_));
 AOI221_X1 _40499_ (.A(_15766_),
    .B1(_13623_),
    .B2(_12027_),
    .C1(_12808_),
    .C2(_15329_),
    .ZN(_15767_));
 XNOR2_X1 _40500_ (.A(_12306_),
    .B(_13628_),
    .ZN(_15768_));
 OAI21_X1 _40501_ (.A(_15767_),
    .B1(_15768_),
    .B2(_12241_),
    .ZN(_15769_));
 MUX2_X1 _40502_ (.A(\core.keymem.prev_key1_reg[61] ),
    .B(_15769_),
    .S(_15728_),
    .Z(_02970_));
 NAND2_X1 _40503_ (.A1(\core.keymem.prev_key1_reg[62] ),
    .A2(_15498_),
    .ZN(_15770_));
 OAI21_X1 _40504_ (.A(_13441_),
    .B1(_12610_),
    .B2(_12262_),
    .ZN(_15771_));
 AOI21_X1 _40505_ (.A(_15771_),
    .B1(_13635_),
    .B2(_14245_),
    .ZN(_15772_));
 AOI21_X1 _40506_ (.A(_15772_),
    .B1(_14438_),
    .B2(_14439_),
    .ZN(_15773_));
 OAI21_X1 _40507_ (.A(_15770_),
    .B1(_15773_),
    .B2(_15509_),
    .ZN(_02971_));
 MUX2_X1 _40508_ (.A(_00080_),
    .B(_13657_),
    .S(_12844_),
    .Z(_15774_));
 AOI21_X1 _40509_ (.A(_14441_),
    .B1(_13639_),
    .B2(_14245_),
    .ZN(_15775_));
 OAI221_X1 _40510_ (.A(_15625_),
    .B1(_15774_),
    .B2(_15433_),
    .C1(_15775_),
    .C2(_06680_),
    .ZN(_15776_));
 OR2_X1 _40511_ (.A1(\core.keymem.prev_key1_reg[63] ),
    .A2(_15625_),
    .ZN(_15777_));
 AND2_X1 _40512_ (.A1(_15776_),
    .A2(_15777_),
    .ZN(_02972_));
 OR3_X1 _40513_ (.A1(_13132_),
    .A2(_12614_),
    .A3(_12617_),
    .ZN(_15778_));
 OAI21_X1 _40514_ (.A(_15778_),
    .B1(_12620_),
    .B2(_15433_),
    .ZN(_15779_));
 MUX2_X1 _40515_ (.A(\core.keymem.prev_key1_reg[64] ),
    .B(_15779_),
    .S(_15728_),
    .Z(_02973_));
 OAI21_X1 _40516_ (.A(_13664_),
    .B1(_13670_),
    .B2(_15433_),
    .ZN(_15780_));
 MUX2_X1 _40517_ (.A(\core.keymem.prev_key1_reg[65] ),
    .B(_15780_),
    .S(_15728_),
    .Z(_02974_));
 NOR2_X1 _40518_ (.A1(_12860_),
    .A2(_12316_),
    .ZN(_15781_));
 OAI21_X1 _40519_ (.A(_13441_),
    .B1(_14448_),
    .B2(_15781_),
    .ZN(_15782_));
 NAND2_X1 _40520_ (.A1(_15431_),
    .A2(_15782_),
    .ZN(_15783_));
 MUX2_X1 _40521_ (.A(\core.key[66] ),
    .B(_13676_),
    .S(_14367_),
    .Z(_15784_));
 AOI21_X1 _40522_ (.A(_15783_),
    .B1(_15784_),
    .B2(_14439_),
    .ZN(_15785_));
 INV_X1 _40523_ (.A(\core.keymem.prev_key1_reg[66] ),
    .ZN(_15786_));
 AOI21_X1 _40524_ (.A(_15785_),
    .B1(_15592_),
    .B2(_15786_),
    .ZN(_02975_));
 NOR2_X1 _40525_ (.A1(_14205_),
    .A2(_12410_),
    .ZN(_15787_));
 NOR2_X1 _40526_ (.A1(_15345_),
    .A2(_15787_),
    .ZN(_15788_));
 NOR2_X1 _40527_ (.A1(_15435_),
    .A2(_15788_),
    .ZN(_15789_));
 OAI21_X1 _40528_ (.A(_15470_),
    .B1(_15789_),
    .B2(_13687_),
    .ZN(_15790_));
 INV_X1 _40529_ (.A(\core.keymem.prev_key1_reg[67] ),
    .ZN(_15791_));
 OAI21_X1 _40530_ (.A(_15790_),
    .B1(_15440_),
    .B2(_15791_),
    .ZN(_02976_));
 NOR2_X1 _40531_ (.A1(_12680_),
    .A2(_12416_),
    .ZN(_15792_));
 OR2_X1 _40532_ (.A1(_15348_),
    .A2(_15792_),
    .ZN(_15793_));
 OAI21_X1 _40533_ (.A(_12630_),
    .B1(_12632_),
    .B2(_13415_),
    .ZN(_15794_));
 AOI221_X1 _40534_ (.A(_15446_),
    .B1(_15793_),
    .B2(_12972_),
    .C1(_14404_),
    .C2(_15794_),
    .ZN(_15795_));
 INV_X1 _40535_ (.A(\core.keymem.prev_key1_reg[68] ),
    .ZN(_15796_));
 AOI21_X1 _40536_ (.A(_15795_),
    .B1(_15592_),
    .B2(_15796_),
    .ZN(_02977_));
 AOI21_X1 _40537_ (.A(_13697_),
    .B1(_14464_),
    .B2(\core.key[69] ),
    .ZN(_15797_));
 AOI21_X1 _40538_ (.A(_15351_),
    .B1(_13698_),
    .B2(_15657_),
    .ZN(_15798_));
 OAI22_X1 _40539_ (.A1(_15672_),
    .A2(_15797_),
    .B1(_15798_),
    .B2(_15745_),
    .ZN(_15799_));
 MUX2_X1 _40540_ (.A(_12434_),
    .B(_15799_),
    .S(_15728_),
    .Z(_02978_));
 NOR2_X1 _40541_ (.A1(_00378_),
    .A2(_15741_),
    .ZN(_15800_));
 NAND2_X1 _40542_ (.A1(_13703_),
    .A2(_13708_),
    .ZN(_15801_));
 OAI21_X2 _40543_ (.A(_15470_),
    .B1(_15800_),
    .B2(_15801_),
    .ZN(_15802_));
 OAI21_X1 _40544_ (.A(_15802_),
    .B1(_15440_),
    .B2(_06824_),
    .ZN(_02979_));
 AOI21_X1 _40545_ (.A(_13132_),
    .B1(_00087_),
    .B2(_14282_),
    .ZN(_15803_));
 OAI21_X1 _40546_ (.A(_15803_),
    .B1(_12643_),
    .B2(_14304_),
    .ZN(_15804_));
 AOI21_X1 _40547_ (.A(_12644_),
    .B1(_12646_),
    .B2(_14267_),
    .ZN(_15805_));
 OAI21_X1 _40548_ (.A(_15804_),
    .B1(_15805_),
    .B2(_15433_),
    .ZN(_15806_));
 MUX2_X1 _40549_ (.A(_12464_),
    .B(_15806_),
    .S(_15439_),
    .Z(_02980_));
 AOI21_X1 _40550_ (.A(_15357_),
    .B1(_12657_),
    .B2(_12871_),
    .ZN(_15807_));
 OAI21_X1 _40551_ (.A(_15431_),
    .B1(_15807_),
    .B2(_06679_),
    .ZN(_15808_));
 OAI21_X1 _40552_ (.A(_12651_),
    .B1(_12654_),
    .B2(_14278_),
    .ZN(_15809_));
 AOI21_X1 _40553_ (.A(_15808_),
    .B1(_15809_),
    .B2(_12336_),
    .ZN(_15810_));
 INV_X1 _40554_ (.A(\core.keymem.prev_key1_reg[71] ),
    .ZN(_15811_));
 AOI21_X1 _40555_ (.A(_15810_),
    .B1(_15592_),
    .B2(_15811_),
    .ZN(_02981_));
 NAND2_X1 _40556_ (.A1(_13331_),
    .A2(_12664_),
    .ZN(_15812_));
 AOI21_X1 _40557_ (.A(_12156_),
    .B1(_00089_),
    .B2(_12193_),
    .ZN(_15813_));
 MUX2_X1 _40558_ (.A(\core.key[72] ),
    .B(_12672_),
    .S(_12170_),
    .Z(_15814_));
 AOI221_X2 _40559_ (.A(_15441_),
    .B1(_15812_),
    .B2(_15813_),
    .C1(_15814_),
    .C2(_12335_),
    .ZN(_15815_));
 INV_X1 _40560_ (.A(\core.keymem.prev_key1_reg[72] ),
    .ZN(_15816_));
 AOI21_X1 _40561_ (.A(_15815_),
    .B1(_15592_),
    .B2(_15816_),
    .ZN(_02982_));
 NAND2_X1 _40562_ (.A1(_12683_),
    .A2(_15498_),
    .ZN(_15817_));
 NAND2_X1 _40563_ (.A1(_12347_),
    .A2(_12685_),
    .ZN(_15818_));
 AND3_X1 _40564_ (.A1(_12808_),
    .A2(_12681_),
    .A3(_15818_),
    .ZN(_15819_));
 AOI221_X1 _40565_ (.A(_15819_),
    .B1(_12679_),
    .B2(_12311_),
    .C1(\core.key[73] ),
    .C2(_12269_),
    .ZN(_15820_));
 OAI21_X1 _40566_ (.A(_15817_),
    .B1(_15820_),
    .B2(_15509_),
    .ZN(_02983_));
 NAND2_X1 _40567_ (.A1(\core.keymem.prev_key1_reg[74] ),
    .A2(_15498_),
    .ZN(_15821_));
 OAI21_X1 _40568_ (.A(_15821_),
    .B1(_15448_),
    .B2(_13725_),
    .ZN(_02984_));
 NOR2_X1 _40569_ (.A1(_12680_),
    .A2(_12886_),
    .ZN(_15822_));
 OR2_X1 _40570_ (.A1(_15366_),
    .A2(_15822_),
    .ZN(_15823_));
 AOI221_X2 _40571_ (.A(_15441_),
    .B1(_15823_),
    .B2(_12972_),
    .C1(_14404_),
    .C2(_13730_),
    .ZN(_15824_));
 INV_X1 _40572_ (.A(\core.keymem.prev_key1_reg[75] ),
    .ZN(_15825_));
 AOI21_X1 _40573_ (.A(_15824_),
    .B1(_15592_),
    .B2(_15825_),
    .ZN(_02985_));
 NAND2_X1 _40574_ (.A1(\core.keymem.prev_key1_reg[76] ),
    .A2(_15498_),
    .ZN(_15826_));
 OAI21_X1 _40575_ (.A(_13734_),
    .B1(_12502_),
    .B2(_14212_),
    .ZN(_15827_));
 NOR2_X1 _40576_ (.A1(_14289_),
    .A2(_15827_),
    .ZN(_15828_));
 OAI21_X1 _40577_ (.A(_13736_),
    .B1(_13739_),
    .B2(_14278_),
    .ZN(_15829_));
 AOI21_X1 _40578_ (.A(_15828_),
    .B1(_15829_),
    .B2(_14439_),
    .ZN(_15830_));
 OAI21_X1 _40579_ (.A(_15826_),
    .B1(_15830_),
    .B2(_15509_),
    .ZN(_02986_));
 AOI21_X1 _40580_ (.A(_13746_),
    .B1(_14464_),
    .B2(\core.key[77] ),
    .ZN(_15831_));
 AOI21_X1 _40581_ (.A(_13743_),
    .B1(_12968_),
    .B2(_15657_),
    .ZN(_15832_));
 OAI22_X1 _40582_ (.A1(_15672_),
    .A2(_15831_),
    .B1(_15832_),
    .B2(_15745_),
    .ZN(_15833_));
 MUX2_X1 _40583_ (.A(\core.keymem.prev_key1_reg[77] ),
    .B(_15833_),
    .S(_15439_),
    .Z(_02987_));
 NOR2_X1 _40584_ (.A1(_14277_),
    .A2(_12699_),
    .ZN(_15834_));
 AOI21_X1 _40585_ (.A(_15834_),
    .B1(_14464_),
    .B2(\core.key[78] ),
    .ZN(_15835_));
 AOI21_X1 _40586_ (.A(_15375_),
    .B1(_12704_),
    .B2(_15657_),
    .ZN(_15836_));
 OAI22_X1 _40587_ (.A1(_15672_),
    .A2(_15835_),
    .B1(_15836_),
    .B2(_15745_),
    .ZN(_15837_));
 MUX2_X1 _40588_ (.A(_12701_),
    .B(_15837_),
    .S(_15439_),
    .Z(_02988_));
 NOR2_X1 _40589_ (.A1(_14277_),
    .A2(_12512_),
    .ZN(_15838_));
 AOI21_X1 _40590_ (.A(_15838_),
    .B1(_14464_),
    .B2(\core.key[79] ),
    .ZN(_15839_));
 AOI21_X1 _40591_ (.A(_14475_),
    .B1(_12516_),
    .B2(_15657_),
    .ZN(_15840_));
 OAI22_X1 _40592_ (.A1(_15672_),
    .A2(_15839_),
    .B1(_15840_),
    .B2(_15745_),
    .ZN(_15841_));
 MUX2_X1 _40593_ (.A(\core.keymem.prev_key1_reg[79] ),
    .B(_15841_),
    .S(_15439_),
    .Z(_02989_));
 NAND2_X1 _40594_ (.A1(\core.keymem.prev_key1_reg[7] ),
    .A2(_15541_),
    .ZN(_15842_));
 MUX2_X1 _40595_ (.A(_00380_),
    .B(_13760_),
    .S(_14222_),
    .Z(_15843_));
 NAND2_X1 _40596_ (.A1(_14439_),
    .A2(_13765_),
    .ZN(_15844_));
 OAI221_X1 _40597_ (.A(_15842_),
    .B1(_15843_),
    .B2(_15477_),
    .C1(_15443_),
    .C2(_15844_),
    .ZN(_02990_));
 INV_X1 _40598_ (.A(_00097_),
    .ZN(_15845_));
 OAI21_X1 _40599_ (.A(_12972_),
    .B1(_15845_),
    .B2(_13875_),
    .ZN(_15846_));
 AOI21_X1 _40600_ (.A(_15846_),
    .B1(_12528_),
    .B2(_12186_),
    .ZN(_15847_));
 NOR3_X1 _40601_ (.A1(_12715_),
    .A2(_15447_),
    .A3(_15847_),
    .ZN(_15848_));
 AOI21_X1 _40602_ (.A(_15848_),
    .B1(_15448_),
    .B2(_15381_),
    .ZN(_02991_));
 NOR2_X1 _40603_ (.A1(_14282_),
    .A2(_13038_),
    .ZN(_15849_));
 NOR2_X1 _40604_ (.A1(_15384_),
    .A2(_15849_),
    .ZN(_15850_));
 OAI22_X1 _40605_ (.A1(_15672_),
    .A2(_13772_),
    .B1(_15850_),
    .B2(_15745_),
    .ZN(_15851_));
 MUX2_X1 _40606_ (.A(\core.keymem.prev_key1_reg[81] ),
    .B(_15851_),
    .S(_15439_),
    .Z(_02992_));
 NOR2_X1 _40607_ (.A1(_12860_),
    .A2(_13090_),
    .ZN(_15852_));
 NOR2_X1 _40608_ (.A1(_15387_),
    .A2(_15852_),
    .ZN(_15853_));
 OAI21_X1 _40609_ (.A(_15431_),
    .B1(_15853_),
    .B2(_06679_),
    .ZN(_15854_));
 OAI21_X1 _40610_ (.A(_13778_),
    .B1(_13780_),
    .B2(_14278_),
    .ZN(_15855_));
 AOI21_X1 _40611_ (.A(_15854_),
    .B1(_15855_),
    .B2(_12336_),
    .ZN(_15856_));
 INV_X1 _40612_ (.A(\core.keymem.prev_key1_reg[82] ),
    .ZN(_15857_));
 AOI21_X1 _40613_ (.A(_15856_),
    .B1(_15448_),
    .B2(_15857_),
    .ZN(_02993_));
 NOR2_X1 _40614_ (.A1(_12860_),
    .A2(_13100_),
    .ZN(_15858_));
 NOR2_X1 _40615_ (.A1(_13785_),
    .A2(_15858_),
    .ZN(_15859_));
 OAI21_X1 _40616_ (.A(_15431_),
    .B1(_15859_),
    .B2(_06679_),
    .ZN(_15860_));
 NAND2_X1 _40617_ (.A1(\core.key[83] ),
    .A2(_14464_),
    .ZN(_15861_));
 OAI21_X1 _40618_ (.A(_15861_),
    .B1(_13787_),
    .B2(_14278_),
    .ZN(_15862_));
 AOI21_X1 _40619_ (.A(_15860_),
    .B1(_15862_),
    .B2(_12336_),
    .ZN(_15863_));
 INV_X1 _40620_ (.A(\core.keymem.prev_key1_reg[83] ),
    .ZN(_15864_));
 AOI21_X1 _40621_ (.A(_15863_),
    .B1(_15448_),
    .B2(_15864_),
    .ZN(_02994_));
 NAND2_X1 _40622_ (.A1(\core.keymem.prev_key1_reg[84] ),
    .A2(_15498_),
    .ZN(_15865_));
 AOI21_X1 _40623_ (.A(_12721_),
    .B1(_12545_),
    .B2(_15451_),
    .ZN(_15866_));
 NOR2_X1 _40624_ (.A1(_14289_),
    .A2(_15866_),
    .ZN(_15867_));
 AOI21_X1 _40625_ (.A(_15867_),
    .B1(_12723_),
    .B2(_14439_),
    .ZN(_15868_));
 OAI21_X1 _40626_ (.A(_15865_),
    .B1(_15868_),
    .B2(_15509_),
    .ZN(_02995_));
 NOR2_X1 _40627_ (.A1(_14277_),
    .A2(_12573_),
    .ZN(_15869_));
 AOI21_X1 _40628_ (.A(_15869_),
    .B1(_14464_),
    .B2(\core.key[85] ),
    .ZN(_15870_));
 NOR2_X1 _40629_ (.A1(_12860_),
    .A2(_13795_),
    .ZN(_15871_));
 NOR2_X1 _40630_ (.A1(_13793_),
    .A2(_15871_),
    .ZN(_15872_));
 OAI22_X1 _40631_ (.A1(_15672_),
    .A2(_15870_),
    .B1(_15872_),
    .B2(_15745_),
    .ZN(_15873_));
 MUX2_X1 _40632_ (.A(_12579_),
    .B(_15873_),
    .S(_15439_),
    .Z(_02996_));
 NAND2_X1 _40633_ (.A1(\core.key[86] ),
    .A2(_14277_),
    .ZN(_15874_));
 AND2_X1 _40634_ (.A1(_12739_),
    .A2(_15874_),
    .ZN(_15875_));
 AOI21_X1 _40635_ (.A(_15396_),
    .B1(_12729_),
    .B2(_15657_),
    .ZN(_15876_));
 OAI22_X1 _40636_ (.A1(_15433_),
    .A2(_15875_),
    .B1(_15876_),
    .B2(_15745_),
    .ZN(_15877_));
 MUX2_X1 _40637_ (.A(_12727_),
    .B(_15877_),
    .S(_15439_),
    .Z(_02997_));
 AOI21_X1 _40638_ (.A(_14487_),
    .B1(_12265_),
    .B2(_15657_),
    .ZN(_15878_));
 OAI22_X1 _40639_ (.A1(_15433_),
    .A2(_13802_),
    .B1(_15878_),
    .B2(_15745_),
    .ZN(_15879_));
 MUX2_X1 _40640_ (.A(\core.keymem.prev_key1_reg[87] ),
    .B(_15879_),
    .S(_15439_),
    .Z(_02998_));
 NAND2_X1 _40641_ (.A1(_13204_),
    .A2(_15541_),
    .ZN(_15880_));
 NOR2_X1 _40642_ (.A1(_14242_),
    .A2(_13808_),
    .ZN(_15881_));
 NOR2_X1 _40643_ (.A1(_15401_),
    .A2(_15881_),
    .ZN(_15882_));
 OAI21_X1 _40644_ (.A(_13806_),
    .B1(_13201_),
    .B2(_14278_),
    .ZN(_15883_));
 OAI221_X1 _40645_ (.A(_15880_),
    .B1(_15882_),
    .B2(_15477_),
    .C1(_15883_),
    .C2(_15708_),
    .ZN(_02999_));
 OAI21_X1 _40646_ (.A(_15431_),
    .B1(_12155_),
    .B2(_14242_),
    .ZN(_15884_));
 AOI21_X1 _40647_ (.A(_13132_),
    .B1(_15403_),
    .B2(_12155_),
    .ZN(_15885_));
 OAI22_X1 _40648_ (.A1(_00107_),
    .A2(_15741_),
    .B1(_15885_),
    .B2(_14304_),
    .ZN(_15886_));
 AOI22_X1 _40649_ (.A1(_13213_),
    .A2(_15884_),
    .B1(_15886_),
    .B2(_15625_),
    .ZN(_15887_));
 OR2_X1 _40650_ (.A1(_13813_),
    .A2(_13814_),
    .ZN(_15888_));
 AOI21_X1 _40651_ (.A(_15887_),
    .B1(_15482_),
    .B2(_15888_),
    .ZN(_03000_));
 OAI21_X1 _40652_ (.A(_15625_),
    .B1(_13455_),
    .B2(_12884_),
    .ZN(_15889_));
 NAND2_X1 _40653_ (.A1(_07261_),
    .A2(_15889_),
    .ZN(_15890_));
 NAND3_X1 _40654_ (.A1(_12951_),
    .A2(\core.key[8] ),
    .A3(_12946_),
    .ZN(_15891_));
 OAI21_X1 _40655_ (.A(_15891_),
    .B1(_15405_),
    .B2(_06678_),
    .ZN(_15892_));
 AND2_X1 _40656_ (.A1(_13828_),
    .A2(_13835_),
    .ZN(_15893_));
 XNOR2_X1 _40657_ (.A(_12672_),
    .B(_15893_),
    .ZN(_15894_));
 NOR2_X1 _40658_ (.A1(_07261_),
    .A2(_12263_),
    .ZN(_15895_));
 AOI221_X1 _40659_ (.A(_15892_),
    .B1(_15894_),
    .B2(_12311_),
    .C1(_13455_),
    .C2(_15895_),
    .ZN(_15896_));
 OAI21_X1 _40660_ (.A(_15890_),
    .B1(_15896_),
    .B2(_15509_),
    .ZN(_03001_));
 NAND2_X1 _40661_ (.A1(_12279_),
    .A2(_15443_),
    .ZN(_15897_));
 OAI21_X1 _40662_ (.A(_14362_),
    .B1(_14242_),
    .B2(_13858_),
    .ZN(_15898_));
 NOR3_X1 _40663_ (.A1(_12279_),
    .A2(_11800_),
    .A3(_12901_),
    .ZN(_15899_));
 OR3_X1 _40664_ (.A1(_06679_),
    .A2(_15408_),
    .A3(_15899_),
    .ZN(_15900_));
 NAND3_X1 _40665_ (.A1(_15432_),
    .A2(_15898_),
    .A3(_15900_),
    .ZN(_15901_));
 NAND4_X1 _40666_ (.A1(_12279_),
    .A2(_14226_),
    .A3(_12901_),
    .A4(_15898_),
    .ZN(_15902_));
 NAND3_X1 _40667_ (.A1(_15897_),
    .A2(_15901_),
    .A3(_15902_),
    .ZN(_03002_));
 OAI21_X1 _40668_ (.A(_13865_),
    .B1(_13267_),
    .B2(_14464_),
    .ZN(_15903_));
 OAI21_X1 _40669_ (.A(_15435_),
    .B1(_14238_),
    .B2(_15903_),
    .ZN(_15904_));
 OR3_X1 _40670_ (.A1(_13277_),
    .A2(_12860_),
    .A3(_12168_),
    .ZN(_15905_));
 NOR2_X1 _40671_ (.A1(_06679_),
    .A2(_15411_),
    .ZN(_15906_));
 AOI21_X1 _40672_ (.A(_15442_),
    .B1(_15905_),
    .B2(_15906_),
    .ZN(_15907_));
 AND3_X1 _40673_ (.A1(_13277_),
    .A2(_12186_),
    .A3(_12168_),
    .ZN(_15908_));
 OAI21_X1 _40674_ (.A(_15904_),
    .B1(_15907_),
    .B2(_15908_),
    .ZN(_15909_));
 OAI21_X1 _40675_ (.A(_15909_),
    .B1(_15440_),
    .B2(_13862_),
    .ZN(_03003_));
 NOR2_X1 _40676_ (.A1(_13876_),
    .A2(_15454_),
    .ZN(_15910_));
 NAND3_X1 _40677_ (.A1(_14245_),
    .A2(_13872_),
    .A3(_13873_),
    .ZN(_15911_));
 NOR3_X1 _40678_ (.A1(_13317_),
    .A2(_12860_),
    .A3(_12912_),
    .ZN(_15912_));
 OAI21_X1 _40679_ (.A(_12972_),
    .B1(_00113_),
    .B2(_12185_),
    .ZN(_15913_));
 OAI21_X1 _40680_ (.A(_15430_),
    .B1(_15912_),
    .B2(_15913_),
    .ZN(_15914_));
 NAND3_X1 _40681_ (.A1(_13317_),
    .A2(_14313_),
    .A3(_12912_),
    .ZN(_15915_));
 AOI22_X1 _40682_ (.A1(_06680_),
    .A2(_15911_),
    .B1(_15914_),
    .B2(_15915_),
    .ZN(_15916_));
 OR2_X1 _40683_ (.A1(_15910_),
    .A2(_15916_),
    .ZN(_03004_));
 NOR2_X1 _40684_ (.A1(_00115_),
    .A2(_15741_),
    .ZN(_15917_));
 AOI21_X1 _40685_ (.A(_15917_),
    .B1(_13881_),
    .B2(_14265_),
    .ZN(_15918_));
 NAND2_X1 _40686_ (.A1(_12336_),
    .A2(_13883_),
    .ZN(_15919_));
 OAI21_X1 _40687_ (.A(_15918_),
    .B1(_15919_),
    .B2(_13887_),
    .ZN(_15920_));
 MUX2_X1 _40688_ (.A(_12294_),
    .B(_15920_),
    .S(_15439_),
    .Z(_03005_));
 NAND2_X1 _40689_ (.A1(_15451_),
    .A2(_13891_),
    .ZN(_15921_));
 OAI21_X1 _40690_ (.A(_14362_),
    .B1(_13890_),
    .B2(_15921_),
    .ZN(_15922_));
 NOR3_X1 _40691_ (.A1(_13336_),
    .A2(_11800_),
    .A3(_12196_),
    .ZN(_15923_));
 OR3_X1 _40692_ (.A1(_06679_),
    .A2(_15417_),
    .A3(_15923_),
    .ZN(_15924_));
 NAND3_X1 _40693_ (.A1(_15432_),
    .A2(_15922_),
    .A3(_15924_),
    .ZN(_15925_));
 AND2_X1 _40694_ (.A1(_14245_),
    .A2(_12196_),
    .ZN(_15926_));
 AOI21_X1 _40695_ (.A(_15541_),
    .B1(_15926_),
    .B2(_15922_),
    .ZN(_15927_));
 OAI21_X1 _40696_ (.A(_15925_),
    .B1(_15927_),
    .B2(_13893_),
    .ZN(_03006_));
 NAND2_X1 _40697_ (.A1(_12186_),
    .A2(_13898_),
    .ZN(_15928_));
 NOR2_X1 _40698_ (.A1(_13897_),
    .A2(_15928_),
    .ZN(_15929_));
 NOR3_X1 _40699_ (.A1(_13387_),
    .A2(_11800_),
    .A3(_12943_),
    .ZN(_15930_));
 NOR3_X1 _40700_ (.A1(_14274_),
    .A2(_15420_),
    .A3(_15930_),
    .ZN(_15931_));
 NOR2_X1 _40701_ (.A1(_15442_),
    .A2(_15931_),
    .ZN(_15932_));
 AND3_X1 _40702_ (.A1(_13387_),
    .A2(_14222_),
    .A3(_12943_),
    .ZN(_15933_));
 OAI22_X1 _40703_ (.A1(_14293_),
    .A2(_15929_),
    .B1(_15932_),
    .B2(_15933_),
    .ZN(_15934_));
 OAI21_X1 _40704_ (.A(_15934_),
    .B1(_15432_),
    .B2(_13900_),
    .ZN(_03007_));
 MUX2_X1 _40705_ (.A(_12758_),
    .B(_12351_),
    .S(_11875_),
    .Z(_15935_));
 AOI221_X1 _40706_ (.A(_15441_),
    .B1(_15935_),
    .B2(_12972_),
    .C1(_14404_),
    .C2(_13904_),
    .ZN(_15936_));
 AOI21_X1 _40707_ (.A(_15936_),
    .B1(_15448_),
    .B2(_12350_),
    .ZN(_03008_));
 NAND2_X1 _40708_ (.A1(\core.keymem.prev_key1_reg[97] ),
    .A2(_15498_),
    .ZN(_15937_));
 NAND2_X1 _40709_ (.A1(_12775_),
    .A2(_12764_),
    .ZN(_15938_));
 OAI21_X1 _40710_ (.A(_15937_),
    .B1(_15938_),
    .B2(_15509_),
    .ZN(_03009_));
 NAND2_X1 _40711_ (.A1(\core.keymem.prev_key1_reg[98] ),
    .A2(_15541_),
    .ZN(_15939_));
 AOI21_X1 _40712_ (.A(_12782_),
    .B1(_14238_),
    .B2(_00123_),
    .ZN(_15940_));
 OAI21_X1 _40713_ (.A(_15454_),
    .B1(_15940_),
    .B2(_06680_),
    .ZN(_15941_));
 AOI21_X1 _40714_ (.A(_14293_),
    .B1(_14226_),
    .B2(_12785_),
    .ZN(_15942_));
 OAI21_X1 _40715_ (.A(_15939_),
    .B1(_15941_),
    .B2(_15942_),
    .ZN(_03010_));
 NAND2_X1 _40716_ (.A1(\core.keymem.prev_key1_reg[99] ),
    .A2(_15541_),
    .ZN(_15943_));
 OAI21_X1 _40717_ (.A(_15454_),
    .B1(_12791_),
    .B2(_06680_),
    .ZN(_15944_));
 OAI21_X1 _40718_ (.A(_15943_),
    .B1(_15944_),
    .B2(_12798_),
    .ZN(_03011_));
 INV_X1 _40719_ (.A(\core.keymem.prev_key1_reg[9] ),
    .ZN(_15945_));
 NAND3_X1 _40720_ (.A1(_15945_),
    .A2(_14265_),
    .A3(_13460_),
    .ZN(_15946_));
 OR2_X1 _40721_ (.A1(_12786_),
    .A2(_13911_),
    .ZN(_15947_));
 NOR2_X1 _40722_ (.A1(_14277_),
    .A2(_13915_),
    .ZN(_15948_));
 OAI221_X1 _40723_ (.A(_15946_),
    .B1(_15947_),
    .B2(_15948_),
    .C1(_15741_),
    .C2(_00404_),
    .ZN(_15949_));
 OAI21_X1 _40724_ (.A(_15625_),
    .B1(_13460_),
    .B2(_12884_),
    .ZN(_15950_));
 AOI22_X1 _40725_ (.A1(_15432_),
    .A2(_15949_),
    .B1(_15950_),
    .B2(\core.keymem.prev_key1_reg[9] ),
    .ZN(_15951_));
 INV_X1 _40726_ (.A(_15951_),
    .ZN(_03012_));
 AOI21_X1 _40727_ (.A(_11798_),
    .B1(_11900_),
    .B2(_22104_),
    .ZN(_15952_));
 OR2_X2 _40728_ (.A1(_11916_),
    .A2(_15952_),
    .ZN(_15953_));
 BUF_X2 _40729_ (.A(_15953_),
    .Z(_15954_));
 OR2_X1 _40730_ (.A1(_11805_),
    .A2(_15954_),
    .ZN(_15955_));
 MUX2_X1 _40731_ (.A(_11952_),
    .B(_12937_),
    .S(_15954_),
    .Z(_15956_));
 OAI22_X1 _40732_ (.A1(_12106_),
    .A2(_15955_),
    .B1(_15956_),
    .B2(_16224_),
    .ZN(_15957_));
 INV_X1 _40733_ (.A(_15957_),
    .ZN(_03013_));
 XOR2_X1 _40734_ (.A(_12106_),
    .B(_12937_),
    .Z(_15958_));
 NAND3_X1 _40735_ (.A1(_11792_),
    .A2(_15954_),
    .A3(_15958_),
    .ZN(_15959_));
 NAND2_X1 _40736_ (.A1(_12751_),
    .A2(_12132_),
    .ZN(_15960_));
 OAI21_X1 _40737_ (.A(_15959_),
    .B1(_15960_),
    .B2(_15954_),
    .ZN(_03014_));
 MUX2_X1 _40738_ (.A(_11952_),
    .B(_12132_),
    .S(_15953_),
    .Z(_15961_));
 OAI22_X1 _40739_ (.A1(\core.keymem.rcon_reg[2] ),
    .A2(_15955_),
    .B1(_15961_),
    .B2(_16224_),
    .ZN(_15962_));
 INV_X1 _40740_ (.A(_15962_),
    .ZN(_03015_));
 XOR2_X1 _40741_ (.A(_12937_),
    .B(\core.keymem.rcon_reg[2] ),
    .Z(_15963_));
 MUX2_X1 _40742_ (.A(_11952_),
    .B(_15963_),
    .S(_15953_),
    .Z(_15964_));
 OAI22_X1 _40743_ (.A1(_12166_),
    .A2(_15955_),
    .B1(_15964_),
    .B2(_16224_),
    .ZN(_15965_));
 INV_X1 _40744_ (.A(_15965_),
    .ZN(_03016_));
 XOR2_X1 _40745_ (.A(_12937_),
    .B(_12166_),
    .Z(_15966_));
 NAND3_X1 _40746_ (.A1(_11792_),
    .A2(_15954_),
    .A3(_15966_),
    .ZN(_15967_));
 NAND2_X1 _40747_ (.A1(_12751_),
    .A2(_12908_),
    .ZN(_15968_));
 OAI21_X1 _40748_ (.A(_15967_),
    .B1(_15968_),
    .B2(_15954_),
    .ZN(_03017_));
 NAND3_X1 _40749_ (.A1(_11792_),
    .A2(_12908_),
    .A3(_15954_),
    .ZN(_15969_));
 NAND2_X1 _40750_ (.A1(_12751_),
    .A2(\core.keymem.rcon_logic.tmp_rcon[6] ),
    .ZN(_15970_));
 OAI21_X1 _40751_ (.A(_15969_),
    .B1(_15970_),
    .B2(_15954_),
    .ZN(_03018_));
 NAND3_X1 _40752_ (.A1(_11792_),
    .A2(\core.keymem.rcon_logic.tmp_rcon[6] ),
    .A3(_15954_),
    .ZN(_15971_));
 NAND2_X1 _40753_ (.A1(_12751_),
    .A2(_12194_),
    .ZN(_15972_));
 OAI21_X1 _40754_ (.A(_15971_),
    .B1(_15972_),
    .B2(_15954_),
    .ZN(_03019_));
 MUX2_X1 _40755_ (.A(_11952_),
    .B(_12194_),
    .S(_15953_),
    .Z(_15973_));
 OAI22_X1 _40756_ (.A1(_12937_),
    .A2(_15955_),
    .B1(_15973_),
    .B2(_16224_),
    .ZN(_15974_));
 INV_X1 _40757_ (.A(_15974_),
    .ZN(_03020_));
 AOI21_X1 _40758_ (.A(\core.keymem.key_mem_ctrl_reg[3] ),
    .B1(_16214_),
    .B2(\core.key_ready ),
    .ZN(_15975_));
 INV_X1 _40759_ (.A(_15975_),
    .ZN(_03021_));
 NOR2_X2 _40760_ (.A1(_16229_),
    .A2(\core.keymem.key_mem_ctrl_reg[2] ),
    .ZN(_15976_));
 NAND2_X1 _40761_ (.A1(_12917_),
    .A2(_15976_),
    .ZN(_15977_));
 NAND3_X1 _40762_ (.A1(_16286_),
    .A2(_12176_),
    .A3(_00326_),
    .ZN(_15978_));
 NAND2_X1 _40763_ (.A1(_15977_),
    .A2(_15978_),
    .ZN(_03022_));
 NAND2_X1 _40764_ (.A1(\core.keymem.round_ctr_reg[1] ),
    .A2(_15976_),
    .ZN(_15979_));
 NAND2_X1 _40765_ (.A1(_11792_),
    .A2(_00326_),
    .ZN(_15980_));
 OR2_X1 _40766_ (.A1(_15976_),
    .A2(_15980_),
    .ZN(_15981_));
 INV_X1 _40767_ (.A(_22107_),
    .ZN(_15982_));
 OAI21_X1 _40768_ (.A(_15979_),
    .B1(_15981_),
    .B2(_15982_),
    .ZN(_03023_));
 NOR2_X1 _40769_ (.A1(_13920_),
    .A2(_15980_),
    .ZN(_15983_));
 OAI21_X1 _40770_ (.A(_16218_),
    .B1(_15976_),
    .B2(_15983_),
    .ZN(_15984_));
 NAND2_X1 _40771_ (.A1(_12802_),
    .A2(_13920_),
    .ZN(_15985_));
 OAI21_X1 _40772_ (.A(_15984_),
    .B1(_15985_),
    .B2(_15981_),
    .ZN(_03024_));
 NAND2_X1 _40773_ (.A1(_11794_),
    .A2(_15976_),
    .ZN(_15986_));
 NAND3_X1 _40774_ (.A1(_16218_),
    .A2(_12917_),
    .A3(\core.keymem.round_ctr_reg[1] ),
    .ZN(_15987_));
 XNOR2_X1 _40775_ (.A(_00319_),
    .B(_15987_),
    .ZN(_15988_));
 OAI21_X1 _40776_ (.A(_15986_),
    .B1(_15988_),
    .B2(_15981_),
    .ZN(_03025_));
 OAI21_X1 _40777_ (.A(\core.aes_core_ctrl_reg[0] ),
    .B1(_16206_),
    .B2(_16210_),
    .ZN(_15989_));
 NAND2_X1 _40778_ (.A1(\core.ready ),
    .A2(_15989_),
    .ZN(_15990_));
 NAND2_X1 _40779_ (.A1(_16205_),
    .A2(_15990_),
    .ZN(_03026_));
 AOI22_X1 _40780_ (.A1(\core.aes_core_ctrl_reg[1] ),
    .A2(_16204_),
    .B1(_15989_),
    .B2(\core.result_valid ),
    .ZN(_15991_));
 INV_X1 _40781_ (.A(_15991_),
    .ZN(_03027_));
 BUF_X4 _40782_ (.A(_16203_),
    .Z(_15992_));
 BUF_X4 _40783_ (.A(_15992_),
    .Z(_15993_));
 NAND2_X4 _40784_ (.A1(_16335_),
    .A2(_16293_),
    .ZN(_15994_));
 OR3_X2 _40785_ (.A1(net6),
    .A2(net7),
    .A3(net5),
    .ZN(_15995_));
 NOR2_X4 _40786_ (.A1(net4),
    .A2(_15995_),
    .ZN(_15996_));
 NAND2_X2 _40787_ (.A1(_22100_),
    .A2(_15996_),
    .ZN(_15997_));
 NOR3_X4 _40788_ (.A1(_16297_),
    .A2(_15994_),
    .A3(_15997_),
    .ZN(_15998_));
 MUX2_X2 _40789_ (.A(_15993_),
    .B(_16289_),
    .S(_15998_),
    .Z(_03028_));
 INV_X2 _40790_ (.A(net4),
    .ZN(_15999_));
 AOI21_X2 _40791_ (.A(_22095_),
    .B1(_16294_),
    .B2(_22102_),
    .ZN(_16000_));
 NOR4_X4 _40792_ (.A1(_15999_),
    .A2(_16297_),
    .A3(_15995_),
    .A4(_16000_),
    .ZN(_16001_));
 NAND3_X4 _40793_ (.A1(_22094_),
    .A2(_16299_),
    .A3(_16001_),
    .ZN(_16002_));
 CLKBUF_X3 _40794_ (.A(_16002_),
    .Z(_16003_));
 MUX2_X1 _40795_ (.A(_16289_),
    .B(\core.key[224] ),
    .S(_16003_),
    .Z(_03029_));
 MUX2_X1 _40796_ (.A(_16302_),
    .B(\core.key[234] ),
    .S(_16003_),
    .Z(_03030_));
 MUX2_X1 _40797_ (.A(_16303_),
    .B(\core.key[235] ),
    .S(_16003_),
    .Z(_03031_));
 MUX2_X1 _40798_ (.A(_16304_),
    .B(\core.key[236] ),
    .S(_16003_),
    .Z(_03032_));
 MUX2_X1 _40799_ (.A(_16305_),
    .B(\core.key[237] ),
    .S(_16003_),
    .Z(_03033_));
 MUX2_X1 _40800_ (.A(_16306_),
    .B(\core.key[238] ),
    .S(_16003_),
    .Z(_03034_));
 MUX2_X1 _40801_ (.A(_16307_),
    .B(\core.key[239] ),
    .S(_16003_),
    .Z(_03035_));
 MUX2_X1 _40802_ (.A(_16308_),
    .B(\core.key[240] ),
    .S(_16003_),
    .Z(_03036_));
 MUX2_X1 _40803_ (.A(_16309_),
    .B(\core.key[241] ),
    .S(_16003_),
    .Z(_03037_));
 MUX2_X1 _40804_ (.A(_16310_),
    .B(\core.key[242] ),
    .S(_16003_),
    .Z(_03038_));
 BUF_X4 _40805_ (.A(_16002_),
    .Z(_16004_));
 MUX2_X1 _40806_ (.A(_16311_),
    .B(\core.key[243] ),
    .S(_16004_),
    .Z(_03039_));
 MUX2_X1 _40807_ (.A(_16313_),
    .B(\core.key[225] ),
    .S(_16004_),
    .Z(_03040_));
 MUX2_X1 _40808_ (.A(_16314_),
    .B(\core.key[244] ),
    .S(_16004_),
    .Z(_03041_));
 MUX2_X1 _40809_ (.A(_16315_),
    .B(\core.key[245] ),
    .S(_16004_),
    .Z(_03042_));
 MUX2_X1 _40810_ (.A(_16316_),
    .B(\core.key[246] ),
    .S(_16004_),
    .Z(_03043_));
 MUX2_X1 _40811_ (.A(_16317_),
    .B(\core.key[247] ),
    .S(_16004_),
    .Z(_03044_));
 MUX2_X1 _40812_ (.A(_16318_),
    .B(\core.key[248] ),
    .S(_16004_),
    .Z(_03045_));
 MUX2_X1 _40813_ (.A(_16319_),
    .B(\core.key[249] ),
    .S(_16004_),
    .Z(_03046_));
 MUX2_X1 _40814_ (.A(_16320_),
    .B(\core.key[250] ),
    .S(_16004_),
    .Z(_03047_));
 MUX2_X1 _40815_ (.A(_16321_),
    .B(\core.key[251] ),
    .S(_16004_),
    .Z(_03048_));
 BUF_X4 _40816_ (.A(_16002_),
    .Z(_16005_));
 MUX2_X1 _40817_ (.A(_16322_),
    .B(\core.key[252] ),
    .S(_16005_),
    .Z(_03049_));
 MUX2_X1 _40818_ (.A(_16324_),
    .B(\core.key[253] ),
    .S(_16005_),
    .Z(_03050_));
 MUX2_X1 _40819_ (.A(_16325_),
    .B(\core.key[226] ),
    .S(_16005_),
    .Z(_03051_));
 MUX2_X1 _40820_ (.A(_16326_),
    .B(\core.key[254] ),
    .S(_16005_),
    .Z(_03052_));
 MUX2_X1 _40821_ (.A(_16327_),
    .B(\core.key[255] ),
    .S(_16005_),
    .Z(_03053_));
 MUX2_X1 _40822_ (.A(_16328_),
    .B(\core.key[227] ),
    .S(_16005_),
    .Z(_03054_));
 MUX2_X1 _40823_ (.A(_16329_),
    .B(\core.key[228] ),
    .S(_16005_),
    .Z(_03055_));
 MUX2_X1 _40824_ (.A(_16330_),
    .B(\core.key[229] ),
    .S(_16005_),
    .Z(_03056_));
 MUX2_X1 _40825_ (.A(_16331_),
    .B(\core.key[230] ),
    .S(_16005_),
    .Z(_03057_));
 MUX2_X1 _40826_ (.A(_16332_),
    .B(\core.key[231] ),
    .S(_16005_),
    .Z(_03058_));
 MUX2_X1 _40827_ (.A(_16333_),
    .B(\core.key[232] ),
    .S(_16002_),
    .Z(_03059_));
 MUX2_X1 _40828_ (.A(_16334_),
    .B(\core.key[233] ),
    .S(_16002_),
    .Z(_03060_));
 NAND2_X4 _40829_ (.A1(_22094_),
    .A2(_16001_),
    .ZN(_16006_));
 NOR3_X4 _40830_ (.A1(_16335_),
    .A2(_16293_),
    .A3(_16006_),
    .ZN(_16007_));
 BUF_X4 _40831_ (.A(_16007_),
    .Z(_16008_));
 MUX2_X1 _40832_ (.A(\core.key[192] ),
    .B(_16289_),
    .S(_16008_),
    .Z(_03061_));
 MUX2_X1 _40833_ (.A(\core.key[202] ),
    .B(_16302_),
    .S(_16008_),
    .Z(_03062_));
 MUX2_X1 _40834_ (.A(\core.key[203] ),
    .B(_16303_),
    .S(_16008_),
    .Z(_03063_));
 MUX2_X1 _40835_ (.A(\core.key[204] ),
    .B(_16304_),
    .S(_16008_),
    .Z(_03064_));
 MUX2_X1 _40836_ (.A(\core.key[205] ),
    .B(_16305_),
    .S(_16008_),
    .Z(_03065_));
 MUX2_X1 _40837_ (.A(\core.key[206] ),
    .B(_16306_),
    .S(_16008_),
    .Z(_03066_));
 MUX2_X1 _40838_ (.A(\core.key[207] ),
    .B(_16307_),
    .S(_16008_),
    .Z(_03067_));
 MUX2_X1 _40839_ (.A(\core.key[208] ),
    .B(_16308_),
    .S(_16008_),
    .Z(_03068_));
 MUX2_X1 _40840_ (.A(\core.key[209] ),
    .B(_16309_),
    .S(_16008_),
    .Z(_03069_));
 MUX2_X1 _40841_ (.A(\core.key[210] ),
    .B(_16310_),
    .S(_16008_),
    .Z(_03070_));
 BUF_X4 _40842_ (.A(_16007_),
    .Z(_16009_));
 MUX2_X1 _40843_ (.A(\core.key[211] ),
    .B(_16311_),
    .S(_16009_),
    .Z(_03071_));
 MUX2_X1 _40844_ (.A(\core.key[193] ),
    .B(_16313_),
    .S(_16009_),
    .Z(_03072_));
 MUX2_X1 _40845_ (.A(\core.key[212] ),
    .B(_16314_),
    .S(_16009_),
    .Z(_03073_));
 MUX2_X1 _40846_ (.A(\core.key[213] ),
    .B(_16315_),
    .S(_16009_),
    .Z(_03074_));
 MUX2_X1 _40847_ (.A(\core.key[214] ),
    .B(_16316_),
    .S(_16009_),
    .Z(_03075_));
 MUX2_X1 _40848_ (.A(\core.key[215] ),
    .B(_16317_),
    .S(_16009_),
    .Z(_03076_));
 MUX2_X1 _40849_ (.A(\core.key[216] ),
    .B(_16318_),
    .S(_16009_),
    .Z(_03077_));
 MUX2_X1 _40850_ (.A(\core.key[217] ),
    .B(_16319_),
    .S(_16009_),
    .Z(_03078_));
 MUX2_X1 _40851_ (.A(\core.key[218] ),
    .B(_16320_),
    .S(_16009_),
    .Z(_03079_));
 MUX2_X1 _40852_ (.A(\core.key[219] ),
    .B(_16321_),
    .S(_16009_),
    .Z(_03080_));
 CLKBUF_X3 _40853_ (.A(_16007_),
    .Z(_16010_));
 MUX2_X1 _40854_ (.A(\core.key[220] ),
    .B(_16322_),
    .S(_16010_),
    .Z(_03081_));
 MUX2_X1 _40855_ (.A(\core.key[221] ),
    .B(_16324_),
    .S(_16010_),
    .Z(_03082_));
 MUX2_X1 _40856_ (.A(\core.key[194] ),
    .B(_16325_),
    .S(_16010_),
    .Z(_03083_));
 MUX2_X1 _40857_ (.A(\core.key[222] ),
    .B(_16326_),
    .S(_16010_),
    .Z(_03084_));
 MUX2_X1 _40858_ (.A(\core.key[223] ),
    .B(_16327_),
    .S(_16010_),
    .Z(_03085_));
 MUX2_X1 _40859_ (.A(\core.key[195] ),
    .B(_16328_),
    .S(_16010_),
    .Z(_03086_));
 MUX2_X1 _40860_ (.A(\core.key[196] ),
    .B(_16329_),
    .S(_16010_),
    .Z(_03087_));
 MUX2_X1 _40861_ (.A(\core.key[197] ),
    .B(_16330_),
    .S(_16010_),
    .Z(_03088_));
 MUX2_X1 _40862_ (.A(\core.key[198] ),
    .B(_16331_),
    .S(_16010_),
    .Z(_03089_));
 MUX2_X1 _40863_ (.A(\core.key[199] ),
    .B(_16332_),
    .S(_16010_),
    .Z(_03090_));
 MUX2_X1 _40864_ (.A(\core.key[200] ),
    .B(_16333_),
    .S(_16007_),
    .Z(_03091_));
 MUX2_X1 _40865_ (.A(\core.key[201] ),
    .B(_16334_),
    .S(_16007_),
    .Z(_03092_));
 NOR2_X4 _40866_ (.A1(_15994_),
    .A2(_16006_),
    .ZN(_16011_));
 BUF_X4 _40867_ (.A(_16011_),
    .Z(_16012_));
 MUX2_X1 _40868_ (.A(\core.key[160] ),
    .B(_16289_),
    .S(_16012_),
    .Z(_03093_));
 MUX2_X1 _40869_ (.A(\core.key[170] ),
    .B(_16302_),
    .S(_16012_),
    .Z(_03094_));
 MUX2_X1 _40870_ (.A(\core.key[171] ),
    .B(_16303_),
    .S(_16012_),
    .Z(_03095_));
 MUX2_X1 _40871_ (.A(\core.key[172] ),
    .B(_16304_),
    .S(_16012_),
    .Z(_03096_));
 MUX2_X1 _40872_ (.A(\core.key[173] ),
    .B(_16305_),
    .S(_16012_),
    .Z(_03097_));
 MUX2_X1 _40873_ (.A(\core.key[174] ),
    .B(_16306_),
    .S(_16012_),
    .Z(_03098_));
 MUX2_X1 _40874_ (.A(\core.key[175] ),
    .B(_16307_),
    .S(_16012_),
    .Z(_03099_));
 MUX2_X1 _40875_ (.A(\core.key[176] ),
    .B(_16308_),
    .S(_16012_),
    .Z(_03100_));
 MUX2_X1 _40876_ (.A(\core.key[177] ),
    .B(_16309_),
    .S(_16012_),
    .Z(_03101_));
 MUX2_X1 _40877_ (.A(\core.key[178] ),
    .B(_16310_),
    .S(_16012_),
    .Z(_03102_));
 BUF_X4 _40878_ (.A(_16011_),
    .Z(_16013_));
 MUX2_X1 _40879_ (.A(\core.key[179] ),
    .B(_16311_),
    .S(_16013_),
    .Z(_03103_));
 MUX2_X1 _40880_ (.A(\core.key[161] ),
    .B(_16313_),
    .S(_16013_),
    .Z(_03104_));
 MUX2_X1 _40881_ (.A(\core.key[180] ),
    .B(_16314_),
    .S(_16013_),
    .Z(_03105_));
 MUX2_X1 _40882_ (.A(\core.key[181] ),
    .B(_16315_),
    .S(_16013_),
    .Z(_03106_));
 MUX2_X1 _40883_ (.A(\core.key[182] ),
    .B(_16316_),
    .S(_16013_),
    .Z(_03107_));
 MUX2_X1 _40884_ (.A(\core.key[183] ),
    .B(_16317_),
    .S(_16013_),
    .Z(_03108_));
 MUX2_X1 _40885_ (.A(\core.key[184] ),
    .B(_16318_),
    .S(_16013_),
    .Z(_03109_));
 MUX2_X1 _40886_ (.A(\core.key[185] ),
    .B(_16319_),
    .S(_16013_),
    .Z(_03110_));
 MUX2_X1 _40887_ (.A(\core.key[186] ),
    .B(_16320_),
    .S(_16013_),
    .Z(_03111_));
 MUX2_X1 _40888_ (.A(\core.key[187] ),
    .B(_16321_),
    .S(_16013_),
    .Z(_03112_));
 BUF_X4 _40889_ (.A(_16011_),
    .Z(_16014_));
 MUX2_X1 _40890_ (.A(\core.key[188] ),
    .B(_16322_),
    .S(_16014_),
    .Z(_03113_));
 MUX2_X1 _40891_ (.A(\core.key[189] ),
    .B(_16324_),
    .S(_16014_),
    .Z(_03114_));
 MUX2_X1 _40892_ (.A(\core.key[162] ),
    .B(_16325_),
    .S(_16014_),
    .Z(_03115_));
 MUX2_X1 _40893_ (.A(\core.key[190] ),
    .B(_16326_),
    .S(_16014_),
    .Z(_03116_));
 MUX2_X1 _40894_ (.A(\core.key[191] ),
    .B(_16327_),
    .S(_16014_),
    .Z(_03117_));
 MUX2_X1 _40895_ (.A(\core.key[163] ),
    .B(_16328_),
    .S(_16014_),
    .Z(_03118_));
 MUX2_X1 _40896_ (.A(\core.key[164] ),
    .B(_16329_),
    .S(_16014_),
    .Z(_03119_));
 MUX2_X1 _40897_ (.A(\core.key[165] ),
    .B(_16330_),
    .S(_16014_),
    .Z(_03120_));
 MUX2_X1 _40898_ (.A(\core.key[166] ),
    .B(_16331_),
    .S(_16014_),
    .Z(_03121_));
 MUX2_X1 _40899_ (.A(\core.key[167] ),
    .B(_16332_),
    .S(_16014_),
    .Z(_03122_));
 MUX2_X1 _40900_ (.A(\core.key[168] ),
    .B(_16333_),
    .S(_16011_),
    .Z(_03123_));
 MUX2_X1 _40901_ (.A(\core.key[169] ),
    .B(_16334_),
    .S(_16011_),
    .Z(_03124_));
 NOR3_X4 _40902_ (.A1(_16291_),
    .A2(_16293_),
    .A3(_16006_),
    .ZN(_16015_));
 BUF_X4 _40903_ (.A(_16015_),
    .Z(_16016_));
 MUX2_X1 _40904_ (.A(\core.key[128] ),
    .B(_16289_),
    .S(_16016_),
    .Z(_03125_));
 MUX2_X1 _40905_ (.A(\core.key[138] ),
    .B(_16302_),
    .S(_16016_),
    .Z(_03126_));
 MUX2_X1 _40906_ (.A(\core.key[139] ),
    .B(_16303_),
    .S(_16016_),
    .Z(_03127_));
 MUX2_X1 _40907_ (.A(\core.key[140] ),
    .B(_16304_),
    .S(_16016_),
    .Z(_03128_));
 MUX2_X1 _40908_ (.A(\core.key[141] ),
    .B(_16305_),
    .S(_16016_),
    .Z(_03129_));
 MUX2_X1 _40909_ (.A(\core.key[142] ),
    .B(_16306_),
    .S(_16016_),
    .Z(_03130_));
 MUX2_X1 _40910_ (.A(\core.key[143] ),
    .B(_16307_),
    .S(_16016_),
    .Z(_03131_));
 MUX2_X1 _40911_ (.A(\core.key[144] ),
    .B(_16308_),
    .S(_16016_),
    .Z(_03132_));
 MUX2_X1 _40912_ (.A(\core.key[145] ),
    .B(_16309_),
    .S(_16016_),
    .Z(_03133_));
 MUX2_X1 _40913_ (.A(\core.key[146] ),
    .B(_16310_),
    .S(_16016_),
    .Z(_03134_));
 BUF_X4 _40914_ (.A(_16015_),
    .Z(_16017_));
 MUX2_X1 _40915_ (.A(\core.key[147] ),
    .B(_16311_),
    .S(_16017_),
    .Z(_03135_));
 MUX2_X1 _40916_ (.A(\core.key[129] ),
    .B(_16313_),
    .S(_16017_),
    .Z(_03136_));
 MUX2_X1 _40917_ (.A(\core.key[148] ),
    .B(_16314_),
    .S(_16017_),
    .Z(_03137_));
 MUX2_X1 _40918_ (.A(\core.key[149] ),
    .B(_16315_),
    .S(_16017_),
    .Z(_03138_));
 MUX2_X1 _40919_ (.A(\core.key[150] ),
    .B(_16316_),
    .S(_16017_),
    .Z(_03139_));
 MUX2_X1 _40920_ (.A(\core.key[151] ),
    .B(_16317_),
    .S(_16017_),
    .Z(_03140_));
 MUX2_X1 _40921_ (.A(\core.key[152] ),
    .B(_16318_),
    .S(_16017_),
    .Z(_03141_));
 MUX2_X1 _40922_ (.A(\core.key[153] ),
    .B(_16319_),
    .S(_16017_),
    .Z(_03142_));
 MUX2_X1 _40923_ (.A(\core.key[154] ),
    .B(_16320_),
    .S(_16017_),
    .Z(_03143_));
 MUX2_X1 _40924_ (.A(\core.key[155] ),
    .B(_16321_),
    .S(_16017_),
    .Z(_03144_));
 BUF_X4 _40925_ (.A(_16015_),
    .Z(_16018_));
 MUX2_X1 _40926_ (.A(\core.key[156] ),
    .B(_16322_),
    .S(_16018_),
    .Z(_03145_));
 MUX2_X1 _40927_ (.A(\core.key[157] ),
    .B(_16324_),
    .S(_16018_),
    .Z(_03146_));
 MUX2_X1 _40928_ (.A(\core.key[130] ),
    .B(_16325_),
    .S(_16018_),
    .Z(_03147_));
 MUX2_X1 _40929_ (.A(\core.key[158] ),
    .B(_16326_),
    .S(_16018_),
    .Z(_03148_));
 MUX2_X1 _40930_ (.A(\core.key[159] ),
    .B(_16327_),
    .S(_16018_),
    .Z(_03149_));
 MUX2_X1 _40931_ (.A(\core.key[131] ),
    .B(_16328_),
    .S(_16018_),
    .Z(_03150_));
 MUX2_X1 _40932_ (.A(\core.key[132] ),
    .B(_16329_),
    .S(_16018_),
    .Z(_03151_));
 MUX2_X1 _40933_ (.A(\core.key[133] ),
    .B(_16330_),
    .S(_16018_),
    .Z(_03152_));
 MUX2_X1 _40934_ (.A(\core.key[134] ),
    .B(_16331_),
    .S(_16018_),
    .Z(_03153_));
 MUX2_X1 _40935_ (.A(\core.key[135] ),
    .B(_16332_),
    .S(_16018_),
    .Z(_03154_));
 MUX2_X1 _40936_ (.A(\core.key[136] ),
    .B(_16333_),
    .S(_16015_),
    .Z(_03155_));
 MUX2_X1 _40937_ (.A(\core.key[137] ),
    .B(_16334_),
    .S(_16015_),
    .Z(_03156_));
 AND2_X1 _40938_ (.A1(net2),
    .A2(_16001_),
    .ZN(_16019_));
 BUF_X4 _40939_ (.A(_16019_),
    .Z(_16020_));
 NAND2_X4 _40940_ (.A1(_16299_),
    .A2(_16020_),
    .ZN(_16021_));
 BUF_X4 _40941_ (.A(_16021_),
    .Z(_16022_));
 MUX2_X1 _40942_ (.A(net18),
    .B(\core.key[96] ),
    .S(_16022_),
    .Z(_03157_));
 MUX2_X1 _40943_ (.A(_16302_),
    .B(\core.key[106] ),
    .S(_16022_),
    .Z(_03158_));
 MUX2_X1 _40944_ (.A(_16303_),
    .B(\core.key[107] ),
    .S(_16022_),
    .Z(_03159_));
 MUX2_X1 _40945_ (.A(_16304_),
    .B(\core.key[108] ),
    .S(_16022_),
    .Z(_03160_));
 MUX2_X1 _40946_ (.A(_16305_),
    .B(\core.key[109] ),
    .S(_16022_),
    .Z(_03161_));
 MUX2_X1 _40947_ (.A(_16306_),
    .B(\core.key[110] ),
    .S(_16022_),
    .Z(_03162_));
 MUX2_X1 _40948_ (.A(_16307_),
    .B(\core.key[111] ),
    .S(_16022_),
    .Z(_03163_));
 MUX2_X1 _40949_ (.A(_16308_),
    .B(\core.key[112] ),
    .S(_16022_),
    .Z(_03164_));
 MUX2_X1 _40950_ (.A(_16309_),
    .B(\core.key[113] ),
    .S(_16022_),
    .Z(_03165_));
 MUX2_X1 _40951_ (.A(_16310_),
    .B(\core.key[114] ),
    .S(_16022_),
    .Z(_03166_));
 BUF_X4 _40952_ (.A(_16021_),
    .Z(_16023_));
 MUX2_X1 _40953_ (.A(_16311_),
    .B(\core.key[115] ),
    .S(_16023_),
    .Z(_03167_));
 MUX2_X1 _40954_ (.A(net29),
    .B(\core.key[97] ),
    .S(_16023_),
    .Z(_03168_));
 MUX2_X1 _40955_ (.A(_16314_),
    .B(\core.key[116] ),
    .S(_16023_),
    .Z(_03169_));
 MUX2_X1 _40956_ (.A(_16315_),
    .B(\core.key[117] ),
    .S(_16023_),
    .Z(_03170_));
 MUX2_X1 _40957_ (.A(_16316_),
    .B(\core.key[118] ),
    .S(_16023_),
    .Z(_03171_));
 MUX2_X1 _40958_ (.A(_16317_),
    .B(\core.key[119] ),
    .S(_16023_),
    .Z(_03172_));
 MUX2_X1 _40959_ (.A(_16318_),
    .B(\core.key[120] ),
    .S(_16023_),
    .Z(_03173_));
 MUX2_X1 _40960_ (.A(_16319_),
    .B(\core.key[121] ),
    .S(_16023_),
    .Z(_03174_));
 MUX2_X1 _40961_ (.A(_16320_),
    .B(\core.key[122] ),
    .S(_16023_),
    .Z(_03175_));
 MUX2_X1 _40962_ (.A(_16321_),
    .B(\core.key[123] ),
    .S(_16023_),
    .Z(_03176_));
 CLKBUF_X3 _40963_ (.A(_16021_),
    .Z(_16024_));
 MUX2_X1 _40964_ (.A(_16322_),
    .B(\core.key[124] ),
    .S(_16024_),
    .Z(_03177_));
 MUX2_X1 _40965_ (.A(_16324_),
    .B(\core.key[125] ),
    .S(_16024_),
    .Z(_03178_));
 MUX2_X1 _40966_ (.A(_16325_),
    .B(\core.key[98] ),
    .S(_16024_),
    .Z(_03179_));
 MUX2_X1 _40967_ (.A(_16326_),
    .B(\core.key[126] ),
    .S(_16024_),
    .Z(_03180_));
 MUX2_X1 _40968_ (.A(_16327_),
    .B(\core.key[127] ),
    .S(_16024_),
    .Z(_03181_));
 MUX2_X1 _40969_ (.A(_16328_),
    .B(\core.key[99] ),
    .S(_16024_),
    .Z(_03182_));
 MUX2_X1 _40970_ (.A(_16329_),
    .B(\core.key[100] ),
    .S(_16024_),
    .Z(_03183_));
 MUX2_X1 _40971_ (.A(_16330_),
    .B(\core.key[101] ),
    .S(_16024_),
    .Z(_03184_));
 MUX2_X1 _40972_ (.A(_16331_),
    .B(\core.key[102] ),
    .S(_16024_),
    .Z(_03185_));
 MUX2_X1 _40973_ (.A(_16332_),
    .B(\core.key[103] ),
    .S(_16024_),
    .Z(_03186_));
 MUX2_X1 _40974_ (.A(_16333_),
    .B(\core.key[104] ),
    .S(_16021_),
    .Z(_03187_));
 MUX2_X1 _40975_ (.A(_16334_),
    .B(\core.key[105] ),
    .S(_16021_),
    .Z(_03188_));
 NAND2_X4 _40976_ (.A1(_16336_),
    .A2(_16020_),
    .ZN(_16025_));
 BUF_X4 _40977_ (.A(_16025_),
    .Z(_16026_));
 MUX2_X1 _40978_ (.A(net18),
    .B(\core.key[64] ),
    .S(_16026_),
    .Z(_03189_));
 MUX2_X1 _40979_ (.A(_16302_),
    .B(\core.key[74] ),
    .S(_16026_),
    .Z(_03190_));
 MUX2_X1 _40980_ (.A(_16303_),
    .B(\core.key[75] ),
    .S(_16026_),
    .Z(_03191_));
 MUX2_X1 _40981_ (.A(_16304_),
    .B(\core.key[76] ),
    .S(_16026_),
    .Z(_03192_));
 MUX2_X1 _40982_ (.A(_16305_),
    .B(\core.key[77] ),
    .S(_16026_),
    .Z(_03193_));
 MUX2_X1 _40983_ (.A(_16306_),
    .B(\core.key[78] ),
    .S(_16026_),
    .Z(_03194_));
 MUX2_X1 _40984_ (.A(_16307_),
    .B(\core.key[79] ),
    .S(_16026_),
    .Z(_03195_));
 MUX2_X1 _40985_ (.A(_16308_),
    .B(\core.key[80] ),
    .S(_16026_),
    .Z(_03196_));
 MUX2_X1 _40986_ (.A(_16309_),
    .B(\core.key[81] ),
    .S(_16026_),
    .Z(_03197_));
 MUX2_X1 _40987_ (.A(_16310_),
    .B(\core.key[82] ),
    .S(_16026_),
    .Z(_03198_));
 BUF_X4 _40988_ (.A(_16025_),
    .Z(_16027_));
 MUX2_X1 _40989_ (.A(_16311_),
    .B(\core.key[83] ),
    .S(_16027_),
    .Z(_03199_));
 MUX2_X1 _40990_ (.A(net29),
    .B(\core.key[65] ),
    .S(_16027_),
    .Z(_03200_));
 MUX2_X1 _40991_ (.A(_16314_),
    .B(\core.key[84] ),
    .S(_16027_),
    .Z(_03201_));
 MUX2_X1 _40992_ (.A(_16315_),
    .B(\core.key[85] ),
    .S(_16027_),
    .Z(_03202_));
 MUX2_X1 _40993_ (.A(_16316_),
    .B(\core.key[86] ),
    .S(_16027_),
    .Z(_03203_));
 MUX2_X1 _40994_ (.A(_16317_),
    .B(\core.key[87] ),
    .S(_16027_),
    .Z(_03204_));
 MUX2_X1 _40995_ (.A(_16318_),
    .B(\core.key[88] ),
    .S(_16027_),
    .Z(_03205_));
 MUX2_X1 _40996_ (.A(_16319_),
    .B(\core.key[89] ),
    .S(_16027_),
    .Z(_03206_));
 MUX2_X1 _40997_ (.A(_16320_),
    .B(\core.key[90] ),
    .S(_16027_),
    .Z(_03207_));
 MUX2_X1 _40998_ (.A(_16321_),
    .B(\core.key[91] ),
    .S(_16027_),
    .Z(_03208_));
 CLKBUF_X3 _40999_ (.A(_16025_),
    .Z(_16028_));
 MUX2_X1 _41000_ (.A(_16322_),
    .B(\core.key[92] ),
    .S(_16028_),
    .Z(_03209_));
 MUX2_X1 _41001_ (.A(_16324_),
    .B(\core.key[93] ),
    .S(_16028_),
    .Z(_03210_));
 MUX2_X1 _41002_ (.A(_16325_),
    .B(\core.key[66] ),
    .S(_16028_),
    .Z(_03211_));
 MUX2_X1 _41003_ (.A(_16326_),
    .B(\core.key[94] ),
    .S(_16028_),
    .Z(_03212_));
 MUX2_X1 _41004_ (.A(_16327_),
    .B(\core.key[95] ),
    .S(_16028_),
    .Z(_03213_));
 MUX2_X1 _41005_ (.A(_16328_),
    .B(\core.key[67] ),
    .S(_16028_),
    .Z(_03214_));
 MUX2_X1 _41006_ (.A(_16329_),
    .B(\core.key[68] ),
    .S(_16028_),
    .Z(_03215_));
 MUX2_X1 _41007_ (.A(_16330_),
    .B(\core.key[69] ),
    .S(_16028_),
    .Z(_03216_));
 MUX2_X1 _41008_ (.A(_16331_),
    .B(\core.key[70] ),
    .S(_16028_),
    .Z(_03217_));
 MUX2_X1 _41009_ (.A(_16332_),
    .B(\core.key[71] ),
    .S(_16028_),
    .Z(_03218_));
 MUX2_X1 _41010_ (.A(_16333_),
    .B(\core.key[72] ),
    .S(_16025_),
    .Z(_03219_));
 MUX2_X1 _41011_ (.A(_16334_),
    .B(\core.key[73] ),
    .S(_16025_),
    .Z(_03220_));
 NAND2_X4 _41012_ (.A1(_16342_),
    .A2(_16020_),
    .ZN(_16029_));
 BUF_X4 _41013_ (.A(_16029_),
    .Z(_16030_));
 MUX2_X1 _41014_ (.A(net18),
    .B(\core.key[32] ),
    .S(_16030_),
    .Z(_03221_));
 MUX2_X1 _41015_ (.A(net19),
    .B(\core.key[42] ),
    .S(_16030_),
    .Z(_03222_));
 MUX2_X1 _41016_ (.A(net20),
    .B(\core.key[43] ),
    .S(_16030_),
    .Z(_03223_));
 MUX2_X1 _41017_ (.A(net21),
    .B(\core.key[44] ),
    .S(_16030_),
    .Z(_03224_));
 MUX2_X1 _41018_ (.A(net22),
    .B(\core.key[45] ),
    .S(_16030_),
    .Z(_03225_));
 MUX2_X1 _41019_ (.A(net23),
    .B(\core.key[46] ),
    .S(_16030_),
    .Z(_03226_));
 MUX2_X1 _41020_ (.A(net24),
    .B(\core.key[47] ),
    .S(_16030_),
    .Z(_03227_));
 MUX2_X1 _41021_ (.A(net25),
    .B(\core.key[48] ),
    .S(_16030_),
    .Z(_03228_));
 MUX2_X1 _41022_ (.A(net26),
    .B(\core.key[49] ),
    .S(_16030_),
    .Z(_03229_));
 MUX2_X1 _41023_ (.A(net27),
    .B(\core.key[50] ),
    .S(_16030_),
    .Z(_03230_));
 BUF_X4 _41024_ (.A(_16029_),
    .Z(_16031_));
 MUX2_X1 _41025_ (.A(net28),
    .B(\core.key[51] ),
    .S(_16031_),
    .Z(_03231_));
 MUX2_X1 _41026_ (.A(net29),
    .B(\core.key[33] ),
    .S(_16031_),
    .Z(_03232_));
 MUX2_X1 _41027_ (.A(net30),
    .B(\core.key[52] ),
    .S(_16031_),
    .Z(_03233_));
 MUX2_X1 _41028_ (.A(net31),
    .B(\core.key[53] ),
    .S(_16031_),
    .Z(_03234_));
 MUX2_X1 _41029_ (.A(net32),
    .B(\core.key[54] ),
    .S(_16031_),
    .Z(_03235_));
 MUX2_X1 _41030_ (.A(net33),
    .B(\core.key[55] ),
    .S(_16031_),
    .Z(_03236_));
 MUX2_X1 _41031_ (.A(net34),
    .B(\core.key[56] ),
    .S(_16031_),
    .Z(_03237_));
 MUX2_X1 _41032_ (.A(net35),
    .B(\core.key[57] ),
    .S(_16031_),
    .Z(_03238_));
 MUX2_X1 _41033_ (.A(net36),
    .B(\core.key[58] ),
    .S(_16031_),
    .Z(_03239_));
 MUX2_X1 _41034_ (.A(net37),
    .B(\core.key[59] ),
    .S(_16031_),
    .Z(_03240_));
 BUF_X4 _41035_ (.A(_16029_),
    .Z(_16032_));
 MUX2_X1 _41036_ (.A(net38),
    .B(\core.key[60] ),
    .S(_16032_),
    .Z(_03241_));
 MUX2_X1 _41037_ (.A(net39),
    .B(\core.key[61] ),
    .S(_16032_),
    .Z(_03242_));
 MUX2_X1 _41038_ (.A(net40),
    .B(\core.key[34] ),
    .S(_16032_),
    .Z(_03243_));
 MUX2_X1 _41039_ (.A(net41),
    .B(\core.key[62] ),
    .S(_16032_),
    .Z(_03244_));
 MUX2_X1 _41040_ (.A(net42),
    .B(\core.key[63] ),
    .S(_16032_),
    .Z(_03245_));
 MUX2_X1 _41041_ (.A(net43),
    .B(\core.key[35] ),
    .S(_16032_),
    .Z(_03246_));
 MUX2_X1 _41042_ (.A(net44),
    .B(\core.key[36] ),
    .S(_16032_),
    .Z(_03247_));
 MUX2_X1 _41043_ (.A(net45),
    .B(\core.key[37] ),
    .S(_16032_),
    .Z(_03248_));
 MUX2_X1 _41044_ (.A(net46),
    .B(\core.key[38] ),
    .S(_16032_),
    .Z(_03249_));
 MUX2_X1 _41045_ (.A(net47),
    .B(\core.key[39] ),
    .S(_16032_),
    .Z(_03250_));
 MUX2_X1 _41046_ (.A(net48),
    .B(\core.key[40] ),
    .S(_16029_),
    .Z(_03251_));
 MUX2_X1 _41047_ (.A(net49),
    .B(\core.key[41] ),
    .S(_16029_),
    .Z(_03252_));
 NAND2_X4 _41048_ (.A1(_16294_),
    .A2(_16020_),
    .ZN(_16033_));
 BUF_X4 _41049_ (.A(_16033_),
    .Z(_16034_));
 MUX2_X1 _41050_ (.A(net18),
    .B(\core.key[0] ),
    .S(_16034_),
    .Z(_03253_));
 MUX2_X1 _41051_ (.A(net19),
    .B(\core.key[10] ),
    .S(_16034_),
    .Z(_03254_));
 MUX2_X1 _41052_ (.A(net20),
    .B(\core.key[11] ),
    .S(_16034_),
    .Z(_03255_));
 MUX2_X1 _41053_ (.A(net21),
    .B(\core.key[12] ),
    .S(_16034_),
    .Z(_03256_));
 MUX2_X1 _41054_ (.A(net22),
    .B(\core.key[13] ),
    .S(_16034_),
    .Z(_03257_));
 MUX2_X1 _41055_ (.A(net23),
    .B(\core.key[14] ),
    .S(_16034_),
    .Z(_03258_));
 MUX2_X1 _41056_ (.A(net24),
    .B(\core.key[15] ),
    .S(_16034_),
    .Z(_03259_));
 MUX2_X1 _41057_ (.A(net25),
    .B(\core.key[16] ),
    .S(_16034_),
    .Z(_03260_));
 MUX2_X1 _41058_ (.A(net26),
    .B(\core.key[17] ),
    .S(_16034_),
    .Z(_03261_));
 MUX2_X1 _41059_ (.A(net27),
    .B(\core.key[18] ),
    .S(_16034_),
    .Z(_03262_));
 BUF_X4 _41060_ (.A(_16033_),
    .Z(_16035_));
 MUX2_X1 _41061_ (.A(net28),
    .B(\core.key[19] ),
    .S(_16035_),
    .Z(_03263_));
 MUX2_X1 _41062_ (.A(net29),
    .B(\core.key[1] ),
    .S(_16035_),
    .Z(_03264_));
 MUX2_X1 _41063_ (.A(net30),
    .B(\core.key[20] ),
    .S(_16035_),
    .Z(_03265_));
 MUX2_X1 _41064_ (.A(net31),
    .B(\core.key[21] ),
    .S(_16035_),
    .Z(_03266_));
 MUX2_X1 _41065_ (.A(net32),
    .B(\core.key[22] ),
    .S(_16035_),
    .Z(_03267_));
 MUX2_X1 _41066_ (.A(net33),
    .B(\core.key[23] ),
    .S(_16035_),
    .Z(_03268_));
 MUX2_X1 _41067_ (.A(net34),
    .B(\core.key[24] ),
    .S(_16035_),
    .Z(_03269_));
 MUX2_X1 _41068_ (.A(net35),
    .B(\core.key[25] ),
    .S(_16035_),
    .Z(_03270_));
 MUX2_X1 _41069_ (.A(net36),
    .B(\core.key[26] ),
    .S(_16035_),
    .Z(_03271_));
 MUX2_X1 _41070_ (.A(net37),
    .B(\core.key[27] ),
    .S(_16035_),
    .Z(_03272_));
 BUF_X4 _41071_ (.A(_16033_),
    .Z(_16036_));
 MUX2_X1 _41072_ (.A(net38),
    .B(\core.key[28] ),
    .S(_16036_),
    .Z(_03273_));
 MUX2_X1 _41073_ (.A(net39),
    .B(\core.key[29] ),
    .S(_16036_),
    .Z(_03274_));
 MUX2_X1 _41074_ (.A(net40),
    .B(\core.key[2] ),
    .S(_16036_),
    .Z(_03275_));
 MUX2_X1 _41075_ (.A(net41),
    .B(\core.key[30] ),
    .S(_16036_),
    .Z(_03276_));
 MUX2_X1 _41076_ (.A(net42),
    .B(\core.key[31] ),
    .S(_16036_),
    .Z(_03277_));
 MUX2_X1 _41077_ (.A(net43),
    .B(\core.key[3] ),
    .S(_16036_),
    .Z(_03278_));
 MUX2_X1 _41078_ (.A(net44),
    .B(\core.key[4] ),
    .S(_16036_),
    .Z(_03279_));
 MUX2_X1 _41079_ (.A(net45),
    .B(\core.key[5] ),
    .S(_16036_),
    .Z(_03280_));
 MUX2_X1 _41080_ (.A(net46),
    .B(\core.key[6] ),
    .S(_16036_),
    .Z(_03281_));
 MUX2_X1 _41081_ (.A(net47),
    .B(\core.key[7] ),
    .S(_16036_),
    .Z(_03282_));
 MUX2_X1 _41082_ (.A(net48),
    .B(\core.key[8] ),
    .S(_16033_),
    .Z(_03283_));
 MUX2_X1 _41083_ (.A(net49),
    .B(\core.key[9] ),
    .S(_16033_),
    .Z(_03284_));
 MUX2_X1 _41084_ (.A(_06680_),
    .B(_16313_),
    .S(_15998_),
    .Z(_03285_));
 MUX2_X1 _41085_ (.A(\core.dec_block.block_w3_reg[0] ),
    .B(\core.enc_block.block_w3_reg[0] ),
    .S(_15993_),
    .Z(\core.muxed_new_block[0] ));
 MUX2_X1 _41086_ (.A(\core.dec_block.block_w0_reg[4] ),
    .B(_10368_),
    .S(_15993_),
    .Z(\core.muxed_new_block[100] ));
 MUX2_X1 _41087_ (.A(\core.dec_block.block_w0_reg[5] ),
    .B(_10425_),
    .S(_15993_),
    .Z(\core.muxed_new_block[101] ));
 MUX2_X1 _41088_ (.A(\core.dec_block.block_w0_reg[6] ),
    .B(_10482_),
    .S(_15993_),
    .Z(\core.muxed_new_block[102] ));
 MUX2_X1 _41089_ (.A(_16581_),
    .B(_10537_),
    .S(_15993_),
    .Z(\core.muxed_new_block[103] ));
 MUX2_X1 _41090_ (.A(\core.dec_block.block_w0_reg[8] ),
    .B(_10624_),
    .S(_15993_),
    .Z(\core.muxed_new_block[104] ));
 MUX2_X1 _41091_ (.A(\core.dec_block.block_w0_reg[9] ),
    .B(_10682_),
    .S(_15993_),
    .Z(\core.muxed_new_block[105] ));
 MUX2_X1 _41092_ (.A(\core.dec_block.block_w0_reg[10] ),
    .B(_07258_),
    .S(_15993_),
    .Z(\core.muxed_new_block[106] ));
 BUF_X4 _41093_ (.A(_15992_),
    .Z(_16037_));
 MUX2_X1 _41094_ (.A(\core.dec_block.block_w0_reg[11] ),
    .B(_07659_),
    .S(_16037_),
    .Z(\core.muxed_new_block[107] ));
 MUX2_X1 _41095_ (.A(\core.dec_block.block_w0_reg[12] ),
    .B(_07813_),
    .S(_16037_),
    .Z(\core.muxed_new_block[108] ));
 MUX2_X1 _41096_ (.A(\core.dec_block.block_w0_reg[13] ),
    .B(_07913_),
    .S(_16037_),
    .Z(\core.muxed_new_block[109] ));
 MUX2_X1 _41097_ (.A(\core.dec_block.block_w3_reg[10] ),
    .B(_10721_),
    .S(_16037_),
    .Z(\core.muxed_new_block[10] ));
 MUX2_X1 _41098_ (.A(_17246_),
    .B(_08056_),
    .S(_16037_),
    .Z(\core.muxed_new_block[110] ));
 MUX2_X1 _41099_ (.A(\core.dec_block.block_w0_reg[15] ),
    .B(_08121_),
    .S(_16037_),
    .Z(\core.muxed_new_block[111] ));
 MUX2_X1 _41100_ (.A(\core.dec_block.block_w0_reg[16] ),
    .B(_08612_),
    .S(_16037_),
    .Z(\core.muxed_new_block[112] ));
 MUX2_X1 _41101_ (.A(\core.dec_block.block_w0_reg[17] ),
    .B(_08614_),
    .S(_16037_),
    .Z(\core.muxed_new_block[113] ));
 MUX2_X1 _41102_ (.A(\core.dec_block.block_w0_reg[18] ),
    .B(_08729_),
    .S(_16037_),
    .Z(\core.muxed_new_block[114] ));
 MUX2_X1 _41103_ (.A(\core.dec_block.block_w0_reg[19] ),
    .B(_08905_),
    .S(_16037_),
    .Z(\core.muxed_new_block[115] ));
 CLKBUF_X3 _41104_ (.A(_15992_),
    .Z(_16038_));
 MUX2_X1 _41105_ (.A(\core.dec_block.block_w0_reg[20] ),
    .B(_09012_),
    .S(_16038_),
    .Z(\core.muxed_new_block[116] ));
 MUX2_X1 _41106_ (.A(\core.dec_block.block_w0_reg[21] ),
    .B(_09139_),
    .S(_16038_),
    .Z(\core.muxed_new_block[117] ));
 MUX2_X1 _41107_ (.A(\core.dec_block.block_w0_reg[22] ),
    .B(_09183_),
    .S(_16038_),
    .Z(\core.muxed_new_block[118] ));
 MUX2_X1 _41108_ (.A(_18574_),
    .B(_09227_),
    .S(_16038_),
    .Z(\core.muxed_new_block[119] ));
 MUX2_X1 _41109_ (.A(_17216_),
    .B(_10739_),
    .S(_16038_),
    .Z(\core.muxed_new_block[11] ));
 MUX2_X1 _41110_ (.A(\core.dec_block.block_w0_reg[24] ),
    .B(_07234_),
    .S(_16038_),
    .Z(\core.muxed_new_block[120] ));
 MUX2_X1 _41111_ (.A(\core.dec_block.block_w0_reg[25] ),
    .B(_08999_),
    .S(_16038_),
    .Z(\core.muxed_new_block[121] ));
 MUX2_X1 _41112_ (.A(\core.dec_block.block_w0_reg[26] ),
    .B(_07643_),
    .S(_16038_),
    .Z(\core.muxed_new_block[122] ));
 MUX2_X1 _41113_ (.A(\core.dec_block.block_w0_reg[27] ),
    .B(_07795_),
    .S(_16038_),
    .Z(\core.muxed_new_block[123] ));
 MUX2_X1 _41114_ (.A(\core.dec_block.block_w0_reg[28] ),
    .B(\core.enc_block.block_w0_reg[28] ),
    .S(_16038_),
    .Z(\core.muxed_new_block[124] ));
 BUF_X4 _41115_ (.A(_15992_),
    .Z(_16039_));
 MUX2_X1 _41116_ (.A(\core.dec_block.block_w0_reg[29] ),
    .B(_08041_),
    .S(_16039_),
    .Z(\core.muxed_new_block[125] ));
 MUX2_X1 _41117_ (.A(\core.dec_block.block_w0_reg[30] ),
    .B(_08107_),
    .S(_16039_),
    .Z(\core.muxed_new_block[126] ));
 MUX2_X1 _41118_ (.A(_04003_),
    .B(_07235_),
    .S(_16039_),
    .Z(\core.muxed_new_block[127] ));
 MUX2_X1 _41119_ (.A(\core.dec_block.block_w3_reg[12] ),
    .B(_10841_),
    .S(_16039_),
    .Z(\core.muxed_new_block[12] ));
 MUX2_X1 _41120_ (.A(\core.dec_block.block_w3_reg[13] ),
    .B(_10854_),
    .S(_16039_),
    .Z(\core.muxed_new_block[13] ));
 MUX2_X1 _41121_ (.A(_17248_),
    .B(_10865_),
    .S(_16039_),
    .Z(\core.muxed_new_block[14] ));
 MUX2_X1 _41122_ (.A(\core.dec_block.block_w3_reg[15] ),
    .B(_10722_),
    .S(_16039_),
    .Z(\core.muxed_new_block[15] ));
 MUX2_X1 _41123_ (.A(\core.dec_block.block_w3_reg[16] ),
    .B(_11052_),
    .S(_16039_),
    .Z(\core.muxed_new_block[16] ));
 MUX2_X1 _41124_ (.A(\core.dec_block.block_w3_reg[17] ),
    .B(_11179_),
    .S(_16039_),
    .Z(\core.muxed_new_block[17] ));
 MUX2_X1 _41125_ (.A(\core.dec_block.block_w3_reg[18] ),
    .B(_11064_),
    .S(_16039_),
    .Z(\core.muxed_new_block[18] ));
 CLKBUF_X3 _41126_ (.A(_15992_),
    .Z(_16040_));
 MUX2_X1 _41127_ (.A(\core.dec_block.block_w3_reg[19] ),
    .B(_11080_),
    .S(_16040_),
    .Z(\core.muxed_new_block[19] ));
 MUX2_X1 _41128_ (.A(\core.dec_block.block_w3_reg[1] ),
    .B(_07645_),
    .S(_16040_),
    .Z(\core.muxed_new_block[1] ));
 MUX2_X1 _41129_ (.A(\core.dec_block.block_w3_reg[20] ),
    .B(\core.enc_block.block_w3_reg[20] ),
    .S(_16040_),
    .Z(\core.muxed_new_block[20] ));
 MUX2_X1 _41130_ (.A(\core.dec_block.block_w3_reg[21] ),
    .B(_11109_),
    .S(_16040_),
    .Z(\core.muxed_new_block[21] ));
 MUX2_X1 _41131_ (.A(\core.dec_block.block_w3_reg[22] ),
    .B(_11123_),
    .S(_16040_),
    .Z(\core.muxed_new_block[22] ));
 MUX2_X1 _41132_ (.A(_18576_),
    .B(_11136_),
    .S(_16040_),
    .Z(\core.muxed_new_block[23] ));
 MUX2_X1 _41133_ (.A(\core.dec_block.block_w3_reg[24] ),
    .B(_11418_),
    .S(_16040_),
    .Z(\core.muxed_new_block[24] ));
 MUX2_X1 _41134_ (.A(\core.dec_block.block_w3_reg[25] ),
    .B(_11560_),
    .S(_16040_),
    .Z(\core.muxed_new_block[25] ));
 MUX2_X1 _41135_ (.A(\core.dec_block.block_w3_reg[26] ),
    .B(\core.enc_block.block_w3_reg[26] ),
    .S(_16040_),
    .Z(\core.muxed_new_block[26] ));
 MUX2_X1 _41136_ (.A(\core.dec_block.block_w3_reg[27] ),
    .B(_11443_),
    .S(_16040_),
    .Z(\core.muxed_new_block[27] ));
 CLKBUF_X3 _41137_ (.A(_15992_),
    .Z(_16041_));
 MUX2_X1 _41138_ (.A(\core.dec_block.block_w3_reg[28] ),
    .B(_11457_),
    .S(_16041_),
    .Z(\core.muxed_new_block[28] ));
 MUX2_X1 _41139_ (.A(\core.dec_block.block_w3_reg[29] ),
    .B(_11473_),
    .S(_16041_),
    .Z(\core.muxed_new_block[29] ));
 MUX2_X1 _41140_ (.A(\core.dec_block.block_w3_reg[2] ),
    .B(_07648_),
    .S(_16041_),
    .Z(\core.muxed_new_block[2] ));
 MUX2_X1 _41141_ (.A(\core.dec_block.block_w3_reg[30] ),
    .B(_11487_),
    .S(_16041_),
    .Z(\core.muxed_new_block[30] ));
 MUX2_X1 _41142_ (.A(\core.dec_block.block_w3_reg[31] ),
    .B(_11417_),
    .S(_16041_),
    .Z(\core.muxed_new_block[31] ));
 MUX2_X1 _41143_ (.A(\core.dec_block.block_w2_reg[0] ),
    .B(_06861_),
    .S(_16041_),
    .Z(\core.muxed_new_block[32] ));
 MUX2_X1 _41144_ (.A(\core.dec_block.block_w2_reg[1] ),
    .B(_06800_),
    .S(_16041_),
    .Z(\core.muxed_new_block[33] ));
 MUX2_X1 _41145_ (.A(\core.dec_block.block_w2_reg[2] ),
    .B(_06788_),
    .S(_16041_),
    .Z(\core.muxed_new_block[34] ));
 MUX2_X1 _41146_ (.A(\core.dec_block.block_w2_reg[3] ),
    .B(_06714_),
    .S(_16041_),
    .Z(\core.muxed_new_block[35] ));
 MUX2_X1 _41147_ (.A(\core.dec_block.block_w2_reg[4] ),
    .B(_06768_),
    .S(_16041_),
    .Z(\core.muxed_new_block[36] ));
 CLKBUF_X3 _41148_ (.A(_15992_),
    .Z(_16042_));
 MUX2_X1 _41149_ (.A(\core.dec_block.block_w2_reg[5] ),
    .B(_06761_),
    .S(_16042_),
    .Z(\core.muxed_new_block[37] ));
 MUX2_X1 _41150_ (.A(_16589_),
    .B(_06748_),
    .S(_16042_),
    .Z(\core.muxed_new_block[38] ));
 MUX2_X1 _41151_ (.A(\core.dec_block.block_w2_reg[7] ),
    .B(_06737_),
    .S(_16042_),
    .Z(\core.muxed_new_block[39] ));
 MUX2_X1 _41152_ (.A(\core.dec_block.block_w3_reg[3] ),
    .B(_07790_),
    .S(_16042_),
    .Z(\core.muxed_new_block[3] ));
 MUX2_X1 _41153_ (.A(\core.dec_block.block_w2_reg[8] ),
    .B(_07237_),
    .S(_16042_),
    .Z(\core.muxed_new_block[40] ));
 MUX2_X1 _41154_ (.A(\core.dec_block.block_w2_reg[9] ),
    .B(_07292_),
    .S(_16042_),
    .Z(\core.muxed_new_block[41] ));
 MUX2_X1 _41155_ (.A(\core.dec_block.block_w2_reg[10] ),
    .B(_07274_),
    .S(_16042_),
    .Z(\core.muxed_new_block[42] ));
 MUX2_X1 _41156_ (.A(\core.dec_block.block_w2_reg[11] ),
    .B(_07283_),
    .S(_16042_),
    .Z(\core.muxed_new_block[43] ));
 MUX2_X1 _41157_ (.A(\core.dec_block.block_w2_reg[12] ),
    .B(_07317_),
    .S(_16042_),
    .Z(\core.muxed_new_block[44] ));
 MUX2_X1 _41158_ (.A(\core.dec_block.block_w2_reg[13] ),
    .B(_07306_),
    .S(_16042_),
    .Z(\core.muxed_new_block[45] ));
 BUF_X4 _41159_ (.A(_15992_),
    .Z(_16043_));
 MUX2_X1 _41160_ (.A(\core.dec_block.block_w2_reg[14] ),
    .B(_07329_),
    .S(_16043_),
    .Z(\core.muxed_new_block[46] ));
 MUX2_X1 _41161_ (.A(\core.dec_block.block_w2_reg[15] ),
    .B(_07338_),
    .S(_16043_),
    .Z(\core.muxed_new_block[47] ));
 MUX2_X1 _41162_ (.A(\core.dec_block.block_w2_reg[16] ),
    .B(_08178_),
    .S(_16043_),
    .Z(\core.muxed_new_block[48] ));
 MUX2_X1 _41163_ (.A(\core.dec_block.block_w2_reg[17] ),
    .B(_08185_),
    .S(_16043_),
    .Z(\core.muxed_new_block[49] ));
 MUX2_X1 _41164_ (.A(\core.dec_block.block_w3_reg[4] ),
    .B(_07897_),
    .S(_16043_),
    .Z(\core.muxed_new_block[4] ));
 MUX2_X1 _41165_ (.A(\core.dec_block.block_w2_reg[18] ),
    .B(_08199_),
    .S(_16043_),
    .Z(\core.muxed_new_block[50] ));
 MUX2_X1 _41166_ (.A(\core.dec_block.block_w2_reg[19] ),
    .B(_08207_),
    .S(_16043_),
    .Z(\core.muxed_new_block[51] ));
 MUX2_X1 _41167_ (.A(\core.dec_block.block_w2_reg[20] ),
    .B(_08218_),
    .S(_16043_),
    .Z(\core.muxed_new_block[52] ));
 MUX2_X1 _41168_ (.A(\core.dec_block.block_w2_reg[21] ),
    .B(_08225_),
    .S(_16043_),
    .Z(\core.muxed_new_block[53] ));
 MUX2_X1 _41169_ (.A(\core.dec_block.block_w2_reg[22] ),
    .B(_08243_),
    .S(_16043_),
    .Z(\core.muxed_new_block[54] ));
 CLKBUF_X3 _41170_ (.A(_15992_),
    .Z(_16044_));
 MUX2_X1 _41171_ (.A(_17537_),
    .B(_08236_),
    .S(_16044_),
    .Z(\core.muxed_new_block[55] ));
 MUX2_X1 _41172_ (.A(\core.dec_block.block_w2_reg[24] ),
    .B(_09321_),
    .S(_16044_),
    .Z(\core.muxed_new_block[56] ));
 MUX2_X1 _41173_ (.A(\core.dec_block.block_w2_reg[25] ),
    .B(_09310_),
    .S(_16044_),
    .Z(\core.muxed_new_block[57] ));
 MUX2_X1 _41174_ (.A(\core.dec_block.block_w2_reg[26] ),
    .B(_09243_),
    .S(_16044_),
    .Z(\core.muxed_new_block[58] ));
 MUX2_X1 _41175_ (.A(\core.dec_block.block_w2_reg[27] ),
    .B(_09231_),
    .S(_16044_),
    .Z(\core.muxed_new_block[59] ));
 MUX2_X1 _41176_ (.A(\core.dec_block.block_w3_reg[5] ),
    .B(_08043_),
    .S(_16044_),
    .Z(\core.muxed_new_block[5] ));
 MUX2_X1 _41177_ (.A(\core.dec_block.block_w2_reg[28] ),
    .B(\core.enc_block.block_w2_reg[28] ),
    .S(_16044_),
    .Z(\core.muxed_new_block[60] ));
 MUX2_X1 _41178_ (.A(\core.dec_block.block_w2_reg[29] ),
    .B(_09275_),
    .S(_16044_),
    .Z(\core.muxed_new_block[61] ));
 MUX2_X1 _41179_ (.A(\core.dec_block.block_w2_reg[30] ),
    .B(_09262_),
    .S(_16044_),
    .Z(\core.muxed_new_block[62] ));
 MUX2_X1 _41180_ (.A(\core.dec_block.block_w2_reg[31] ),
    .B(_09255_),
    .S(_16044_),
    .Z(\core.muxed_new_block[63] ));
 CLKBUF_X3 _41181_ (.A(_15992_),
    .Z(_16045_));
 MUX2_X1 _41182_ (.A(\core.dec_block.block_w1_reg[0] ),
    .B(_06863_),
    .S(_16045_),
    .Z(\core.muxed_new_block[64] ));
 MUX2_X1 _41183_ (.A(\core.dec_block.block_w1_reg[1] ),
    .B(_06802_),
    .S(_16045_),
    .Z(\core.muxed_new_block[65] ));
 MUX2_X1 _41184_ (.A(\core.dec_block.block_w1_reg[2] ),
    .B(_06790_),
    .S(_16045_),
    .Z(\core.muxed_new_block[66] ));
 MUX2_X1 _41185_ (.A(\core.dec_block.block_w1_reg[3] ),
    .B(_06721_),
    .S(_16045_),
    .Z(\core.muxed_new_block[67] ));
 MUX2_X1 _41186_ (.A(\core.dec_block.block_w1_reg[4] ),
    .B(_06770_),
    .S(_16045_),
    .Z(\core.muxed_new_block[68] ));
 MUX2_X1 _41187_ (.A(\core.dec_block.block_w1_reg[5] ),
    .B(_06763_),
    .S(_16045_),
    .Z(\core.muxed_new_block[69] ));
 MUX2_X1 _41188_ (.A(\core.dec_block.block_w3_reg[6] ),
    .B(_08110_),
    .S(_16045_),
    .Z(\core.muxed_new_block[6] ));
 MUX2_X1 _41189_ (.A(\core.dec_block.block_w1_reg[6] ),
    .B(_06751_),
    .S(_16045_),
    .Z(\core.muxed_new_block[70] ));
 MUX2_X1 _41190_ (.A(\core.dec_block.block_w1_reg[7] ),
    .B(_06740_),
    .S(_16045_),
    .Z(\core.muxed_new_block[71] ));
 MUX2_X1 _41191_ (.A(\core.dec_block.block_w1_reg[8] ),
    .B(_07267_),
    .S(_16045_),
    .Z(\core.muxed_new_block[72] ));
 BUF_X4 _41192_ (.A(_16203_),
    .Z(_16046_));
 MUX2_X1 _41193_ (.A(\core.dec_block.block_w1_reg[9] ),
    .B(_07294_),
    .S(_16046_),
    .Z(\core.muxed_new_block[73] ));
 MUX2_X1 _41194_ (.A(\core.dec_block.block_w1_reg[10] ),
    .B(_07276_),
    .S(_16046_),
    .Z(\core.muxed_new_block[74] ));
 MUX2_X1 _41195_ (.A(\core.dec_block.block_w1_reg[11] ),
    .B(_07285_),
    .S(_16046_),
    .Z(\core.muxed_new_block[75] ));
 MUX2_X1 _41196_ (.A(\core.dec_block.block_w1_reg[12] ),
    .B(_07319_),
    .S(_16046_),
    .Z(\core.muxed_new_block[76] ));
 MUX2_X1 _41197_ (.A(\core.dec_block.block_w1_reg[13] ),
    .B(_07308_),
    .S(_16046_),
    .Z(\core.muxed_new_block[77] ));
 MUX2_X1 _41198_ (.A(\core.dec_block.block_w1_reg[14] ),
    .B(_07331_),
    .S(_16046_),
    .Z(\core.muxed_new_block[78] ));
 MUX2_X1 _41199_ (.A(\core.dec_block.block_w1_reg[15] ),
    .B(_07340_),
    .S(_16046_),
    .Z(\core.muxed_new_block[79] ));
 MUX2_X1 _41200_ (.A(\core.dec_block.block_w3_reg[7] ),
    .B(_07791_),
    .S(_16046_),
    .Z(\core.muxed_new_block[7] ));
 MUX2_X1 _41201_ (.A(\core.dec_block.block_w1_reg[16] ),
    .B(_07238_),
    .S(_16046_),
    .Z(\core.muxed_new_block[80] ));
 MUX2_X1 _41202_ (.A(\core.dec_block.block_w1_reg[17] ),
    .B(_08187_),
    .S(_16046_),
    .Z(\core.muxed_new_block[81] ));
 BUF_X4 _41203_ (.A(_16203_),
    .Z(_16047_));
 MUX2_X1 _41204_ (.A(\core.dec_block.block_w1_reg[18] ),
    .B(_07644_),
    .S(_16047_),
    .Z(\core.muxed_new_block[82] ));
 MUX2_X1 _41205_ (.A(\core.dec_block.block_w1_reg[19] ),
    .B(_07794_),
    .S(_16047_),
    .Z(\core.muxed_new_block[83] ));
 MUX2_X1 _41206_ (.A(\core.dec_block.block_w1_reg[20] ),
    .B(_07895_),
    .S(_16047_),
    .Z(\core.muxed_new_block[84] ));
 MUX2_X1 _41207_ (.A(\core.dec_block.block_w1_reg[21] ),
    .B(_08040_),
    .S(_16047_),
    .Z(\core.muxed_new_block[85] ));
 MUX2_X1 _41208_ (.A(\core.dec_block.block_w1_reg[22] ),
    .B(_08106_),
    .S(_16047_),
    .Z(\core.muxed_new_block[86] ));
 MUX2_X1 _41209_ (.A(_18577_),
    .B(_08165_),
    .S(_16047_),
    .Z(\core.muxed_new_block[87] ));
 MUX2_X1 _41210_ (.A(\core.dec_block.block_w1_reg[24] ),
    .B(_09323_),
    .S(_16047_),
    .Z(\core.muxed_new_block[88] ));
 MUX2_X1 _41211_ (.A(\core.dec_block.block_w1_reg[25] ),
    .B(_09312_),
    .S(_16047_),
    .Z(\core.muxed_new_block[89] ));
 MUX2_X1 _41212_ (.A(\core.dec_block.block_w3_reg[8] ),
    .B(\core.enc_block.block_w3_reg[8] ),
    .S(_16047_),
    .Z(\core.muxed_new_block[8] ));
 MUX2_X1 _41213_ (.A(\core.dec_block.block_w1_reg[26] ),
    .B(_09240_),
    .S(_16047_),
    .Z(\core.muxed_new_block[90] ));
 CLKBUF_X3 _41214_ (.A(_16203_),
    .Z(_16048_));
 MUX2_X1 _41215_ (.A(\core.dec_block.block_w1_reg[27] ),
    .B(_09233_),
    .S(_16048_),
    .Z(\core.muxed_new_block[91] ));
 MUX2_X1 _41216_ (.A(\core.dec_block.block_w1_reg[28] ),
    .B(_09285_),
    .S(_16048_),
    .Z(\core.muxed_new_block[92] ));
 MUX2_X1 _41217_ (.A(\core.dec_block.block_w1_reg[29] ),
    .B(_09277_),
    .S(_16048_),
    .Z(\core.muxed_new_block[93] ));
 MUX2_X1 _41218_ (.A(\core.dec_block.block_w1_reg[30] ),
    .B(_09260_),
    .S(_16048_),
    .Z(\core.muxed_new_block[94] ));
 MUX2_X1 _41219_ (.A(\core.dec_block.block_w1_reg[31] ),
    .B(_09253_),
    .S(_16048_),
    .Z(\core.muxed_new_block[95] ));
 MUX2_X1 _41220_ (.A(\core.dec_block.block_w0_reg[0] ),
    .B(\core.enc_block.block_w0_reg[0] ),
    .S(_16048_),
    .Z(\core.muxed_new_block[96] ));
 MUX2_X1 _41221_ (.A(\core.dec_block.block_w0_reg[1] ),
    .B(\core.enc_block.block_w0_reg[1] ),
    .S(_16048_),
    .Z(\core.muxed_new_block[97] ));
 MUX2_X1 _41222_ (.A(\core.dec_block.block_w0_reg[2] ),
    .B(_10088_),
    .S(_16048_),
    .Z(\core.muxed_new_block[98] ));
 MUX2_X1 _41223_ (.A(\core.dec_block.block_w0_reg[3] ),
    .B(_10274_),
    .S(_16048_),
    .Z(\core.muxed_new_block[99] ));
 MUX2_X1 _41224_ (.A(\core.dec_block.block_w3_reg[9] ),
    .B(_10796_),
    .S(_16048_),
    .Z(\core.muxed_new_block[9] ));
 NAND3_X1 _41225_ (.A1(_22100_),
    .A2(_16299_),
    .A3(_15996_),
    .ZN(_16049_));
 NOR2_X1 _41226_ (.A1(_16297_),
    .A2(_16049_),
    .ZN(_16050_));
 AND2_X1 _41227_ (.A1(_16289_),
    .A2(_16050_),
    .ZN(init_new));
 AND2_X1 _41228_ (.A1(_16313_),
    .A2(_16050_),
    .ZN(next_new));
 INV_X1 _41229_ (.A(net17),
    .ZN(_16051_));
 NAND2_X4 _41230_ (.A1(_16051_),
    .A2(net8),
    .ZN(_16052_));
 NOR2_X4 _41231_ (.A1(_15999_),
    .A2(_16296_),
    .ZN(_16053_));
 NOR2_X2 _41232_ (.A1(net2),
    .A2(_22097_),
    .ZN(_16054_));
 AND2_X1 _41233_ (.A1(_16053_),
    .A2(_16054_),
    .ZN(_16055_));
 CLKBUF_X3 _41234_ (.A(_16055_),
    .Z(_16056_));
 MUX2_X1 _41235_ (.A(\result_reg[96] ),
    .B(\result_reg[64] ),
    .S(_16341_),
    .Z(_16057_));
 CLKBUF_X3 _41236_ (.A(_16292_),
    .Z(_16058_));
 MUX2_X1 _41237_ (.A(\result_reg[32] ),
    .B(\result_reg[0] ),
    .S(_16058_),
    .Z(_16059_));
 CLKBUF_X3 _41238_ (.A(_16335_),
    .Z(_16060_));
 MUX2_X1 _41239_ (.A(_16057_),
    .B(_16059_),
    .S(_16060_),
    .Z(_16061_));
 BUF_X4 _41240_ (.A(_16335_),
    .Z(_16062_));
 NOR2_X2 _41241_ (.A1(_16062_),
    .A2(_15997_),
    .ZN(_16063_));
 BUF_X4 _41242_ (.A(_16341_),
    .Z(_16064_));
 MUX2_X1 _41243_ (.A(_16210_),
    .B(ready_reg),
    .S(_16064_),
    .Z(_16065_));
 AOI22_X2 _41244_ (.A1(_16056_),
    .A2(_16061_),
    .B1(_16063_),
    .B2(_16065_),
    .ZN(_16066_));
 NOR2_X2 _41245_ (.A1(_16052_),
    .A2(_16066_),
    .ZN(net50));
 AND2_X2 _41246_ (.A1(_16051_),
    .A2(net8),
    .ZN(_16067_));
 NAND2_X2 _41247_ (.A1(_22096_),
    .A2(_15996_),
    .ZN(_16068_));
 NOR2_X2 _41248_ (.A1(_15994_),
    .A2(_16068_),
    .ZN(_16069_));
 OAI21_X4 _41249_ (.A(_16067_),
    .B1(_16053_),
    .B2(_16069_),
    .ZN(_16070_));
 CLKBUF_X3 _41250_ (.A(_16054_),
    .Z(_16071_));
 BUF_X4 _41251_ (.A(_16292_),
    .Z(_16072_));
 MUX2_X1 _41252_ (.A(\result_reg[106] ),
    .B(\result_reg[74] ),
    .S(_16072_),
    .Z(_16073_));
 BUF_X4 _41253_ (.A(_16292_),
    .Z(_16074_));
 MUX2_X1 _41254_ (.A(\result_reg[42] ),
    .B(\result_reg[10] ),
    .S(_16074_),
    .Z(_16075_));
 BUF_X4 _41255_ (.A(_16335_),
    .Z(_16076_));
 MUX2_X1 _41256_ (.A(_16073_),
    .B(_16075_),
    .S(_16076_),
    .Z(_16077_));
 NAND2_X1 _41257_ (.A1(_16071_),
    .A2(_16077_),
    .ZN(_16078_));
 BUF_X8 _41258_ (.A(_16053_),
    .Z(_16079_));
 AOI21_X2 _41259_ (.A(_16070_),
    .B1(_16078_),
    .B2(_16079_),
    .ZN(net51));
 AND2_X2 _41260_ (.A1(_16067_),
    .A2(_16056_),
    .ZN(_16080_));
 CLKBUF_X3 _41261_ (.A(_16341_),
    .Z(_16081_));
 MUX2_X1 _41262_ (.A(\result_reg[107] ),
    .B(\result_reg[75] ),
    .S(_16081_),
    .Z(_16082_));
 MUX2_X1 _41263_ (.A(\result_reg[43] ),
    .B(\result_reg[11] ),
    .S(_16064_),
    .Z(_16083_));
 MUX2_X1 _41264_ (.A(_16082_),
    .B(_16083_),
    .S(_16062_),
    .Z(_16084_));
 AND2_X1 _41265_ (.A1(_16080_),
    .A2(_16084_),
    .ZN(net52));
 NAND3_X4 _41266_ (.A1(_16293_),
    .A2(_22096_),
    .A3(_15996_),
    .ZN(_16085_));
 MUX2_X1 _41267_ (.A(\result_reg[108] ),
    .B(\result_reg[76] ),
    .S(_16058_),
    .Z(_16086_));
 MUX2_X1 _41268_ (.A(\result_reg[44] ),
    .B(\result_reg[12] ),
    .S(_16058_),
    .Z(_16087_));
 MUX2_X1 _41269_ (.A(_16086_),
    .B(_16087_),
    .S(_16060_),
    .Z(_16088_));
 NAND2_X1 _41270_ (.A1(_16056_),
    .A2(_16088_),
    .ZN(_16089_));
 AOI21_X4 _41271_ (.A(_16052_),
    .B1(_16085_),
    .B2(_16089_),
    .ZN(net53));
 NOR2_X2 _41272_ (.A1(_16294_),
    .A2(_16068_),
    .ZN(_16090_));
 OAI21_X4 _41273_ (.A(_16067_),
    .B1(_16053_),
    .B2(_16090_),
    .ZN(_16091_));
 MUX2_X1 _41274_ (.A(\result_reg[109] ),
    .B(\result_reg[77] ),
    .S(_16072_),
    .Z(_16092_));
 MUX2_X1 _41275_ (.A(\result_reg[45] ),
    .B(\result_reg[13] ),
    .S(_16074_),
    .Z(_16093_));
 MUX2_X1 _41276_ (.A(_16092_),
    .B(_16093_),
    .S(_16076_),
    .Z(_16094_));
 NAND2_X1 _41277_ (.A1(_16071_),
    .A2(_16094_),
    .ZN(_16095_));
 AOI21_X4 _41278_ (.A(_16091_),
    .B1(_16095_),
    .B2(_16079_),
    .ZN(net54));
 NOR3_X2 _41279_ (.A1(_16335_),
    .A2(_16064_),
    .A3(_16068_),
    .ZN(_16096_));
 OAI21_X4 _41280_ (.A(_16067_),
    .B1(_16053_),
    .B2(_16096_),
    .ZN(_16097_));
 BUF_X4 _41281_ (.A(_16292_),
    .Z(_16098_));
 MUX2_X1 _41282_ (.A(\result_reg[110] ),
    .B(\result_reg[78] ),
    .S(_16098_),
    .Z(_16099_));
 MUX2_X1 _41283_ (.A(\result_reg[46] ),
    .B(\result_reg[14] ),
    .S(_16074_),
    .Z(_16100_));
 MUX2_X1 _41284_ (.A(_16099_),
    .B(_16100_),
    .S(_16076_),
    .Z(_16101_));
 NAND2_X1 _41285_ (.A1(_16071_),
    .A2(_16101_),
    .ZN(_16102_));
 AOI21_X2 _41286_ (.A(_16097_),
    .B1(_16102_),
    .B2(_16079_),
    .ZN(net55));
 MUX2_X1 _41287_ (.A(\result_reg[111] ),
    .B(\result_reg[79] ),
    .S(_16081_),
    .Z(_16103_));
 MUX2_X1 _41288_ (.A(\result_reg[47] ),
    .B(\result_reg[15] ),
    .S(_16064_),
    .Z(_16104_));
 MUX2_X1 _41289_ (.A(_16103_),
    .B(_16104_),
    .S(_16062_),
    .Z(_16105_));
 AND2_X1 _41290_ (.A1(_16080_),
    .A2(_16105_),
    .ZN(net56));
 MUX2_X1 _41291_ (.A(\result_reg[112] ),
    .B(\result_reg[80] ),
    .S(_16098_),
    .Z(_16106_));
 MUX2_X1 _41292_ (.A(\result_reg[48] ),
    .B(\result_reg[16] ),
    .S(_16074_),
    .Z(_16107_));
 MUX2_X1 _41293_ (.A(_16106_),
    .B(_16107_),
    .S(_16076_),
    .Z(_16108_));
 NAND2_X1 _41294_ (.A1(_16071_),
    .A2(_16108_),
    .ZN(_16109_));
 AOI21_X2 _41295_ (.A(_16097_),
    .B1(_16109_),
    .B2(_16079_),
    .ZN(net57));
 MUX2_X1 _41296_ (.A(\result_reg[113] ),
    .B(\result_reg[81] ),
    .S(_16098_),
    .Z(_16110_));
 MUX2_X1 _41297_ (.A(\result_reg[49] ),
    .B(\result_reg[17] ),
    .S(_16074_),
    .Z(_16111_));
 MUX2_X1 _41298_ (.A(_16110_),
    .B(_16111_),
    .S(_16076_),
    .Z(_16112_));
 NAND2_X1 _41299_ (.A1(_16071_),
    .A2(_16112_),
    .ZN(_16113_));
 AOI21_X2 _41300_ (.A(_16070_),
    .B1(_16113_),
    .B2(_16079_),
    .ZN(net58));
 MUX2_X1 _41301_ (.A(\result_reg[114] ),
    .B(\result_reg[82] ),
    .S(_16058_),
    .Z(_16114_));
 MUX2_X1 _41302_ (.A(\result_reg[50] ),
    .B(\result_reg[18] ),
    .S(_16058_),
    .Z(_16115_));
 MUX2_X1 _41303_ (.A(_16114_),
    .B(_16115_),
    .S(_16060_),
    .Z(_16116_));
 NAND2_X1 _41304_ (.A1(_16056_),
    .A2(_16116_),
    .ZN(_16117_));
 AOI21_X4 _41305_ (.A(_16052_),
    .B1(_16085_),
    .B2(_16117_),
    .ZN(net59));
 MUX2_X1 _41306_ (.A(\result_reg[115] ),
    .B(\result_reg[83] ),
    .S(_16098_),
    .Z(_16118_));
 MUX2_X1 _41307_ (.A(\result_reg[51] ),
    .B(\result_reg[19] ),
    .S(_16074_),
    .Z(_16119_));
 MUX2_X1 _41308_ (.A(_16118_),
    .B(_16119_),
    .S(_16076_),
    .Z(_16120_));
 NAND2_X1 _41309_ (.A1(_16071_),
    .A2(_16120_),
    .ZN(_16121_));
 AOI21_X2 _41310_ (.A(_16070_),
    .B1(_16121_),
    .B2(_16079_),
    .ZN(net60));
 MUX2_X1 _41311_ (.A(\result_reg[97] ),
    .B(\result_reg[65] ),
    .S(_16341_),
    .Z(_16122_));
 MUX2_X1 _41312_ (.A(\result_reg[33] ),
    .B(\result_reg[1] ),
    .S(_16341_),
    .Z(_16123_));
 MUX2_X1 _41313_ (.A(_16122_),
    .B(_16123_),
    .S(_16335_),
    .Z(_16124_));
 MUX2_X1 _41314_ (.A(_16206_),
    .B(valid_reg),
    .S(_16064_),
    .Z(_16125_));
 AOI22_X2 _41315_ (.A1(_16056_),
    .A2(_16124_),
    .B1(_16125_),
    .B2(_16063_),
    .ZN(_16126_));
 NOR2_X2 _41316_ (.A1(_16052_),
    .A2(_16126_),
    .ZN(net61));
 MUX2_X1 _41317_ (.A(\result_reg[116] ),
    .B(\result_reg[84] ),
    .S(_16081_),
    .Z(_16127_));
 MUX2_X1 _41318_ (.A(\result_reg[52] ),
    .B(\result_reg[20] ),
    .S(_16064_),
    .Z(_16128_));
 MUX2_X1 _41319_ (.A(_16127_),
    .B(_16128_),
    .S(_16062_),
    .Z(_16129_));
 AND2_X1 _41320_ (.A1(_16080_),
    .A2(_16129_),
    .ZN(net62));
 MUX2_X1 _41321_ (.A(\result_reg[117] ),
    .B(\result_reg[85] ),
    .S(_16098_),
    .Z(_16130_));
 MUX2_X1 _41322_ (.A(\result_reg[53] ),
    .B(\result_reg[21] ),
    .S(_16074_),
    .Z(_16131_));
 MUX2_X1 _41323_ (.A(_16130_),
    .B(_16131_),
    .S(_16076_),
    .Z(_16132_));
 NAND2_X1 _41324_ (.A1(_16071_),
    .A2(_16132_),
    .ZN(_16133_));
 AOI21_X4 _41325_ (.A(_16091_),
    .B1(_16133_),
    .B2(_16079_),
    .ZN(net63));
 MUX2_X1 _41326_ (.A(\result_reg[118] ),
    .B(\result_reg[86] ),
    .S(_16098_),
    .Z(_16134_));
 MUX2_X1 _41327_ (.A(\result_reg[54] ),
    .B(\result_reg[22] ),
    .S(_16072_),
    .Z(_16135_));
 MUX2_X1 _41328_ (.A(_16134_),
    .B(_16135_),
    .S(_16076_),
    .Z(_16136_));
 NAND2_X1 _41329_ (.A1(_16071_),
    .A2(_16136_),
    .ZN(_16137_));
 AOI21_X2 _41330_ (.A(_16097_),
    .B1(_16137_),
    .B2(_16079_),
    .ZN(net64));
 MUX2_X1 _41331_ (.A(\result_reg[119] ),
    .B(\result_reg[87] ),
    .S(_16081_),
    .Z(_16138_));
 MUX2_X1 _41332_ (.A(\result_reg[55] ),
    .B(\result_reg[23] ),
    .S(_16064_),
    .Z(_16139_));
 MUX2_X1 _41333_ (.A(_16138_),
    .B(_16139_),
    .S(_16062_),
    .Z(_16140_));
 AND2_X1 _41334_ (.A1(_16080_),
    .A2(_16140_),
    .ZN(net65));
 MUX2_X1 _41335_ (.A(\result_reg[120] ),
    .B(\result_reg[88] ),
    .S(_16098_),
    .Z(_16141_));
 MUX2_X1 _41336_ (.A(\result_reg[56] ),
    .B(\result_reg[24] ),
    .S(_16072_),
    .Z(_16142_));
 MUX2_X1 _41337_ (.A(_16141_),
    .B(_16142_),
    .S(_16076_),
    .Z(_16143_));
 NAND2_X1 _41338_ (.A1(_16071_),
    .A2(_16143_),
    .ZN(_16144_));
 AOI21_X4 _41339_ (.A(_16097_),
    .B1(_16144_),
    .B2(_16079_),
    .ZN(net66));
 MUX2_X1 _41340_ (.A(\result_reg[121] ),
    .B(\result_reg[89] ),
    .S(_16081_),
    .Z(_16145_));
 MUX2_X1 _41341_ (.A(\result_reg[57] ),
    .B(\result_reg[25] ),
    .S(_16064_),
    .Z(_16146_));
 MUX2_X1 _41342_ (.A(_16145_),
    .B(_16146_),
    .S(_16062_),
    .Z(_16147_));
 AND2_X1 _41343_ (.A1(_16080_),
    .A2(_16147_),
    .ZN(net67));
 MUX2_X1 _41344_ (.A(\result_reg[122] ),
    .B(\result_reg[90] ),
    .S(_16081_),
    .Z(_16148_));
 MUX2_X1 _41345_ (.A(\result_reg[58] ),
    .B(\result_reg[26] ),
    .S(_16064_),
    .Z(_16149_));
 MUX2_X1 _41346_ (.A(_16148_),
    .B(_16149_),
    .S(_16062_),
    .Z(_16150_));
 AND2_X1 _41347_ (.A1(_16080_),
    .A2(_16150_),
    .ZN(net68));
 MUX2_X1 _41348_ (.A(\result_reg[123] ),
    .B(\result_reg[91] ),
    .S(_16081_),
    .Z(_16151_));
 MUX2_X1 _41349_ (.A(\result_reg[59] ),
    .B(\result_reg[27] ),
    .S(_16064_),
    .Z(_16152_));
 MUX2_X1 _41350_ (.A(_16151_),
    .B(_16152_),
    .S(_16062_),
    .Z(_16153_));
 AND2_X1 _41351_ (.A1(_16080_),
    .A2(_16153_),
    .ZN(net69));
 MUX2_X1 _41352_ (.A(\result_reg[124] ),
    .B(\result_reg[92] ),
    .S(_16098_),
    .Z(_16154_));
 MUX2_X1 _41353_ (.A(\result_reg[60] ),
    .B(\result_reg[28] ),
    .S(_16072_),
    .Z(_16155_));
 MUX2_X1 _41354_ (.A(_16154_),
    .B(_16155_),
    .S(_16060_),
    .Z(_16156_));
 NAND2_X1 _41355_ (.A1(_16071_),
    .A2(_16156_),
    .ZN(_16157_));
 AOI21_X2 _41356_ (.A(_16070_),
    .B1(_16157_),
    .B2(_16079_),
    .ZN(net70));
 MUX2_X1 _41357_ (.A(\result_reg[125] ),
    .B(\result_reg[93] ),
    .S(_16098_),
    .Z(_16158_));
 MUX2_X1 _41358_ (.A(\result_reg[61] ),
    .B(\result_reg[29] ),
    .S(_16072_),
    .Z(_16159_));
 MUX2_X1 _41359_ (.A(_16158_),
    .B(_16159_),
    .S(_16060_),
    .Z(_16160_));
 NAND2_X1 _41360_ (.A1(_16054_),
    .A2(_16160_),
    .ZN(_16161_));
 AOI21_X4 _41361_ (.A(_16091_),
    .B1(_16161_),
    .B2(_16053_),
    .ZN(net71));
 INV_X1 _41362_ (.A(_16049_),
    .ZN(_16162_));
 MUX2_X1 _41363_ (.A(\result_reg[98] ),
    .B(\result_reg[66] ),
    .S(_16341_),
    .Z(_16163_));
 MUX2_X1 _41364_ (.A(\result_reg[34] ),
    .B(\result_reg[2] ),
    .S(_16341_),
    .Z(_16164_));
 MUX2_X1 _41365_ (.A(_16163_),
    .B(_16164_),
    .S(_16335_),
    .Z(_16165_));
 AOI22_X2 _41366_ (.A1(_15993_),
    .A2(_16162_),
    .B1(_16056_),
    .B2(_16165_),
    .ZN(_16166_));
 NOR2_X2 _41367_ (.A1(_16052_),
    .A2(_16166_),
    .ZN(net72));
 MUX2_X1 _41368_ (.A(\result_reg[126] ),
    .B(\result_reg[94] ),
    .S(_16098_),
    .Z(_16167_));
 MUX2_X1 _41369_ (.A(\result_reg[62] ),
    .B(\result_reg[30] ),
    .S(_16072_),
    .Z(_16168_));
 MUX2_X1 _41370_ (.A(_16167_),
    .B(_16168_),
    .S(_16060_),
    .Z(_16169_));
 NAND2_X1 _41371_ (.A1(_16054_),
    .A2(_16169_),
    .ZN(_16170_));
 AOI21_X4 _41372_ (.A(_16097_),
    .B1(_16170_),
    .B2(_16053_),
    .ZN(net73));
 MUX2_X1 _41373_ (.A(\result_reg[127] ),
    .B(\result_reg[95] ),
    .S(_16074_),
    .Z(_16171_));
 MUX2_X1 _41374_ (.A(\result_reg[63] ),
    .B(\result_reg[31] ),
    .S(_16081_),
    .Z(_16172_));
 MUX2_X1 _41375_ (.A(_16171_),
    .B(_16172_),
    .S(_16062_),
    .Z(_16173_));
 AND2_X1 _41376_ (.A1(_16080_),
    .A2(_16173_),
    .ZN(net74));
 MUX2_X1 _41377_ (.A(\result_reg[99] ),
    .B(\result_reg[67] ),
    .S(_16341_),
    .Z(_16174_));
 MUX2_X1 _41378_ (.A(\result_reg[35] ),
    .B(\result_reg[3] ),
    .S(_16341_),
    .Z(_16175_));
 MUX2_X1 _41379_ (.A(_16174_),
    .B(_16175_),
    .S(_16335_),
    .Z(_16176_));
 AOI22_X2 _41380_ (.A1(_15428_),
    .A2(_16162_),
    .B1(_16056_),
    .B2(_16176_),
    .ZN(_16177_));
 NOR2_X2 _41381_ (.A1(_16052_),
    .A2(_16177_),
    .ZN(net75));
 MUX2_X1 _41382_ (.A(\result_reg[100] ),
    .B(\result_reg[68] ),
    .S(_16058_),
    .Z(_16178_));
 MUX2_X1 _41383_ (.A(\result_reg[36] ),
    .B(\result_reg[4] ),
    .S(_16072_),
    .Z(_16179_));
 MUX2_X1 _41384_ (.A(_16178_),
    .B(_16179_),
    .S(_16060_),
    .Z(_16180_));
 NAND2_X1 _41385_ (.A1(_16054_),
    .A2(_16180_),
    .ZN(_16181_));
 AOI21_X4 _41386_ (.A(_16070_),
    .B1(_16181_),
    .B2(_16053_),
    .ZN(net76));
 MUX2_X1 _41387_ (.A(\result_reg[101] ),
    .B(\result_reg[69] ),
    .S(_16058_),
    .Z(_16182_));
 MUX2_X1 _41388_ (.A(\result_reg[37] ),
    .B(\result_reg[5] ),
    .S(_16072_),
    .Z(_16183_));
 MUX2_X1 _41389_ (.A(_16182_),
    .B(_16183_),
    .S(_16060_),
    .Z(_16184_));
 NAND2_X1 _41390_ (.A1(_16054_),
    .A2(_16184_),
    .ZN(_16185_));
 AOI21_X4 _41391_ (.A(_16091_),
    .B1(_16185_),
    .B2(_16053_),
    .ZN(net77));
 MUX2_X1 _41392_ (.A(\result_reg[102] ),
    .B(\result_reg[70] ),
    .S(_16074_),
    .Z(_16186_));
 MUX2_X1 _41393_ (.A(\result_reg[38] ),
    .B(\result_reg[6] ),
    .S(_16081_),
    .Z(_16187_));
 MUX2_X1 _41394_ (.A(_16186_),
    .B(_16187_),
    .S(_16062_),
    .Z(_16188_));
 AND2_X1 _41395_ (.A1(_16080_),
    .A2(_16188_),
    .ZN(net78));
 MUX2_X1 _41396_ (.A(\result_reg[103] ),
    .B(\result_reg[71] ),
    .S(_16074_),
    .Z(_16189_));
 MUX2_X1 _41397_ (.A(\result_reg[39] ),
    .B(\result_reg[7] ),
    .S(_16081_),
    .Z(_16190_));
 MUX2_X1 _41398_ (.A(_16189_),
    .B(_16190_),
    .S(_16076_),
    .Z(_16191_));
 AND2_X1 _41399_ (.A1(_16080_),
    .A2(_16191_),
    .ZN(net79));
 MUX2_X1 _41400_ (.A(\result_reg[104] ),
    .B(\result_reg[72] ),
    .S(_16058_),
    .Z(_16192_));
 MUX2_X1 _41401_ (.A(\result_reg[40] ),
    .B(\result_reg[8] ),
    .S(_16072_),
    .Z(_16193_));
 MUX2_X1 _41402_ (.A(_16192_),
    .B(_16193_),
    .S(_16060_),
    .Z(_16194_));
 NAND2_X1 _41403_ (.A1(_16054_),
    .A2(_16194_),
    .ZN(_16195_));
 AOI21_X4 _41404_ (.A(_16097_),
    .B1(_16195_),
    .B2(_16053_),
    .ZN(net80));
 MUX2_X1 _41405_ (.A(\result_reg[105] ),
    .B(\result_reg[73] ),
    .S(_16058_),
    .Z(_16196_));
 MUX2_X1 _41406_ (.A(\result_reg[41] ),
    .B(\result_reg[9] ),
    .S(_16058_),
    .Z(_16197_));
 MUX2_X1 _41407_ (.A(_16196_),
    .B(_16197_),
    .S(_16060_),
    .Z(_16198_));
 NAND2_X1 _41408_ (.A1(_16056_),
    .A2(_16198_),
    .ZN(_16199_));
 AOI21_X4 _41409_ (.A(_16052_),
    .B1(_16085_),
    .B2(_16199_),
    .ZN(net81));
 HA_X1 _41410_ (.A(\core.enc_block.round[2] ),
    .B(_22091_),
    .CO(_22092_),
    .S(_22093_));
 HA_X1 _41411_ (.A(_22094_),
    .B(_22095_),
    .CO(_22096_),
    .S(_22097_));
 HA_X1 _41412_ (.A(_22094_),
    .B(_22095_),
    .CO(_22098_),
    .S(_22099_));
 HA_X1 _41413_ (.A(_22094_),
    .B(net3),
    .CO(_22100_),
    .S(_22101_));
 HA_X1 _41414_ (.A(net2),
    .B(_22095_),
    .CO(_22102_),
    .S(_22103_));
 HA_X1 _41415_ (.A(_22104_),
    .B(_22105_),
    .CO(_22106_),
    .S(_22107_));
 HA_X1 _41416_ (.A(_22104_),
    .B(\core.keymem.round_ctr_reg[1] ),
    .CO(_22108_),
    .S(_22109_));
 HA_X1 _41417_ (.A(\core.keymem.round_ctr_reg[0] ),
    .B(_22105_),
    .CO(_22110_),
    .S(_22111_));
 HA_X1 _41418_ (.A(\core.keymem.round_ctr_reg[0] ),
    .B(\core.keymem.round_ctr_reg[1] ),
    .CO(_22112_),
    .S(_22113_));
 HA_X1 _41419_ (.A(\core.enc_block.round[0] ),
    .B(\core.enc_block.round[1] ),
    .CO(_22114_),
    .S(_22115_));
 HA_X1 _41420_ (.A(_22116_),
    .B(_22117_),
    .CO(_22118_),
    .S(_22119_));
 HA_X1 _41421_ (.A(_22116_),
    .B(\core.enc_block.sword_ctr_reg[1] ),
    .CO(_22120_),
    .S(_22121_));
 HA_X1 _41422_ (.A(\core.enc_block.sword_ctr_reg[0] ),
    .B(_22117_),
    .CO(_22122_),
    .S(_22123_));
 HA_X1 _41423_ (.A(\core.enc_block.sword_ctr_reg[0] ),
    .B(\core.enc_block.sword_ctr_reg[1] ),
    .CO(_22124_),
    .S(_22125_));
 HA_X1 _41424_ (.A(_22126_),
    .B(_22127_),
    .CO(_22128_),
    .S(_22129_));
 HA_X1 _41425_ (.A(_22130_),
    .B(_22131_),
    .CO(_22132_),
    .S(_22133_));
 HA_X1 _41426_ (.A(_22130_),
    .B(\core.dec_block.sword_ctr_reg[1] ),
    .CO(_22134_),
    .S(_22135_));
 HA_X1 _41427_ (.A(\core.dec_block.sword_ctr_reg[0] ),
    .B(_22131_),
    .CO(_22136_),
    .S(_22137_));
 HA_X1 _41428_ (.A(\core.dec_block.sword_ctr_reg[0] ),
    .B(\core.dec_block.sword_ctr_reg[1] ),
    .CO(_22138_),
    .S(_22139_));
 DFFR_X2 \block_reg[0][0]$_DFFE_PN0P_  (.D(_00439_),
    .RN(net90),
    .CK(clknet_leaf_297_clk),
    .Q(\block_reg[0][0] ),
    .QN(_21954_));
 DFFR_X2 \block_reg[0][10]$_DFFE_PN0P_  (.D(_00440_),
    .RN(net92),
    .CK(clknet_leaf_270_clk),
    .Q(\block_reg[0][10] ),
    .QN(_21953_));
 DFFR_X2 \block_reg[0][11]$_DFFE_PN0P_  (.D(_00441_),
    .RN(net91),
    .CK(clknet_leaf_270_clk),
    .Q(\block_reg[0][11] ),
    .QN(_21952_));
 DFFR_X1 \block_reg[0][12]$_DFFE_PN0P_  (.D(_00442_),
    .RN(net92),
    .CK(clknet_leaf_271_clk),
    .Q(\block_reg[0][12] ),
    .QN(_21951_));
 DFFR_X1 \block_reg[0][13]$_DFFE_PN0P_  (.D(_00443_),
    .RN(net92),
    .CK(clknet_leaf_270_clk),
    .Q(\block_reg[0][13] ),
    .QN(_21950_));
 DFFR_X1 \block_reg[0][14]$_DFFE_PN0P_  (.D(_00444_),
    .RN(net91),
    .CK(clknet_leaf_290_clk),
    .Q(\block_reg[0][14] ),
    .QN(_21949_));
 DFFR_X2 \block_reg[0][15]$_DFFE_PN0P_  (.D(_00445_),
    .RN(net92),
    .CK(clknet_leaf_271_clk),
    .Q(\block_reg[0][15] ),
    .QN(_21948_));
 DFFR_X2 \block_reg[0][16]$_DFFE_PN0P_  (.D(_00446_),
    .RN(net90),
    .CK(clknet_leaf_297_clk),
    .Q(\block_reg[0][16] ),
    .QN(_21947_));
 DFFR_X2 \block_reg[0][17]$_DFFE_PN0P_  (.D(_00447_),
    .RN(net91),
    .CK(clknet_leaf_289_clk),
    .Q(\block_reg[0][17] ),
    .QN(_21946_));
 DFFR_X2 \block_reg[0][18]$_DFFE_PN0P_  (.D(_00448_),
    .RN(net91),
    .CK(clknet_leaf_273_clk),
    .Q(\block_reg[0][18] ),
    .QN(_21945_));
 DFFR_X2 \block_reg[0][19]$_DFFE_PN0P_  (.D(_00449_),
    .RN(net91),
    .CK(clknet_leaf_285_clk),
    .Q(\block_reg[0][19] ),
    .QN(_21944_));
 DFFR_X1 \block_reg[0][1]$_DFFE_PN0P_  (.D(_00450_),
    .RN(net85),
    .CK(clknet_leaf_361_clk),
    .Q(\block_reg[0][1] ),
    .QN(_21943_));
 DFFR_X2 \block_reg[0][20]$_DFFE_PN0P_  (.D(_00451_),
    .RN(net93),
    .CK(clknet_leaf_373_clk),
    .Q(\block_reg[0][20] ),
    .QN(_21942_));
 DFFR_X2 \block_reg[0][21]$_DFFE_PN0P_  (.D(_00452_),
    .RN(net93),
    .CK(clknet_leaf_362_clk),
    .Q(\block_reg[0][21] ),
    .QN(_21941_));
 DFFR_X2 \block_reg[0][22]$_DFFE_PN0P_  (.D(_00453_),
    .RN(net93),
    .CK(clknet_leaf_372_clk),
    .Q(\block_reg[0][22] ),
    .QN(_21940_));
 DFFR_X2 \block_reg[0][23]$_DFFE_PN0P_  (.D(_00454_),
    .RN(net91),
    .CK(clknet_leaf_286_clk),
    .Q(\block_reg[0][23] ),
    .QN(_21939_));
 DFFR_X2 \block_reg[0][24]$_DFFE_PN0P_  (.D(_00455_),
    .RN(net91),
    .CK(clknet_leaf_285_clk),
    .Q(\block_reg[0][24] ),
    .QN(_21938_));
 DFFR_X1 \block_reg[0][25]$_DFFE_PN0P_  (.D(_00456_),
    .RN(net93),
    .CK(clknet_leaf_372_clk),
    .Q(\block_reg[0][25] ),
    .QN(_21937_));
 DFFR_X2 \block_reg[0][26]$_DFFE_PN0P_  (.D(_00457_),
    .RN(net93),
    .CK(clknet_leaf_361_clk),
    .Q(\block_reg[0][26] ),
    .QN(_21936_));
 DFFR_X2 \block_reg[0][27]$_DFFE_PN0P_  (.D(_00458_),
    .RN(net93),
    .CK(clknet_leaf_363_clk),
    .Q(\block_reg[0][27] ),
    .QN(_21935_));
 DFFR_X2 \block_reg[0][28]$_DFFE_PN0P_  (.D(_00459_),
    .RN(net89),
    .CK(clknet_leaf_363_clk),
    .Q(\block_reg[0][28] ),
    .QN(_21934_));
 DFFR_X2 \block_reg[0][29]$_DFFE_PN0P_  (.D(_00460_),
    .RN(net91),
    .CK(clknet_leaf_288_clk),
    .Q(\block_reg[0][29] ),
    .QN(_21933_));
 DFFR_X2 \block_reg[0][2]$_DFFE_PN0P_  (.D(_00461_),
    .RN(net93),
    .CK(clknet_leaf_373_clk),
    .Q(\block_reg[0][2] ),
    .QN(_21932_));
 DFFR_X1 \block_reg[0][30]$_DFFE_PN0P_  (.D(_00462_),
    .RN(net93),
    .CK(clknet_leaf_363_clk),
    .Q(\block_reg[0][30] ),
    .QN(_21931_));
 DFFR_X2 \block_reg[0][31]$_DFFE_PN0P_  (.D(_00463_),
    .RN(net89),
    .CK(clknet_leaf_363_clk),
    .Q(\block_reg[0][31] ),
    .QN(_21930_));
 DFFR_X2 \block_reg[0][3]$_DFFE_PN0P_  (.D(_00464_),
    .RN(net89),
    .CK(clknet_leaf_372_clk),
    .Q(\block_reg[0][3] ),
    .QN(_21929_));
 DFFR_X1 \block_reg[0][4]$_DFFE_PN0P_  (.D(_00465_),
    .RN(net93),
    .CK(clknet_leaf_362_clk),
    .Q(\block_reg[0][4] ),
    .QN(_21928_));
 DFFR_X2 \block_reg[0][5]$_DFFE_PN0P_  (.D(_00466_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[0][5] ),
    .QN(_21927_));
 DFFR_X2 \block_reg[0][6]$_DFFE_PN0P_  (.D(_00467_),
    .RN(net91),
    .CK(clknet_leaf_285_clk),
    .Q(\block_reg[0][6] ),
    .QN(_21926_));
 DFFR_X2 \block_reg[0][7]$_DFFE_PN0P_  (.D(_00468_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[0][7] ),
    .QN(_21925_));
 DFFR_X2 \block_reg[0][8]$_DFFE_PN0P_  (.D(_00469_),
    .RN(net91),
    .CK(clknet_leaf_296_clk),
    .Q(\block_reg[0][8] ),
    .QN(_21924_));
 DFFR_X2 \block_reg[0][9]$_DFFE_PN0P_  (.D(_00470_),
    .RN(net90),
    .CK(clknet_leaf_293_clk),
    .Q(\block_reg[0][9] ),
    .QN(_21923_));
 DFFR_X2 \block_reg[1][0]$_DFFE_PN0P_  (.D(_00471_),
    .RN(net91),
    .CK(clknet_leaf_289_clk),
    .Q(\block_reg[1][0] ),
    .QN(_21922_));
 DFFR_X2 \block_reg[1][10]$_DFFE_PN0P_  (.D(_00472_),
    .RN(net91),
    .CK(clknet_leaf_290_clk),
    .Q(\block_reg[1][10] ),
    .QN(_21921_));
 DFFR_X2 \block_reg[1][11]$_DFFE_PN0P_  (.D(_00473_),
    .RN(net90),
    .CK(clknet_leaf_291_clk),
    .Q(\block_reg[1][11] ),
    .QN(_21920_));
 DFFR_X1 \block_reg[1][12]$_DFFE_PN0P_  (.D(_00474_),
    .RN(net90),
    .CK(clknet_leaf_291_clk),
    .Q(\block_reg[1][12] ),
    .QN(_21919_));
 DFFR_X2 \block_reg[1][13]$_DFFE_PN0P_  (.D(_00475_),
    .RN(net91),
    .CK(clknet_leaf_290_clk),
    .Q(\block_reg[1][13] ),
    .QN(_21918_));
 DFFR_X2 \block_reg[1][14]$_DFFE_PN0P_  (.D(_00476_),
    .RN(net91),
    .CK(clknet_leaf_292_clk),
    .Q(\block_reg[1][14] ),
    .QN(_21917_));
 DFFR_X2 \block_reg[1][15]$_DFFE_PN0P_  (.D(_00477_),
    .RN(net91),
    .CK(clknet_leaf_290_clk),
    .Q(\block_reg[1][15] ),
    .QN(_21916_));
 DFFR_X2 \block_reg[1][16]$_DFFE_PN0P_  (.D(_00478_),
    .RN(net90),
    .CK(clknet_leaf_297_clk),
    .Q(\block_reg[1][16] ),
    .QN(_21915_));
 DFFR_X1 \block_reg[1][17]$_DFFE_PN0P_  (.D(_00479_),
    .RN(net91),
    .CK(clknet_leaf_289_clk),
    .Q(\block_reg[1][17] ),
    .QN(_21914_));
 DFFR_X2 \block_reg[1][18]$_DFFE_PN0P_  (.D(_00480_),
    .RN(net91),
    .CK(clknet_leaf_289_clk),
    .Q(\block_reg[1][18] ),
    .QN(_21913_));
 DFFR_X2 \block_reg[1][19]$_DFFE_PN0P_  (.D(_00481_),
    .RN(net91),
    .CK(clknet_leaf_285_clk),
    .Q(\block_reg[1][19] ),
    .QN(_21912_));
 DFFR_X2 \block_reg[1][1]$_DFFE_PN0P_  (.D(_00482_),
    .RN(net91),
    .CK(clknet_leaf_292_clk),
    .Q(\block_reg[1][1] ),
    .QN(_21911_));
 DFFR_X2 \block_reg[1][20]$_DFFE_PN0P_  (.D(_00483_),
    .RN(net91),
    .CK(clknet_leaf_286_clk),
    .Q(\block_reg[1][20] ),
    .QN(_21910_));
 DFFR_X2 \block_reg[1][21]$_DFFE_PN0P_  (.D(_00484_),
    .RN(net93),
    .CK(clknet_leaf_362_clk),
    .Q(\block_reg[1][21] ),
    .QN(_21909_));
 DFFR_X2 \block_reg[1][22]$_DFFE_PN0P_  (.D(_00485_),
    .RN(net93),
    .CK(clknet_leaf_372_clk),
    .Q(\block_reg[1][22] ),
    .QN(_21908_));
 DFFR_X2 \block_reg[1][23]$_DFFE_PN0P_  (.D(_00486_),
    .RN(net91),
    .CK(clknet_leaf_286_clk),
    .Q(\block_reg[1][23] ),
    .QN(_21907_));
 DFFR_X1 \block_reg[1][24]$_DFFE_PN0P_  (.D(_00487_),
    .RN(net91),
    .CK(clknet_leaf_286_clk),
    .Q(\block_reg[1][24] ),
    .QN(_21906_));
 DFFR_X2 \block_reg[1][25]$_DFFE_PN0P_  (.D(_00488_),
    .RN(net93),
    .CK(clknet_leaf_372_clk),
    .Q(\block_reg[1][25] ),
    .QN(_21905_));
 DFFR_X2 \block_reg[1][26]$_DFFE_PN0P_  (.D(_00489_),
    .RN(net93),
    .CK(clknet_leaf_362_clk),
    .Q(\block_reg[1][26] ),
    .QN(_21904_));
 DFFR_X2 \block_reg[1][27]$_DFFE_PN0P_  (.D(_00490_),
    .RN(net93),
    .CK(clknet_leaf_362_clk),
    .Q(\block_reg[1][27] ),
    .QN(_21903_));
 DFFR_X2 \block_reg[1][28]$_DFFE_PN0P_  (.D(_00491_),
    .RN(net85),
    .CK(clknet_leaf_364_clk),
    .Q(\block_reg[1][28] ),
    .QN(_21902_));
 DFFR_X1 \block_reg[1][29]$_DFFE_PN0P_  (.D(_00492_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[1][29] ),
    .QN(_21901_));
 DFFR_X2 \block_reg[1][2]$_DFFE_PN0P_  (.D(_00493_),
    .RN(net93),
    .CK(clknet_leaf_373_clk),
    .Q(\block_reg[1][2] ),
    .QN(_21900_));
 DFFR_X2 \block_reg[1][30]$_DFFE_PN0P_  (.D(_00494_),
    .RN(net93),
    .CK(clknet_leaf_363_clk),
    .Q(\block_reg[1][30] ),
    .QN(_21899_));
 DFFR_X2 \block_reg[1][31]$_DFFE_PN0P_  (.D(_00495_),
    .RN(net85),
    .CK(clknet_leaf_363_clk),
    .Q(\block_reg[1][31] ),
    .QN(_21898_));
 DFFR_X2 \block_reg[1][3]$_DFFE_PN0P_  (.D(_00496_),
    .RN(net85),
    .CK(clknet_leaf_371_clk),
    .Q(\block_reg[1][3] ),
    .QN(_21897_));
 DFFR_X2 \block_reg[1][4]$_DFFE_PN0P_  (.D(_00497_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[1][4] ),
    .QN(_21896_));
 DFFR_X2 \block_reg[1][5]$_DFFE_PN0P_  (.D(_00498_),
    .RN(net91),
    .CK(clknet_leaf_288_clk),
    .Q(\block_reg[1][5] ),
    .QN(_21895_));
 DFFR_X2 \block_reg[1][6]$_DFFE_PN0P_  (.D(_00499_),
    .RN(net91),
    .CK(clknet_leaf_284_clk),
    .Q(\block_reg[1][6] ),
    .QN(_21894_));
 DFFR_X1 \block_reg[1][7]$_DFFE_PN0P_  (.D(_00500_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[1][7] ),
    .QN(_21893_));
 DFFR_X2 \block_reg[1][8]$_DFFE_PN0P_  (.D(_00501_),
    .RN(net91),
    .CK(clknet_leaf_296_clk),
    .Q(\block_reg[1][8] ),
    .QN(_21892_));
 DFFR_X2 \block_reg[1][9]$_DFFE_PN0P_  (.D(_00502_),
    .RN(net90),
    .CK(clknet_leaf_312_clk),
    .Q(\block_reg[1][9] ),
    .QN(_21891_));
 DFFR_X2 \block_reg[2][0]$_DFFE_PN0P_  (.D(_00503_),
    .RN(net91),
    .CK(clknet_leaf_291_clk),
    .Q(\block_reg[2][0] ),
    .QN(_21890_));
 DFFR_X1 \block_reg[2][10]$_DFFE_PN0P_  (.D(_00504_),
    .RN(net91),
    .CK(clknet_leaf_290_clk),
    .Q(\block_reg[2][10] ),
    .QN(_21889_));
 DFFR_X1 \block_reg[2][11]$_DFFE_PN0P_  (.D(_00505_),
    .RN(net91),
    .CK(clknet_leaf_271_clk),
    .Q(\block_reg[2][11] ),
    .QN(_21888_));
 DFFR_X2 \block_reg[2][12]$_DFFE_PN0P_  (.D(_00506_),
    .RN(net92),
    .CK(clknet_leaf_270_clk),
    .Q(\block_reg[2][12] ),
    .QN(_21887_));
 DFFR_X2 \block_reg[2][13]$_DFFE_PN0P_  (.D(_00507_),
    .RN(net92),
    .CK(clknet_leaf_271_clk),
    .Q(\block_reg[2][13] ),
    .QN(_21886_));
 DFFR_X2 \block_reg[2][14]$_DFFE_PN0P_  (.D(_00508_),
    .RN(net91),
    .CK(clknet_leaf_290_clk),
    .Q(\block_reg[2][14] ),
    .QN(_21885_));
 DFFR_X2 \block_reg[2][15]$_DFFE_PN0P_  (.D(_00509_),
    .RN(net92),
    .CK(clknet_leaf_271_clk),
    .Q(\block_reg[2][15] ),
    .QN(_21884_));
 DFFR_X2 \block_reg[2][16]$_DFFE_PN0P_  (.D(_00510_),
    .RN(net91),
    .CK(clknet_leaf_296_clk),
    .Q(\block_reg[2][16] ),
    .QN(_21883_));
 DFFR_X2 \block_reg[2][17]$_DFFE_PN0P_  (.D(_00511_),
    .RN(net91),
    .CK(clknet_leaf_292_clk),
    .Q(\block_reg[2][17] ),
    .QN(_21882_));
 DFFR_X2 \block_reg[2][18]$_DFFE_PN0P_  (.D(_00512_),
    .RN(net91),
    .CK(clknet_leaf_289_clk),
    .Q(\block_reg[2][18] ),
    .QN(_21881_));
 DFFR_X2 \block_reg[2][19]$_DFFE_PN0P_  (.D(_00513_),
    .RN(net93),
    .CK(clknet_leaf_363_clk),
    .Q(\block_reg[2][19] ),
    .QN(_21880_));
 DFFR_X1 \block_reg[2][1]$_DFFE_PN0P_  (.D(_00514_),
    .RN(net91),
    .CK(clknet_leaf_292_clk),
    .Q(\block_reg[2][1] ),
    .QN(_21879_));
 DFFR_X2 \block_reg[2][20]$_DFFE_PN0P_  (.D(_00515_),
    .RN(net93),
    .CK(clknet_leaf_362_clk),
    .Q(\block_reg[2][20] ),
    .QN(_21878_));
 DFFR_X2 \block_reg[2][21]$_DFFE_PN0P_  (.D(_00516_),
    .RN(net93),
    .CK(clknet_leaf_361_clk),
    .Q(\block_reg[2][21] ),
    .QN(_21877_));
 DFFR_X2 \block_reg[2][22]$_DFFE_PN0P_  (.D(_00517_),
    .RN(net93),
    .CK(clknet_leaf_364_clk),
    .Q(\block_reg[2][22] ),
    .QN(_21876_));
 DFFR_X1 \block_reg[2][23]$_DFFE_PN0P_  (.D(_00518_),
    .RN(net91),
    .CK(clknet_leaf_292_clk),
    .Q(\block_reg[2][23] ),
    .QN(_21875_));
 DFFR_X2 \block_reg[2][24]$_DFFE_PN0P_  (.D(_00519_),
    .RN(net91),
    .CK(clknet_leaf_286_clk),
    .Q(\block_reg[2][24] ),
    .QN(_21874_));
 DFFR_X2 \block_reg[2][25]$_DFFE_PN0P_  (.D(_00520_),
    .RN(net85),
    .CK(clknet_leaf_364_clk),
    .Q(\block_reg[2][25] ),
    .QN(_21873_));
 DFFR_X2 \block_reg[2][26]$_DFFE_PN0P_  (.D(_00521_),
    .RN(net85),
    .CK(clknet_leaf_361_clk),
    .Q(\block_reg[2][26] ),
    .QN(_21872_));
 DFFR_X2 \block_reg[2][27]$_DFFE_PN0P_  (.D(_00522_),
    .RN(net85),
    .CK(clknet_leaf_361_clk),
    .Q(\block_reg[2][27] ),
    .QN(_21871_));
 DFFR_X2 \block_reg[2][28]$_DFFE_PN0P_  (.D(_00523_),
    .RN(net85),
    .CK(clknet_leaf_364_clk),
    .Q(\block_reg[2][28] ),
    .QN(_21870_));
 DFFR_X2 \block_reg[2][29]$_DFFE_PN0P_  (.D(_00524_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[2][29] ),
    .QN(_21869_));
 DFFR_X2 \block_reg[2][2]$_DFFE_PN0P_  (.D(_00525_),
    .RN(net85),
    .CK(clknet_leaf_365_clk),
    .Q(\block_reg[2][2] ),
    .QN(_21868_));
 DFFR_X2 \block_reg[2][30]$_DFFE_PN0P_  (.D(_00526_),
    .RN(net85),
    .CK(clknet_leaf_365_clk),
    .Q(\block_reg[2][30] ),
    .QN(_21867_));
 DFFR_X2 \block_reg[2][31]$_DFFE_PN0P_  (.D(_00527_),
    .RN(net85),
    .CK(clknet_leaf_365_clk),
    .Q(\block_reg[2][31] ),
    .QN(_21866_));
 DFFR_X1 \block_reg[2][3]$_DFFE_PN0P_  (.D(_00528_),
    .RN(net85),
    .CK(clknet_leaf_364_clk),
    .Q(\block_reg[2][3] ),
    .QN(_21865_));
 DFFR_X2 \block_reg[2][4]$_DFFE_PN0P_  (.D(_00529_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[2][4] ),
    .QN(_21864_));
 DFFR_X2 \block_reg[2][5]$_DFFE_PN0P_  (.D(_00530_),
    .RN(net91),
    .CK(clknet_leaf_288_clk),
    .Q(\block_reg[2][5] ),
    .QN(_21863_));
 DFFR_X2 \block_reg[2][6]$_DFFE_PN0P_  (.D(_00531_),
    .RN(net91),
    .CK(clknet_leaf_285_clk),
    .Q(\block_reg[2][6] ),
    .QN(_21862_));
 DFFR_X1 \block_reg[2][7]$_DFFE_PN0P_  (.D(_00532_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[2][7] ),
    .QN(_21861_));
 DFFR_X1 \block_reg[2][8]$_DFFE_PN0P_  (.D(_00533_),
    .RN(net91),
    .CK(clknet_leaf_291_clk),
    .Q(\block_reg[2][8] ),
    .QN(_21860_));
 DFFR_X2 \block_reg[2][9]$_DFFE_PN0P_  (.D(_00534_),
    .RN(net90),
    .CK(clknet_leaf_311_clk),
    .Q(\block_reg[2][9] ),
    .QN(_21859_));
 DFFR_X2 \block_reg[3][0]$_DFFE_PN0P_  (.D(_00535_),
    .RN(net91),
    .CK(clknet_leaf_291_clk),
    .Q(\block_reg[3][0] ),
    .QN(_21858_));
 DFFR_X2 \block_reg[3][10]$_DFFE_PN0P_  (.D(_00536_),
    .RN(net91),
    .CK(clknet_leaf_290_clk),
    .Q(\block_reg[3][10] ),
    .QN(_21857_));
 DFFR_X2 \block_reg[3][11]$_DFFE_PN0P_  (.D(_00537_),
    .RN(net91),
    .CK(clknet_leaf_271_clk),
    .Q(\block_reg[3][11] ),
    .QN(_21856_));
 DFFR_X2 \block_reg[3][12]$_DFFE_PN0P_  (.D(_00538_),
    .RN(net91),
    .CK(clknet_leaf_297_clk),
    .Q(\block_reg[3][12] ),
    .QN(_21855_));
 DFFR_X2 \block_reg[3][13]$_DFFE_PN0P_  (.D(_00539_),
    .RN(net91),
    .CK(clknet_leaf_288_clk),
    .Q(\block_reg[3][13] ),
    .QN(_21854_));
 DFFR_X2 \block_reg[3][14]$_DFFE_PN0P_  (.D(_00540_),
    .RN(net91),
    .CK(clknet_leaf_289_clk),
    .Q(\block_reg[3][14] ),
    .QN(_21853_));
 DFFR_X2 \block_reg[3][15]$_DFFE_PN0P_  (.D(_00541_),
    .RN(net91),
    .CK(clknet_leaf_271_clk),
    .Q(\block_reg[3][15] ),
    .QN(_21852_));
 DFFR_X2 \block_reg[3][16]$_DFFE_PN0P_  (.D(_00542_),
    .RN(net91),
    .CK(clknet_leaf_296_clk),
    .Q(\block_reg[3][16] ),
    .QN(_21851_));
 DFFR_X2 \block_reg[3][17]$_DFFE_PN0P_  (.D(_00543_),
    .RN(net91),
    .CK(clknet_leaf_287_clk),
    .Q(\block_reg[3][17] ),
    .QN(_21850_));
 DFFR_X2 \block_reg[3][18]$_DFFE_PN0P_  (.D(_00544_),
    .RN(net91),
    .CK(clknet_leaf_289_clk),
    .Q(\block_reg[3][18] ),
    .QN(_21849_));
 DFFR_X2 \block_reg[3][19]$_DFFE_PN0P_  (.D(_00545_),
    .RN(net91),
    .CK(clknet_leaf_286_clk),
    .Q(\block_reg[3][19] ),
    .QN(_21848_));
 DFFR_X2 \block_reg[3][1]$_DFFE_PN0P_  (.D(_00546_),
    .RN(net91),
    .CK(clknet_leaf_286_clk),
    .Q(\block_reg[3][1] ),
    .QN(_21847_));
 DFFR_X1 \block_reg[3][20]$_DFFE_PN0P_  (.D(_00547_),
    .RN(net93),
    .CK(clknet_leaf_372_clk),
    .Q(\block_reg[3][20] ),
    .QN(_21846_));
 DFFR_X2 \block_reg[3][21]$_DFFE_PN0P_  (.D(_00548_),
    .RN(net93),
    .CK(clknet_leaf_363_clk),
    .Q(\block_reg[3][21] ),
    .QN(_21845_));
 DFFR_X2 \block_reg[3][22]$_DFFE_PN0P_  (.D(_00549_),
    .RN(net85),
    .CK(clknet_leaf_365_clk),
    .Q(\block_reg[3][22] ),
    .QN(_21844_));
 DFFR_X1 \block_reg[3][23]$_DFFE_PN0P_  (.D(_00550_),
    .RN(net85),
    .CK(clknet_leaf_361_clk),
    .Q(\block_reg[3][23] ),
    .QN(_21843_));
 DFFR_X1 \block_reg[3][24]$_DFFE_PN0P_  (.D(_00551_),
    .RN(net91),
    .CK(clknet_leaf_292_clk),
    .Q(\block_reg[3][24] ),
    .QN(_21842_));
 DFFR_X2 \block_reg[3][25]$_DFFE_PN0P_  (.D(_00552_),
    .RN(net85),
    .CK(clknet_leaf_365_clk),
    .Q(\block_reg[3][25] ),
    .QN(_21841_));
 DFFR_X2 \block_reg[3][26]$_DFFE_PN0P_  (.D(_00553_),
    .RN(net85),
    .CK(clknet_leaf_361_clk),
    .Q(\block_reg[3][26] ),
    .QN(_21840_));
 DFFR_X2 \block_reg[3][27]$_DFFE_PN0P_  (.D(_00554_),
    .RN(net85),
    .CK(clknet_leaf_365_clk),
    .Q(\block_reg[3][27] ),
    .QN(_21839_));
 DFFR_X2 \block_reg[3][28]$_DFFE_PN0P_  (.D(_00555_),
    .RN(net85),
    .CK(clknet_leaf_364_clk),
    .Q(\block_reg[3][28] ),
    .QN(_21838_));
 DFFR_X2 \block_reg[3][29]$_DFFE_PN0P_  (.D(_00556_),
    .RN(net85),
    .CK(clknet_leaf_365_clk),
    .Q(\block_reg[3][29] ),
    .QN(_21837_));
 DFFR_X2 \block_reg[3][2]$_DFFE_PN0P_  (.D(_00557_),
    .RN(net89),
    .CK(clknet_leaf_371_clk),
    .Q(\block_reg[3][2] ),
    .QN(_21836_));
 DFFR_X2 \block_reg[3][30]$_DFFE_PN0P_  (.D(_00558_),
    .RN(net85),
    .CK(clknet_leaf_365_clk),
    .Q(\block_reg[3][30] ),
    .QN(_21835_));
 DFFR_X2 \block_reg[3][31]$_DFFE_PN0P_  (.D(_00559_),
    .RN(net85),
    .CK(clknet_leaf_364_clk),
    .Q(\block_reg[3][31] ),
    .QN(_21834_));
 DFFR_X2 \block_reg[3][3]$_DFFE_PN0P_  (.D(_00560_),
    .RN(net89),
    .CK(clknet_leaf_371_clk),
    .Q(\block_reg[3][3] ),
    .QN(_21833_));
 DFFR_X2 \block_reg[3][4]$_DFFE_PN0P_  (.D(_00561_),
    .RN(net93),
    .CK(clknet_leaf_362_clk),
    .Q(\block_reg[3][4] ),
    .QN(_21832_));
 DFFR_X2 \block_reg[3][5]$_DFFE_PN0P_  (.D(_00562_),
    .RN(net89),
    .CK(clknet_leaf_371_clk),
    .Q(\block_reg[3][5] ),
    .QN(_21831_));
 DFFR_X2 \block_reg[3][6]$_DFFE_PN0P_  (.D(_00563_),
    .RN(net93),
    .CK(clknet_leaf_372_clk),
    .Q(\block_reg[3][6] ),
    .QN(_21830_));
 DFFR_X2 \block_reg[3][7]$_DFFE_PN0P_  (.D(_00564_),
    .RN(net89),
    .CK(clknet_leaf_371_clk),
    .Q(\block_reg[3][7] ),
    .QN(_21829_));
 DFFR_X1 \block_reg[3][8]$_DFFE_PN0P_  (.D(_00565_),
    .RN(net91),
    .CK(clknet_leaf_296_clk),
    .Q(\block_reg[3][8] ),
    .QN(_21828_));
 DFFR_X2 \block_reg[3][9]$_DFFE_PN0P_  (.D(_00566_),
    .RN(net90),
    .CK(clknet_leaf_312_clk),
    .Q(\block_reg[3][9] ),
    .QN(_21955_));
 DFFS_X2 \core.aes_core_ctrl_reg[0]$_DFF_PN1_  (.D(_00006_),
    .SN(net84),
    .CK(clknet_leaf_356_clk),
    .Q(\core.aes_core_ctrl_reg[0] ),
    .QN(_21956_));
 DFFR_X2 \core.aes_core_ctrl_reg[1]$_DFF_PN0_  (.D(_00007_),
    .RN(net84),
    .CK(clknet_leaf_356_clk),
    .Q(\core.aes_core_ctrl_reg[1] ),
    .QN(_21957_));
 DFFR_X1 \core.aes_core_ctrl_reg[2]$_DFF_PN0_  (.D(_00008_),
    .RN(net84),
    .CK(clknet_leaf_355_clk),
    .Q(\core.aes_core_ctrl_reg[2] ),
    .QN(_21827_));
 DFFR_X2 \core.dec_block.block_w0_reg[0]$_DFFE_PN0P_  (.D(_00567_),
    .RN(net91),
    .CK(clknet_leaf_302_clk),
    .Q(\core.dec_block.block_w0_reg[0] ),
    .QN(_21826_));
 DFFR_X2 \core.dec_block.block_w0_reg[10]$_DFFE_PN0P_  (.D(_00568_),
    .RN(net91),
    .CK(clknet_leaf_257_clk),
    .Q(\core.dec_block.block_w0_reg[10] ),
    .QN(_21825_));
 DFFR_X2 \core.dec_block.block_w0_reg[11]$_DFFE_PN0P_  (.D(_00569_),
    .RN(net91),
    .CK(clknet_leaf_257_clk),
    .Q(\core.dec_block.block_w0_reg[11] ),
    .QN(_21824_));
 DFFR_X2 \core.dec_block.block_w0_reg[12]$_DFFE_PN0P_  (.D(_00570_),
    .RN(net94),
    .CK(clknet_leaf_256_clk),
    .Q(\core.dec_block.block_w0_reg[12] ),
    .QN(_21823_));
 DFFR_X2 \core.dec_block.block_w0_reg[13]$_DFFE_PN0P_  (.D(_00571_),
    .RN(net92),
    .CK(clknet_leaf_259_clk),
    .Q(\core.dec_block.block_w0_reg[13] ),
    .QN(_21822_));
 DFFR_X1 \core.dec_block.block_w0_reg[14]$_DFFE_PN0P_  (.D(_00572_),
    .RN(net94),
    .CK(clknet_leaf_253_clk),
    .Q(\core.dec_block.block_w0_reg[14] ),
    .QN(_21821_));
 DFFR_X2 \core.dec_block.block_w0_reg[15]$_DFFE_PN0P_  (.D(_00573_),
    .RN(net94),
    .CK(clknet_leaf_253_clk),
    .Q(\core.dec_block.block_w0_reg[15] ),
    .QN(_21820_));
 DFFR_X2 \core.dec_block.block_w0_reg[16]$_DFFE_PN0P_  (.D(_00574_),
    .RN(net90),
    .CK(clknet_leaf_305_clk),
    .Q(\core.dec_block.block_w0_reg[16] ),
    .QN(_21819_));
 DFFR_X2 \core.dec_block.block_w0_reg[17]$_DFFE_PN0P_  (.D(_00575_),
    .RN(net90),
    .CK(clknet_leaf_306_clk),
    .Q(\core.dec_block.block_w0_reg[17] ),
    .QN(_21818_));
 DFFR_X2 \core.dec_block.block_w0_reg[18]$_DFFE_PN0P_  (.D(_00576_),
    .RN(net90),
    .CK(clknet_leaf_304_clk),
    .Q(\core.dec_block.block_w0_reg[18] ),
    .QN(_21817_));
 DFFR_X1 \core.dec_block.block_w0_reg[19]$_DFFE_PN0P_  (.D(_00577_),
    .RN(net90),
    .CK(clknet_leaf_306_clk),
    .Q(\core.dec_block.block_w0_reg[19] ),
    .QN(_21816_));
 DFFR_X2 \core.dec_block.block_w0_reg[1]$_DFFE_PN0P_  (.D(_00578_),
    .RN(net90),
    .CK(clknet_leaf_300_clk),
    .Q(\core.dec_block.block_w0_reg[1] ),
    .QN(_21815_));
 DFFR_X2 \core.dec_block.block_w0_reg[20]$_DFFE_PN0P_  (.D(_00579_),
    .RN(net90),
    .CK(clknet_leaf_305_clk),
    .Q(\core.dec_block.block_w0_reg[20] ),
    .QN(_21814_));
 DFFR_X2 \core.dec_block.block_w0_reg[21]$_DFFE_PN0P_  (.D(_00580_),
    .RN(net90),
    .CK(clknet_leaf_310_clk),
    .Q(\core.dec_block.block_w0_reg[21] ),
    .QN(_21813_));
 DFFR_X2 \core.dec_block.block_w0_reg[22]$_DFFE_PN0P_  (.D(_00581_),
    .RN(net90),
    .CK(clknet_leaf_305_clk),
    .Q(\core.dec_block.block_w0_reg[22] ),
    .QN(_21812_));
 DFFR_X1 \core.dec_block.block_w0_reg[23]$_DFFE_PN0P_  (.D(_00582_),
    .RN(net91),
    .CK(clknet_leaf_255_clk),
    .Q(\core.dec_block.block_w0_reg[23] ),
    .QN(_21811_));
 DFFR_X2 \core.dec_block.block_w0_reg[24]$_DFFE_PN0P_  (.D(_00583_),
    .RN(net90),
    .CK(clknet_leaf_298_clk),
    .Q(\core.dec_block.block_w0_reg[24] ),
    .QN(_21810_));
 DFFR_X2 \core.dec_block.block_w0_reg[25]$_DFFE_PN0P_  (.D(_00584_),
    .RN(net90),
    .CK(clknet_leaf_295_clk),
    .Q(\core.dec_block.block_w0_reg[25] ),
    .QN(_21809_));
 DFFR_X2 \core.dec_block.block_w0_reg[26]$_DFFE_PN0P_  (.D(_00585_),
    .RN(net90),
    .CK(clknet_leaf_311_clk),
    .Q(\core.dec_block.block_w0_reg[26] ),
    .QN(_21808_));
 DFFR_X2 \core.dec_block.block_w0_reg[27]$_DFFE_PN0P_  (.D(_00586_),
    .RN(net90),
    .CK(clknet_leaf_295_clk),
    .Q(\core.dec_block.block_w0_reg[27] ),
    .QN(_21807_));
 DFFR_X2 \core.dec_block.block_w0_reg[28]$_DFFE_PN0P_  (.D(_00587_),
    .RN(net90),
    .CK(clknet_leaf_311_clk),
    .Q(\core.dec_block.block_w0_reg[28] ),
    .QN(_21806_));
 DFFR_X2 \core.dec_block.block_w0_reg[29]$_DFFE_PN0P_  (.D(_00588_),
    .RN(net90),
    .CK(clknet_leaf_299_clk),
    .Q(\core.dec_block.block_w0_reg[29] ),
    .QN(_21805_));
 DFFR_X2 \core.dec_block.block_w0_reg[2]$_DFFE_PN0P_  (.D(_00589_),
    .RN(net90),
    .CK(clknet_leaf_294_clk),
    .Q(\core.dec_block.block_w0_reg[2] ),
    .QN(_21804_));
 DFFR_X2 \core.dec_block.block_w0_reg[30]$_DFFE_PN0P_  (.D(_00590_),
    .RN(net91),
    .CK(clknet_leaf_255_clk),
    .Q(\core.dec_block.block_w0_reg[30] ),
    .QN(_21803_));
 DFFR_X1 \core.dec_block.block_w0_reg[31]$_DFFE_PN0P_  (.D(_00591_),
    .RN(net90),
    .CK(clknet_leaf_299_clk),
    .Q(\core.dec_block.block_w0_reg[31] ),
    .QN(_21802_));
 DFFR_X2 \core.dec_block.block_w0_reg[3]$_DFFE_PN0P_  (.D(_00592_),
    .RN(net90),
    .CK(clknet_leaf_294_clk),
    .Q(\core.dec_block.block_w0_reg[3] ),
    .QN(_21801_));
 DFFR_X2 \core.dec_block.block_w0_reg[4]$_DFFE_PN0P_  (.D(_00593_),
    .RN(net91),
    .CK(clknet_leaf_255_clk),
    .Q(\core.dec_block.block_w0_reg[4] ),
    .QN(_21800_));
 DFFR_X2 \core.dec_block.block_w0_reg[5]$_DFFE_PN0P_  (.D(_00594_),
    .RN(net91),
    .CK(clknet_leaf_298_clk),
    .Q(\core.dec_block.block_w0_reg[5] ),
    .QN(_21799_));
 DFFR_X2 \core.dec_block.block_w0_reg[6]$_DFFE_PN0P_  (.D(_00595_),
    .RN(net91),
    .CK(clknet_leaf_298_clk),
    .Q(\core.dec_block.block_w0_reg[6] ),
    .QN(_21798_));
 DFFR_X1 \core.dec_block.block_w0_reg[7]$_DFFE_PN0P_  (.D(_00596_),
    .RN(net91),
    .CK(clknet_leaf_257_clk),
    .Q(\core.dec_block.block_w0_reg[7] ),
    .QN(_21797_));
 DFFR_X2 \core.dec_block.block_w0_reg[8]$_DFFE_PN0P_  (.D(_00597_),
    .RN(net91),
    .CK(clknet_leaf_257_clk),
    .Q(\core.dec_block.block_w0_reg[8] ),
    .QN(_21796_));
 DFFR_X2 \core.dec_block.block_w0_reg[9]$_DFFE_PN0P_  (.D(_00598_),
    .RN(net91),
    .CK(clknet_leaf_256_clk),
    .Q(\core.dec_block.block_w0_reg[9] ),
    .QN(_21795_));
 DFFR_X2 \core.dec_block.block_w1_reg[0]$_DFFE_PN0P_  (.D(_00599_),
    .RN(net91),
    .CK(clknet_leaf_302_clk),
    .Q(\core.dec_block.block_w1_reg[0] ),
    .QN(_21794_));
 DFFR_X2 \core.dec_block.block_w1_reg[10]$_DFFE_PN0P_  (.D(_00600_),
    .RN(net91),
    .CK(clknet_leaf_303_clk),
    .Q(\core.dec_block.block_w1_reg[10] ),
    .QN(_21793_));
 DFFR_X2 \core.dec_block.block_w1_reg[11]$_DFFE_PN0P_  (.D(_00601_),
    .RN(net91),
    .CK(clknet_leaf_253_clk),
    .Q(\core.dec_block.block_w1_reg[11] ),
    .QN(_21792_));
 DFFR_X2 \core.dec_block.block_w1_reg[12]$_DFFE_PN0P_  (.D(_00602_),
    .RN(net91),
    .CK(clknet_leaf_255_clk),
    .Q(\core.dec_block.block_w1_reg[12] ),
    .QN(_21791_));
 DFFR_X2 \core.dec_block.block_w1_reg[13]$_DFFE_PN0P_  (.D(_00603_),
    .RN(net91),
    .CK(clknet_leaf_253_clk),
    .Q(\core.dec_block.block_w1_reg[13] ),
    .QN(_21790_));
 DFFR_X2 \core.dec_block.block_w1_reg[14]$_DFFE_PN0P_  (.D(_00604_),
    .RN(net91),
    .CK(clknet_leaf_254_clk),
    .Q(\core.dec_block.block_w1_reg[14] ),
    .QN(_21789_));
 DFFR_X2 \core.dec_block.block_w1_reg[15]$_DFFE_PN0P_  (.D(_00605_),
    .RN(net91),
    .CK(clknet_leaf_253_clk),
    .Q(\core.dec_block.block_w1_reg[15] ),
    .QN(_21788_));
 DFFR_X2 \core.dec_block.block_w1_reg[16]$_DFFE_PN0P_  (.D(_00606_),
    .RN(net91),
    .CK(clknet_leaf_303_clk),
    .Q(\core.dec_block.block_w1_reg[16] ),
    .QN(_21787_));
 DFFR_X2 \core.dec_block.block_w1_reg[17]$_DFFE_PN0P_  (.D(_00607_),
    .RN(net91),
    .CK(clknet_leaf_301_clk),
    .Q(\core.dec_block.block_w1_reg[17] ),
    .QN(_21786_));
 DFFR_X2 \core.dec_block.block_w1_reg[18]$_DFFE_PN0P_  (.D(_00608_),
    .RN(net91),
    .CK(clknet_leaf_303_clk),
    .Q(\core.dec_block.block_w1_reg[18] ),
    .QN(_21785_));
 DFFR_X2 \core.dec_block.block_w1_reg[19]$_DFFE_PN0P_  (.D(_00609_),
    .RN(net90),
    .CK(clknet_leaf_301_clk),
    .Q(\core.dec_block.block_w1_reg[19] ),
    .QN(_21784_));
 DFFR_X2 \core.dec_block.block_w1_reg[1]$_DFFE_PN0P_  (.D(_00610_),
    .RN(net90),
    .CK(clknet_leaf_300_clk),
    .Q(\core.dec_block.block_w1_reg[1] ),
    .QN(_21783_));
 DFFR_X2 \core.dec_block.block_w1_reg[20]$_DFFE_PN0P_  (.D(_00611_),
    .RN(net91),
    .CK(clknet_leaf_302_clk),
    .Q(\core.dec_block.block_w1_reg[20] ),
    .QN(_21782_));
 DFFR_X2 \core.dec_block.block_w1_reg[21]$_DFFE_PN0P_  (.D(_00612_),
    .RN(net90),
    .CK(clknet_leaf_305_clk),
    .Q(\core.dec_block.block_w1_reg[21] ),
    .QN(_21781_));
 DFFR_X2 \core.dec_block.block_w1_reg[22]$_DFFE_PN0P_  (.D(_00613_),
    .RN(net91),
    .CK(clknet_leaf_301_clk),
    .Q(\core.dec_block.block_w1_reg[22] ),
    .QN(_21780_));
 DFFR_X1 \core.dec_block.block_w1_reg[23]$_DFFE_PN0P_  (.D(_00614_),
    .RN(net91),
    .CK(clknet_leaf_255_clk),
    .Q(\core.dec_block.block_w1_reg[23] ),
    .QN(_21779_));
 DFFR_X2 \core.dec_block.block_w1_reg[24]$_DFFE_PN0P_  (.D(_00615_),
    .RN(net91),
    .CK(clknet_leaf_304_clk),
    .Q(\core.dec_block.block_w1_reg[24] ),
    .QN(_21778_));
 DFFR_X2 \core.dec_block.block_w1_reg[25]$_DFFE_PN0P_  (.D(_00616_),
    .RN(net90),
    .CK(clknet_leaf_304_clk),
    .Q(\core.dec_block.block_w1_reg[25] ),
    .QN(_21777_));
 DFFR_X2 \core.dec_block.block_w1_reg[26]$_DFFE_PN0P_  (.D(_00617_),
    .RN(net91),
    .CK(clknet_leaf_303_clk),
    .Q(\core.dec_block.block_w1_reg[26] ),
    .QN(_21776_));
 DFFR_X2 \core.dec_block.block_w1_reg[27]$_DFFE_PN0P_  (.D(_00618_),
    .RN(net90),
    .CK(clknet_leaf_306_clk),
    .Q(\core.dec_block.block_w1_reg[27] ),
    .QN(_21775_));
 DFFR_X2 \core.dec_block.block_w1_reg[28]$_DFFE_PN0P_  (.D(_00619_),
    .RN(net90),
    .CK(clknet_leaf_304_clk),
    .Q(\core.dec_block.block_w1_reg[28] ),
    .QN(_21774_));
 DFFR_X2 \core.dec_block.block_w1_reg[29]$_DFFE_PN0P_  (.D(_00620_),
    .RN(net90),
    .CK(clknet_leaf_301_clk),
    .Q(\core.dec_block.block_w1_reg[29] ),
    .QN(_21773_));
 DFFR_X2 \core.dec_block.block_w1_reg[2]$_DFFE_PN0P_  (.D(_00621_),
    .RN(net90),
    .CK(clknet_leaf_294_clk),
    .Q(\core.dec_block.block_w1_reg[2] ),
    .QN(_21772_));
 DFFR_X2 \core.dec_block.block_w1_reg[30]$_DFFE_PN0P_  (.D(_00622_),
    .RN(net91),
    .CK(clknet_leaf_302_clk),
    .Q(\core.dec_block.block_w1_reg[30] ),
    .QN(_21771_));
 DFFR_X2 \core.dec_block.block_w1_reg[31]$_DFFE_PN0P_  (.D(_00623_),
    .RN(net91),
    .CK(clknet_leaf_303_clk),
    .Q(\core.dec_block.block_w1_reg[31] ),
    .QN(_21770_));
 DFFR_X2 \core.dec_block.block_w1_reg[3]$_DFFE_PN0P_  (.D(_00624_),
    .RN(net90),
    .CK(clknet_leaf_294_clk),
    .Q(\core.dec_block.block_w1_reg[3] ),
    .QN(_21769_));
 DFFR_X2 \core.dec_block.block_w1_reg[4]$_DFFE_PN0P_  (.D(_00625_),
    .RN(net91),
    .CK(clknet_leaf_256_clk),
    .Q(\core.dec_block.block_w1_reg[4] ),
    .QN(_21768_));
 DFFR_X2 \core.dec_block.block_w1_reg[5]$_DFFE_PN0P_  (.D(_00626_),
    .RN(net91),
    .CK(clknet_leaf_299_clk),
    .Q(\core.dec_block.block_w1_reg[5] ),
    .QN(_21767_));
 DFFR_X2 \core.dec_block.block_w1_reg[6]$_DFFE_PN0P_  (.D(_00627_),
    .RN(net91),
    .CK(clknet_leaf_299_clk),
    .Q(\core.dec_block.block_w1_reg[6] ),
    .QN(_21766_));
 DFFR_X2 \core.dec_block.block_w1_reg[7]$_DFFE_PN0P_  (.D(_00628_),
    .RN(net90),
    .CK(clknet_leaf_299_clk),
    .Q(\core.dec_block.block_w1_reg[7] ),
    .QN(_21765_));
 DFFR_X2 \core.dec_block.block_w1_reg[8]$_DFFE_PN0P_  (.D(_00629_),
    .RN(net90),
    .CK(clknet_leaf_299_clk),
    .Q(\core.dec_block.block_w1_reg[8] ),
    .QN(_21764_));
 DFFR_X2 \core.dec_block.block_w1_reg[9]$_DFFE_PN0P_  (.D(_00630_),
    .RN(net91),
    .CK(clknet_leaf_302_clk),
    .Q(\core.dec_block.block_w1_reg[9] ),
    .QN(_21763_));
 DFFR_X2 \core.dec_block.block_w2_reg[0]$_DFFE_PN0P_  (.D(_00631_),
    .RN(net90),
    .CK(clknet_leaf_301_clk),
    .Q(\core.dec_block.block_w2_reg[0] ),
    .QN(_21762_));
 DFFR_X2 \core.dec_block.block_w2_reg[10]$_DFFE_PN0P_  (.D(_00632_),
    .RN(net91),
    .CK(clknet_leaf_257_clk),
    .Q(\core.dec_block.block_w2_reg[10] ),
    .QN(_21761_));
 DFFR_X2 \core.dec_block.block_w2_reg[11]$_DFFE_PN0P_  (.D(_00633_),
    .RN(net91),
    .CK(clknet_leaf_257_clk),
    .Q(\core.dec_block.block_w2_reg[11] ),
    .QN(_21760_));
 DFFR_X2 \core.dec_block.block_w2_reg[12]$_DFFE_PN0P_  (.D(_00634_),
    .RN(net94),
    .CK(clknet_leaf_256_clk),
    .Q(\core.dec_block.block_w2_reg[12] ),
    .QN(_21759_));
 DFFR_X2 \core.dec_block.block_w2_reg[13]$_DFFE_PN0P_  (.D(_00635_),
    .RN(net91),
    .CK(clknet_leaf_256_clk),
    .Q(\core.dec_block.block_w2_reg[13] ),
    .QN(_21758_));
 DFFR_X2 \core.dec_block.block_w2_reg[14]$_DFFE_PN0P_  (.D(_00636_),
    .RN(net91),
    .CK(clknet_leaf_254_clk),
    .Q(\core.dec_block.block_w2_reg[14] ),
    .QN(_21757_));
 DFFR_X2 \core.dec_block.block_w2_reg[15]$_DFFE_PN0P_  (.D(_00637_),
    .RN(net91),
    .CK(clknet_leaf_254_clk),
    .Q(\core.dec_block.block_w2_reg[15] ),
    .QN(_21756_));
 DFFR_X2 \core.dec_block.block_w2_reg[16]$_DFFE_PN0P_  (.D(_00638_),
    .RN(net91),
    .CK(clknet_leaf_303_clk),
    .Q(\core.dec_block.block_w2_reg[16] ),
    .QN(_21755_));
 DFFR_X2 \core.dec_block.block_w2_reg[17]$_DFFE_PN0P_  (.D(_00639_),
    .RN(net91),
    .CK(clknet_leaf_304_clk),
    .Q(\core.dec_block.block_w2_reg[17] ),
    .QN(_21754_));
 DFFR_X2 \core.dec_block.block_w2_reg[18]$_DFFE_PN0P_  (.D(_00640_),
    .RN(net91),
    .CK(clknet_leaf_304_clk),
    .Q(\core.dec_block.block_w2_reg[18] ),
    .QN(_21753_));
 DFFR_X2 \core.dec_block.block_w2_reg[19]$_DFFE_PN0P_  (.D(_00641_),
    .RN(net90),
    .CK(clknet_leaf_305_clk),
    .Q(\core.dec_block.block_w2_reg[19] ),
    .QN(_21752_));
 DFFR_X2 \core.dec_block.block_w2_reg[1]$_DFFE_PN0P_  (.D(_00642_),
    .RN(net90),
    .CK(clknet_leaf_294_clk),
    .Q(\core.dec_block.block_w2_reg[1] ),
    .QN(_21751_));
 DFFR_X2 \core.dec_block.block_w2_reg[20]$_DFFE_PN0P_  (.D(_00643_),
    .RN(net91),
    .CK(clknet_leaf_303_clk),
    .Q(\core.dec_block.block_w2_reg[20] ),
    .QN(_21750_));
 DFFR_X2 \core.dec_block.block_w2_reg[21]$_DFFE_PN0P_  (.D(_00644_),
    .RN(net91),
    .CK(clknet_leaf_301_clk),
    .Q(\core.dec_block.block_w2_reg[21] ),
    .QN(_21749_));
 DFFR_X2 \core.dec_block.block_w2_reg[22]$_DFFE_PN0P_  (.D(_00645_),
    .RN(net90),
    .CK(clknet_leaf_301_clk),
    .Q(\core.dec_block.block_w2_reg[22] ),
    .QN(_21748_));
 DFFR_X1 \core.dec_block.block_w2_reg[23]$_DFFE_PN0P_  (.D(_00646_),
    .RN(net91),
    .CK(clknet_leaf_255_clk),
    .Q(\core.dec_block.block_w2_reg[23] ),
    .QN(_21747_));
 DFFR_X2 \core.dec_block.block_w2_reg[24]$_DFFE_PN0P_  (.D(_00647_),
    .RN(net90),
    .CK(clknet_leaf_295_clk),
    .Q(\core.dec_block.block_w2_reg[24] ),
    .QN(_21746_));
 DFFR_X2 \core.dec_block.block_w2_reg[25]$_DFFE_PN0P_  (.D(_00648_),
    .RN(net90),
    .CK(clknet_leaf_295_clk),
    .Q(\core.dec_block.block_w2_reg[25] ),
    .QN(_21745_));
 DFFR_X2 \core.dec_block.block_w2_reg[26]$_DFFE_PN0P_  (.D(_00649_),
    .RN(net90),
    .CK(clknet_leaf_295_clk),
    .Q(\core.dec_block.block_w2_reg[26] ),
    .QN(_21744_));
 DFFR_X2 \core.dec_block.block_w2_reg[27]$_DFFE_PN0P_  (.D(_00650_),
    .RN(net90),
    .CK(clknet_leaf_295_clk),
    .Q(\core.dec_block.block_w2_reg[27] ),
    .QN(_21743_));
 DFFR_X2 \core.dec_block.block_w2_reg[28]$_DFFE_PN0P_  (.D(_00651_),
    .RN(net90),
    .CK(clknet_leaf_293_clk),
    .Q(\core.dec_block.block_w2_reg[28] ),
    .QN(_21742_));
 DFFR_X2 \core.dec_block.block_w2_reg[29]$_DFFE_PN0P_  (.D(_00652_),
    .RN(net90),
    .CK(clknet_leaf_298_clk),
    .Q(\core.dec_block.block_w2_reg[29] ),
    .QN(_21741_));
 DFFR_X2 \core.dec_block.block_w2_reg[2]$_DFFE_PN0P_  (.D(_00653_),
    .RN(net90),
    .CK(clknet_leaf_293_clk),
    .Q(\core.dec_block.block_w2_reg[2] ),
    .QN(_21740_));
 DFFR_X2 \core.dec_block.block_w2_reg[30]$_DFFE_PN0P_  (.D(_00654_),
    .RN(net91),
    .CK(clknet_leaf_297_clk),
    .Q(\core.dec_block.block_w2_reg[30] ),
    .QN(_21739_));
 DFFR_X2 \core.dec_block.block_w2_reg[31]$_DFFE_PN0P_  (.D(_00655_),
    .RN(net90),
    .CK(clknet_leaf_297_clk),
    .Q(\core.dec_block.block_w2_reg[31] ),
    .QN(_21738_));
 DFFR_X2 \core.dec_block.block_w2_reg[3]$_DFFE_PN0P_  (.D(_00656_),
    .RN(net90),
    .CK(clknet_leaf_293_clk),
    .Q(\core.dec_block.block_w2_reg[3] ),
    .QN(_21737_));
 DFFR_X2 \core.dec_block.block_w2_reg[4]$_DFFE_PN0P_  (.D(_00657_),
    .RN(net90),
    .CK(clknet_leaf_311_clk),
    .Q(\core.dec_block.block_w2_reg[4] ),
    .QN(_21736_));
 DFFR_X2 \core.dec_block.block_w2_reg[5]$_DFFE_PN0P_  (.D(_00658_),
    .RN(net90),
    .CK(clknet_leaf_294_clk),
    .Q(\core.dec_block.block_w2_reg[5] ),
    .QN(_21735_));
 DFFR_X1 \core.dec_block.block_w2_reg[6]$_DFFE_PN0P_  (.D(_00659_),
    .RN(net90),
    .CK(clknet_leaf_294_clk),
    .Q(\core.dec_block.block_w2_reg[6] ),
    .QN(_21734_));
 DFFR_X2 \core.dec_block.block_w2_reg[7]$_DFFE_PN0P_  (.D(_00660_),
    .RN(net90),
    .CK(clknet_leaf_300_clk),
    .Q(\core.dec_block.block_w2_reg[7] ),
    .QN(_21733_));
 DFFR_X2 \core.dec_block.block_w2_reg[8]$_DFFE_PN0P_  (.D(_00661_),
    .RN(net90),
    .CK(clknet_leaf_298_clk),
    .Q(\core.dec_block.block_w2_reg[8] ),
    .QN(_21732_));
 DFFR_X2 \core.dec_block.block_w2_reg[9]$_DFFE_PN0P_  (.D(_00662_),
    .RN(net91),
    .CK(clknet_leaf_298_clk),
    .Q(\core.dec_block.block_w2_reg[9] ),
    .QN(_21731_));
 DFFR_X2 \core.dec_block.block_w3_reg[0]$_DFFE_PN0P_  (.D(_00663_),
    .RN(net90),
    .CK(clknet_leaf_300_clk),
    .Q(\core.dec_block.block_w3_reg[0] ),
    .QN(_21730_));
 DFFR_X2 \core.dec_block.block_w3_reg[10]$_DFFE_PN0P_  (.D(_00664_),
    .RN(net91),
    .CK(clknet_leaf_302_clk),
    .Q(\core.dec_block.block_w3_reg[10] ),
    .QN(_21729_));
 DFFR_X1 \core.dec_block.block_w3_reg[11]$_DFFE_PN0P_  (.D(_00665_),
    .RN(net91),
    .CK(clknet_leaf_254_clk),
    .Q(\core.dec_block.block_w3_reg[11] ),
    .QN(_21728_));
 DFFR_X2 \core.dec_block.block_w3_reg[12]$_DFFE_PN0P_  (.D(_00666_),
    .RN(net91),
    .CK(clknet_leaf_254_clk),
    .Q(\core.dec_block.block_w3_reg[12] ),
    .QN(_21727_));
 DFFR_X2 \core.dec_block.block_w3_reg[13]$_DFFE_PN0P_  (.D(_00667_),
    .RN(net91),
    .CK(clknet_leaf_255_clk),
    .Q(\core.dec_block.block_w3_reg[13] ),
    .QN(_21726_));
 DFFR_X1 \core.dec_block.block_w3_reg[14]$_DFFE_PN0P_  (.D(_00668_),
    .RN(net91),
    .CK(clknet_leaf_254_clk),
    .Q(\core.dec_block.block_w3_reg[14] ),
    .QN(_21725_));
 DFFR_X2 \core.dec_block.block_w3_reg[15]$_DFFE_PN0P_  (.D(_00669_),
    .RN(net91),
    .CK(clknet_leaf_253_clk),
    .Q(\core.dec_block.block_w3_reg[15] ),
    .QN(_21724_));
 DFFR_X2 \core.dec_block.block_w3_reg[16]$_DFFE_PN0P_  (.D(_00670_),
    .RN(net90),
    .CK(clknet_leaf_305_clk),
    .Q(\core.dec_block.block_w3_reg[16] ),
    .QN(_21723_));
 DFFR_X2 \core.dec_block.block_w3_reg[17]$_DFFE_PN0P_  (.D(_00671_),
    .RN(net90),
    .CK(clknet_leaf_305_clk),
    .Q(\core.dec_block.block_w3_reg[17] ),
    .QN(_21722_));
 DFFR_X2 \core.dec_block.block_w3_reg[18]$_DFFE_PN0P_  (.D(_00672_),
    .RN(net90),
    .CK(clknet_leaf_305_clk),
    .Q(\core.dec_block.block_w3_reg[18] ),
    .QN(_21721_));
 DFFR_X2 \core.dec_block.block_w3_reg[19]$_DFFE_PN0P_  (.D(_00673_),
    .RN(net90),
    .CK(clknet_leaf_307_clk),
    .Q(\core.dec_block.block_w3_reg[19] ),
    .QN(_21720_));
 DFFR_X2 \core.dec_block.block_w3_reg[1]$_DFFE_PN0P_  (.D(_00674_),
    .RN(net90),
    .CK(clknet_leaf_310_clk),
    .Q(\core.dec_block.block_w3_reg[1] ),
    .QN(_21719_));
 DFFR_X2 \core.dec_block.block_w3_reg[20]$_DFFE_PN0P_  (.D(_00675_),
    .RN(net90),
    .CK(clknet_leaf_306_clk),
    .Q(\core.dec_block.block_w3_reg[20] ),
    .QN(_21718_));
 DFFR_X2 \core.dec_block.block_w3_reg[21]$_DFFE_PN0P_  (.D(_00676_),
    .RN(net90),
    .CK(clknet_leaf_310_clk),
    .Q(\core.dec_block.block_w3_reg[21] ),
    .QN(_21717_));
 DFFR_X2 \core.dec_block.block_w3_reg[22]$_DFFE_PN0P_  (.D(_00677_),
    .RN(net90),
    .CK(clknet_leaf_310_clk),
    .Q(\core.dec_block.block_w3_reg[22] ),
    .QN(_21716_));
 DFFR_X1 \core.dec_block.block_w3_reg[23]$_DFFE_PN0P_  (.D(_00678_),
    .RN(net90),
    .CK(clknet_leaf_306_clk),
    .Q(\core.dec_block.block_w3_reg[23] ),
    .QN(_21715_));
 DFFR_X2 \core.dec_block.block_w3_reg[24]$_DFFE_PN0P_  (.D(_00679_),
    .RN(net90),
    .CK(clknet_leaf_306_clk),
    .Q(\core.dec_block.block_w3_reg[24] ),
    .QN(_21714_));
 DFFR_X2 \core.dec_block.block_w3_reg[25]$_DFFE_PN0P_  (.D(_00680_),
    .RN(net90),
    .CK(clknet_leaf_308_clk),
    .Q(\core.dec_block.block_w3_reg[25] ),
    .QN(_21713_));
 DFFR_X2 \core.dec_block.block_w3_reg[26]$_DFFE_PN0P_  (.D(_00681_),
    .RN(net90),
    .CK(clknet_leaf_310_clk),
    .Q(\core.dec_block.block_w3_reg[26] ),
    .QN(_21712_));
 DFFR_X2 \core.dec_block.block_w3_reg[27]$_DFFE_PN0P_  (.D(_00682_),
    .RN(net90),
    .CK(clknet_leaf_311_clk),
    .Q(\core.dec_block.block_w3_reg[27] ),
    .QN(_21711_));
 DFFR_X2 \core.dec_block.block_w3_reg[28]$_DFFE_PN0P_  (.D(_00683_),
    .RN(net90),
    .CK(clknet_leaf_308_clk),
    .Q(\core.dec_block.block_w3_reg[28] ),
    .QN(_21710_));
 DFFR_X2 \core.dec_block.block_w3_reg[29]$_DFFE_PN0P_  (.D(_00684_),
    .RN(net90),
    .CK(clknet_leaf_309_clk),
    .Q(\core.dec_block.block_w3_reg[29] ),
    .QN(_21709_));
 DFFR_X2 \core.dec_block.block_w3_reg[2]$_DFFE_PN0P_  (.D(_00685_),
    .RN(net90),
    .CK(clknet_leaf_306_clk),
    .Q(\core.dec_block.block_w3_reg[2] ),
    .QN(_21708_));
 DFFR_X2 \core.dec_block.block_w3_reg[30]$_DFFE_PN0P_  (.D(_00686_),
    .RN(net90),
    .CK(clknet_leaf_309_clk),
    .Q(\core.dec_block.block_w3_reg[30] ),
    .QN(_21707_));
 DFFR_X2 \core.dec_block.block_w3_reg[31]$_DFFE_PN0P_  (.D(_00687_),
    .RN(net90),
    .CK(clknet_leaf_309_clk),
    .Q(\core.dec_block.block_w3_reg[31] ),
    .QN(_21706_));
 DFFR_X2 \core.dec_block.block_w3_reg[3]$_DFFE_PN0P_  (.D(_00688_),
    .RN(net90),
    .CK(clknet_leaf_311_clk),
    .Q(\core.dec_block.block_w3_reg[3] ),
    .QN(_21705_));
 DFFR_X2 \core.dec_block.block_w3_reg[4]$_DFFE_PN0P_  (.D(_00689_),
    .RN(net90),
    .CK(clknet_leaf_310_clk),
    .Q(\core.dec_block.block_w3_reg[4] ),
    .QN(_21704_));
 DFFR_X2 \core.dec_block.block_w3_reg[5]$_DFFE_PN0P_  (.D(_00690_),
    .RN(net90),
    .CK(clknet_leaf_300_clk),
    .Q(\core.dec_block.block_w3_reg[5] ),
    .QN(_21703_));
 DFFR_X2 \core.dec_block.block_w3_reg[6]$_DFFE_PN0P_  (.D(_00691_),
    .RN(net90),
    .CK(clknet_leaf_311_clk),
    .Q(\core.dec_block.block_w3_reg[6] ),
    .QN(_21702_));
 DFFR_X2 \core.dec_block.block_w3_reg[7]$_DFFE_PN0P_  (.D(_00692_),
    .RN(net90),
    .CK(clknet_leaf_311_clk),
    .Q(\core.dec_block.block_w3_reg[7] ),
    .QN(_21701_));
 DFFR_X2 \core.dec_block.block_w3_reg[8]$_DFFE_PN0P_  (.D(_00693_),
    .RN(net90),
    .CK(clknet_leaf_300_clk),
    .Q(\core.dec_block.block_w3_reg[8] ),
    .QN(_21700_));
 DFFR_X2 \core.dec_block.block_w3_reg[9]$_DFFE_PN0P_  (.D(_00694_),
    .RN(net91),
    .CK(clknet_leaf_302_clk),
    .Q(\core.dec_block.block_w3_reg[9] ),
    .QN(_21958_));
 DFFS_X2 \core.dec_block.dec_ctrl_reg[0]$_DFF_PN1_  (.D(_00009_),
    .SN(net94),
    .CK(clknet_leaf_252_clk),
    .Q(\core.dec_block.dec_ctrl_reg[0] ),
    .QN(_00325_));
 DFFR_X2 \core.dec_block.dec_ctrl_reg[1]$_DFF_PN0_  (.D(_00010_),
    .RN(net94),
    .CK(clknet_leaf_252_clk),
    .Q(\core.dec_block.dec_ctrl_reg[1] ),
    .QN(_00324_));
 DFFR_X1 \core.dec_block.dec_ctrl_reg[2]$_DFF_PN0_  (.D(_00000_),
    .RN(net94),
    .CK(clknet_leaf_252_clk),
    .Q(\core.dec_block.dec_ctrl_reg[2] ),
    .QN(_00174_));
 DFFR_X1 \core.dec_block.dec_ctrl_reg[3]$_DFF_PN0_  (.D(_00001_),
    .RN(net94),
    .CK(clknet_leaf_252_clk),
    .Q(\core.dec_block.dec_ctrl_reg[3] ),
    .QN(_21699_));
 DFFS_X2 \core.dec_block.ready_reg$_DFFE_PN1P_  (.D(_00695_),
    .SN(net94),
    .CK(clknet_leaf_259_clk),
    .Q(\core.dec_block.ready ),
    .QN(_21698_));
 DFFR_X1 \core.dec_block.round_ctr_reg[0]$_DFFE_PN0P_  (.D(_00696_),
    .RN(net96),
    .CK(clknet_leaf_261_clk),
    .Q(\core.dec_block.round[0] ),
    .QN(_22126_));
 DFFR_X1 \core.dec_block.round_ctr_reg[1]$_DFFE_PN0P_  (.D(_00697_),
    .RN(net96),
    .CK(clknet_leaf_251_clk),
    .Q(\core.dec_block.round[1] ),
    .QN(_22127_));
 DFFR_X1 \core.dec_block.round_ctr_reg[2]$_DFFE_PN0P_  (.D(_00698_),
    .RN(net94),
    .CK(clknet_leaf_259_clk),
    .Q(\core.dec_block.round[2] ),
    .QN(_21697_));
 DFFR_X1 \core.dec_block.round_ctr_reg[3]$_DFFE_PN0P_  (.D(_00699_),
    .RN(net96),
    .CK(clknet_leaf_251_clk),
    .Q(\core.dec_block.round[3] ),
    .QN(_21696_));
 DFFR_X2 \core.dec_block.sword_ctr_reg[0]$_DFFE_PN0P_  (.D(_00700_),
    .RN(net94),
    .CK(clknet_leaf_252_clk),
    .Q(\core.dec_block.sword_ctr_reg[0] ),
    .QN(_22130_));
 DFFR_X1 \core.dec_block.sword_ctr_reg[1]$_DFFE_PN0P_  (.D(_00701_),
    .RN(net94),
    .CK(clknet_leaf_252_clk),
    .Q(\core.dec_block.sword_ctr_reg[1] ),
    .QN(_22131_));
 DFFR_X2 \core.enc_block.block_w0_reg[0]$_DFFE_PN0P_  (.D(_00702_),
    .RN(net84),
    .CK(clknet_leaf_333_clk),
    .Q(\core.enc_block.block_w0_reg[0] ),
    .QN(_00360_));
 DFFR_X2 \core.enc_block.block_w0_reg[10]$_DFFE_PN0P_  (.D(_00703_),
    .RN(net84),
    .CK(clknet_leaf_342_clk),
    .Q(\core.enc_block.block_w0_reg[10] ),
    .QN(_00399_));
 DFFR_X2 \core.enc_block.block_w0_reg[11]$_DFFE_PN0P_  (.D(_00704_),
    .RN(net84),
    .CK(clknet_leaf_342_clk),
    .Q(\core.enc_block.block_w0_reg[11] ),
    .QN(_00402_));
 DFFR_X1 \core.enc_block.block_w0_reg[12]$_DFFE_PN0P_  (.D(_00705_),
    .RN(net84),
    .CK(clknet_leaf_342_clk),
    .Q(\core.enc_block.block_w0_reg[12] ),
    .QN(_00382_));
 DFFR_X2 \core.enc_block.block_w0_reg[13]$_DFFE_PN0P_  (.D(_00706_),
    .RN(net83),
    .CK(clknet_leaf_339_clk),
    .Q(\core.enc_block.block_w0_reg[13] ),
    .QN(_00385_));
 DFFR_X2 \core.enc_block.block_w0_reg[14]$_DFFE_PN0P_  (.D(_00707_),
    .RN(net83),
    .CK(clknet_leaf_341_clk),
    .Q(\core.enc_block.block_w0_reg[14] ),
    .QN(_00388_));
 DFFR_X1 \core.enc_block.block_w0_reg[15]$_DFFE_PN0P_  (.D(_00708_),
    .RN(net84),
    .CK(clknet_leaf_341_clk),
    .Q(\core.enc_block.block_w0_reg[15] ),
    .QN(_00391_));
 DFFR_X2 \core.enc_block.block_w0_reg[16]$_DFFE_PN0P_  (.D(_00709_),
    .RN(net84),
    .CK(clknet_leaf_332_clk),
    .Q(\core.enc_block.block_w0_reg[16] ),
    .QN(_00423_));
 DFFR_X1 \core.enc_block.block_w0_reg[17]$_DFFE_PN0P_  (.D(_00710_),
    .RN(net84),
    .CK(clknet_leaf_357_clk),
    .Q(\core.enc_block.block_w0_reg[17] ),
    .QN(_00426_));
 DFFR_X1 \core.enc_block.block_w0_reg[18]$_DFFE_PN0P_  (.D(_00711_),
    .RN(net83),
    .CK(clknet_leaf_339_clk),
    .Q(\core.enc_block.block_w0_reg[18] ),
    .QN(_00429_));
 DFFR_X2 \core.enc_block.block_w0_reg[19]$_DFFE_PN0P_  (.D(_00712_),
    .RN(net84),
    .CK(clknet_leaf_312_clk),
    .Q(\core.enc_block.block_w0_reg[19] ),
    .QN(_00432_));
 DFFR_X2 \core.enc_block.block_w0_reg[1]$_DFFE_PN0P_  (.D(_00713_),
    .RN(net84),
    .CK(clknet_leaf_332_clk),
    .Q(\core.enc_block.block_w0_reg[1] ),
    .QN(_00363_));
 DFFR_X2 \core.enc_block.block_w0_reg[20]$_DFFE_PN0P_  (.D(_00714_),
    .RN(net84),
    .CK(clknet_leaf_359_clk),
    .Q(\core.enc_block.block_w0_reg[20] ),
    .QN(_00412_));
 DFFR_X2 \core.enc_block.block_w0_reg[21]$_DFFE_PN0P_  (.D(_00715_),
    .RN(net84),
    .CK(clknet_leaf_312_clk),
    .Q(\core.enc_block.block_w0_reg[21] ),
    .QN(_00415_));
 DFFR_X2 \core.enc_block.block_w0_reg[22]$_DFFE_PN0P_  (.D(_00716_),
    .RN(net83),
    .CK(clknet_leaf_337_clk),
    .Q(\core.enc_block.block_w0_reg[22] ),
    .QN(_00418_));
 DFFR_X2 \core.enc_block.block_w0_reg[23]$_DFFE_PN0P_  (.D(_00717_),
    .RN(net83),
    .CK(clknet_leaf_333_clk),
    .Q(\core.enc_block.block_w0_reg[23] ),
    .QN(_00421_));
 DFFR_X1 \core.enc_block.block_w0_reg[24]$_DFFE_PN0P_  (.D(_00718_),
    .RN(net84),
    .CK(clknet_leaf_343_clk),
    .Q(\core.enc_block.block_w0_reg[24] ),
    .QN(_21695_));
 DFFR_X2 \core.enc_block.block_w0_reg[25]$_DFFE_PN0P_  (.D(_00719_),
    .RN(net83),
    .CK(clknet_leaf_358_clk),
    .Q(\core.enc_block.block_w0_reg[25] ),
    .QN(_00343_));
 DFFR_X1 \core.enc_block.block_w0_reg[26]$_DFFE_PN0P_  (.D(_00720_),
    .RN(net84),
    .CK(clknet_leaf_342_clk),
    .Q(\core.enc_block.block_w0_reg[26] ),
    .QN(_21694_));
 DFFR_X2 \core.enc_block.block_w0_reg[27]$_DFFE_PN0P_  (.D(_00721_),
    .RN(net84),
    .CK(clknet_leaf_342_clk),
    .Q(\core.enc_block.block_w0_reg[27] ),
    .QN(_00347_));
 DFFR_X2 \core.enc_block.block_w0_reg[28]$_DFFE_PN0P_  (.D(_00722_),
    .RN(net84),
    .CK(clknet_leaf_312_clk),
    .Q(\core.enc_block.block_w0_reg[28] ),
    .QN(_00330_));
 DFFR_X2 \core.enc_block.block_w0_reg[29]$_DFFE_PN0P_  (.D(_00723_),
    .RN(net83),
    .CK(clknet_leaf_338_clk),
    .Q(\core.enc_block.block_w0_reg[29] ),
    .QN(_00333_));
 DFFR_X2 \core.enc_block.block_w0_reg[2]$_DFFE_PN0P_  (.D(_00724_),
    .RN(net84),
    .CK(clknet_leaf_343_clk),
    .Q(\core.enc_block.block_w0_reg[2] ),
    .QN(_00366_));
 DFFR_X2 \core.enc_block.block_w0_reg[30]$_DFFE_PN0P_  (.D(_00725_),
    .RN(net84),
    .CK(clknet_leaf_333_clk),
    .Q(\core.enc_block.block_w0_reg[30] ),
    .QN(_00336_));
 DFFR_X2 \core.enc_block.block_w0_reg[31]$_DFFE_PN0P_  (.D(_00726_),
    .RN(net84),
    .CK(clknet_leaf_333_clk),
    .Q(\core.enc_block.block_w0_reg[31] ),
    .QN(_00339_));
 DFFR_X2 \core.enc_block.block_w0_reg[3]$_DFFE_PN0P_  (.D(_00727_),
    .RN(net83),
    .CK(clknet_leaf_334_clk),
    .Q(\core.enc_block.block_w0_reg[3] ),
    .QN(_00369_));
 DFFR_X2 \core.enc_block.block_w0_reg[4]$_DFFE_PN0P_  (.D(_00728_),
    .RN(net84),
    .CK(clknet_leaf_340_clk),
    .Q(\core.enc_block.block_w0_reg[4] ),
    .QN(_00349_));
 DFFR_X2 \core.enc_block.block_w0_reg[5]$_DFFE_PN0P_  (.D(_00729_),
    .RN(net83),
    .CK(clknet_leaf_338_clk),
    .Q(\core.enc_block.block_w0_reg[5] ),
    .QN(_00352_));
 DFFR_X2 \core.enc_block.block_w0_reg[6]$_DFFE_PN0P_  (.D(_00730_),
    .RN(net83),
    .CK(clknet_leaf_336_clk),
    .Q(\core.enc_block.block_w0_reg[6] ),
    .QN(_00355_));
 DFFR_X2 \core.enc_block.block_w0_reg[7]$_DFFE_PN0P_  (.D(_00731_),
    .RN(net84),
    .CK(clknet_leaf_342_clk),
    .Q(\core.enc_block.block_w0_reg[7] ),
    .QN(_00358_));
 DFFR_X2 \core.enc_block.block_w0_reg[8]$_DFFE_PN0P_  (.D(_00732_),
    .RN(net84),
    .CK(clknet_leaf_333_clk),
    .Q(\core.enc_block.block_w0_reg[8] ),
    .QN(_00393_));
 DFFR_X1 \core.enc_block.block_w0_reg[9]$_DFFE_PN0P_  (.D(_00733_),
    .RN(net84),
    .CK(clknet_leaf_332_clk),
    .Q(\core.enc_block.block_w0_reg[9] ),
    .QN(_00396_));
 DFFR_X1 \core.enc_block.block_w1_reg[0]$_DFFE_PN0P_  (.D(_00734_),
    .RN(net84),
    .CK(clknet_leaf_343_clk),
    .Q(\core.enc_block.block_w1_reg[0] ),
    .QN(_21693_));
 DFFR_X1 \core.enc_block.block_w1_reg[10]$_DFFE_PN0P_  (.D(_00735_),
    .RN(net84),
    .CK(clknet_leaf_342_clk),
    .Q(\core.enc_block.block_w1_reg[10] ),
    .QN(_21692_));
 DFFR_X1 \core.enc_block.block_w1_reg[11]$_DFFE_PN0P_  (.D(_00736_),
    .RN(net83),
    .CK(clknet_leaf_337_clk),
    .Q(\core.enc_block.block_w1_reg[11] ),
    .QN(_00303_));
 DFFR_X2 \core.enc_block.block_w1_reg[12]$_DFFE_PN0P_  (.D(_00737_),
    .RN(net83),
    .CK(clknet_leaf_337_clk),
    .Q(\core.enc_block.block_w1_reg[12] ),
    .QN(_00304_));
 DFFR_X1 \core.enc_block.block_w1_reg[13]$_DFFE_PN0P_  (.D(_00738_),
    .RN(net83),
    .CK(clknet_leaf_359_clk),
    .Q(\core.enc_block.block_w1_reg[13] ),
    .QN(_00306_));
 DFFR_X1 \core.enc_block.block_w1_reg[14]$_DFFE_PN0P_  (.D(_00739_),
    .RN(net83),
    .CK(clknet_leaf_338_clk),
    .Q(\core.enc_block.block_w1_reg[14] ),
    .QN(_00307_));
 DFFR_X1 \core.enc_block.block_w1_reg[15]$_DFFE_PN0P_  (.D(_00740_),
    .RN(net83),
    .CK(clknet_leaf_339_clk),
    .Q(\core.enc_block.block_w1_reg[15] ),
    .QN(_21691_));
 DFFR_X1 \core.enc_block.block_w1_reg[16]$_DFFE_PN0P_  (.D(_00741_),
    .RN(net83),
    .CK(clknet_leaf_330_clk),
    .Q(\core.enc_block.block_w1_reg[16] ),
    .QN(_21690_));
 DFFR_X1 \core.enc_block.block_w1_reg[17]$_DFFE_PN0P_  (.D(_00742_),
    .RN(net84),
    .CK(clknet_leaf_356_clk),
    .Q(\core.enc_block.block_w1_reg[17] ),
    .QN(_21689_));
 DFFR_X1 \core.enc_block.block_w1_reg[18]$_DFFE_PN0P_  (.D(_00743_),
    .RN(net84),
    .CK(clknet_leaf_331_clk),
    .Q(\core.enc_block.block_w1_reg[18] ),
    .QN(_21688_));
 DFFR_X1 \core.enc_block.block_w1_reg[19]$_DFFE_PN0P_  (.D(_00744_),
    .RN(net83),
    .CK(clknet_leaf_358_clk),
    .Q(\core.enc_block.block_w1_reg[19] ),
    .QN(_21687_));
 DFFR_X1 \core.enc_block.block_w1_reg[1]$_DFFE_PN0P_  (.D(_00745_),
    .RN(net84),
    .CK(clknet_leaf_341_clk),
    .Q(\core.enc_block.block_w1_reg[1] ),
    .QN(_21686_));
 DFFR_X1 \core.enc_block.block_w1_reg[20]$_DFFE_PN0P_  (.D(_00746_),
    .RN(net84),
    .CK(clknet_leaf_355_clk),
    .Q(\core.enc_block.block_w1_reg[20] ),
    .QN(_21685_));
 DFFR_X1 \core.enc_block.block_w1_reg[21]$_DFFE_PN0P_  (.D(_00747_),
    .RN(net83),
    .CK(clknet_leaf_335_clk),
    .Q(\core.enc_block.block_w1_reg[21] ),
    .QN(_21684_));
 DFFR_X1 \core.enc_block.block_w1_reg[22]$_DFFE_PN0P_  (.D(_00748_),
    .RN(net83),
    .CK(clknet_leaf_335_clk),
    .Q(\core.enc_block.block_w1_reg[22] ),
    .QN(_21683_));
 DFFR_X1 \core.enc_block.block_w1_reg[23]$_DFFE_PN0P_  (.D(_00749_),
    .RN(net84),
    .CK(clknet_leaf_331_clk),
    .Q(\core.enc_block.block_w1_reg[23] ),
    .QN(_21682_));
 DFFR_X1 \core.enc_block.block_w1_reg[24]$_DFFE_PN0P_  (.D(_00750_),
    .RN(net84),
    .CK(clknet_leaf_343_clk),
    .Q(\core.enc_block.block_w1_reg[24] ),
    .QN(_21681_));
 DFFR_X1 \core.enc_block.block_w1_reg[25]$_DFFE_PN0P_  (.D(_00751_),
    .RN(net84),
    .CK(clknet_leaf_343_clk),
    .Q(\core.enc_block.block_w1_reg[25] ),
    .QN(_21680_));
 DFFR_X1 \core.enc_block.block_w1_reg[26]$_DFFE_PN0P_  (.D(_00752_),
    .RN(net83),
    .CK(clknet_leaf_330_clk),
    .Q(\core.enc_block.block_w1_reg[26] ),
    .QN(_21679_));
 DFFR_X1 \core.enc_block.block_w1_reg[27]$_DFFE_PN0P_  (.D(_00753_),
    .RN(net83),
    .CK(clknet_leaf_329_clk),
    .Q(\core.enc_block.block_w1_reg[27] ),
    .QN(_21678_));
 DFFR_X1 \core.enc_block.block_w1_reg[28]$_DFFE_PN0P_  (.D(_00754_),
    .RN(net83),
    .CK(clknet_leaf_334_clk),
    .Q(\core.enc_block.block_w1_reg[28] ),
    .QN(_00311_));
 DFFR_X1 \core.enc_block.block_w1_reg[29]$_DFFE_PN0P_  (.D(_00755_),
    .RN(net84),
    .CK(clknet_leaf_339_clk),
    .Q(\core.enc_block.block_w1_reg[29] ),
    .QN(_21677_));
 DFFR_X1 \core.enc_block.block_w1_reg[2]$_DFFE_PN0P_  (.D(_00756_),
    .RN(net84),
    .CK(clknet_leaf_344_clk),
    .Q(\core.enc_block.block_w1_reg[2] ),
    .QN(_21676_));
 DFFR_X1 \core.enc_block.block_w1_reg[30]$_DFFE_PN0P_  (.D(_00757_),
    .RN(net83),
    .CK(clknet_leaf_336_clk),
    .Q(\core.enc_block.block_w1_reg[30] ),
    .QN(_21675_));
 DFFR_X1 \core.enc_block.block_w1_reg[31]$_DFFE_PN0P_  (.D(_00758_),
    .RN(net84),
    .CK(clknet_leaf_332_clk),
    .Q(\core.enc_block.block_w1_reg[31] ),
    .QN(_21674_));
 DFFR_X1 \core.enc_block.block_w1_reg[3]$_DFFE_PN0P_  (.D(_00759_),
    .RN(net84),
    .CK(clknet_leaf_340_clk),
    .Q(\core.enc_block.block_w1_reg[3] ),
    .QN(_21673_));
 DFFR_X1 \core.enc_block.block_w1_reg[4]$_DFFE_PN0P_  (.D(_00760_),
    .RN(net84),
    .CK(clknet_leaf_340_clk),
    .Q(\core.enc_block.block_w1_reg[4] ),
    .QN(_21672_));
 DFFR_X1 \core.enc_block.block_w1_reg[5]$_DFFE_PN0P_  (.D(_00761_),
    .RN(net84),
    .CK(clknet_leaf_340_clk),
    .Q(\core.enc_block.block_w1_reg[5] ),
    .QN(_21671_));
 DFFR_X1 \core.enc_block.block_w1_reg[6]$_DFFE_PN0P_  (.D(_00762_),
    .RN(net84),
    .CK(clknet_leaf_340_clk),
    .Q(\core.enc_block.block_w1_reg[6] ),
    .QN(_21670_));
 DFFR_X2 \core.enc_block.block_w1_reg[7]$_DFFE_PN0P_  (.D(_00763_),
    .RN(net83),
    .CK(clknet_leaf_341_clk),
    .Q(\core.enc_block.block_w1_reg[7] ),
    .QN(_00308_));
 DFFR_X1 \core.enc_block.block_w1_reg[8]$_DFFE_PN0P_  (.D(_00764_),
    .RN(net84),
    .CK(clknet_leaf_331_clk),
    .Q(\core.enc_block.block_w1_reg[8] ),
    .QN(_21669_));
 DFFR_X1 \core.enc_block.block_w1_reg[9]$_DFFE_PN0P_  (.D(_00765_),
    .RN(net83),
    .CK(clknet_leaf_336_clk),
    .Q(\core.enc_block.block_w1_reg[9] ),
    .QN(_00305_));
 DFFR_X1 \core.enc_block.block_w2_reg[0]$_DFFE_PN0P_  (.D(_00766_),
    .RN(net84),
    .CK(clknet_leaf_341_clk),
    .Q(\core.enc_block.block_w2_reg[0] ),
    .QN(_21668_));
 DFFR_X1 \core.enc_block.block_w2_reg[10]$_DFFE_PN0P_  (.D(_00767_),
    .RN(net84),
    .CK(clknet_leaf_331_clk),
    .Q(\core.enc_block.block_w2_reg[10] ),
    .QN(_21667_));
 DFFR_X1 \core.enc_block.block_w2_reg[11]$_DFFE_PN0P_  (.D(_00768_),
    .RN(net83),
    .CK(clknet_leaf_337_clk),
    .Q(\core.enc_block.block_w2_reg[11] ),
    .QN(_00313_));
 DFFR_X1 \core.enc_block.block_w2_reg[12]$_DFFE_PN0P_  (.D(_00769_),
    .RN(net83),
    .CK(clknet_leaf_337_clk),
    .Q(\core.enc_block.block_w2_reg[12] ),
    .QN(_00314_));
 DFFR_X1 \core.enc_block.block_w2_reg[13]$_DFFE_PN0P_  (.D(_00770_),
    .RN(net84),
    .CK(clknet_leaf_293_clk),
    .Q(\core.enc_block.block_w2_reg[13] ),
    .QN(_00316_));
 DFFR_X1 \core.enc_block.block_w2_reg[14]$_DFFE_PN0P_  (.D(_00771_),
    .RN(net84),
    .CK(clknet_leaf_360_clk),
    .Q(\core.enc_block.block_w2_reg[14] ),
    .QN(_00317_));
 DFFR_X1 \core.enc_block.block_w2_reg[15]$_DFFE_PN0P_  (.D(_00772_),
    .RN(net84),
    .CK(clknet_leaf_360_clk),
    .Q(\core.enc_block.block_w2_reg[15] ),
    .QN(_00315_));
 DFFR_X1 \core.enc_block.block_w2_reg[16]$_DFFE_PN0P_  (.D(_00773_),
    .RN(net84),
    .CK(clknet_leaf_331_clk),
    .Q(\core.enc_block.block_w2_reg[16] ),
    .QN(_21666_));
 DFFR_X1 \core.enc_block.block_w2_reg[17]$_DFFE_PN0P_  (.D(_00774_),
    .RN(net84),
    .CK(clknet_leaf_357_clk),
    .Q(\core.enc_block.block_w2_reg[17] ),
    .QN(_21665_));
 DFFR_X1 \core.enc_block.block_w2_reg[18]$_DFFE_PN0P_  (.D(_00775_),
    .RN(net84),
    .CK(clknet_leaf_356_clk),
    .Q(\core.enc_block.block_w2_reg[18] ),
    .QN(_21664_));
 DFFR_X1 \core.enc_block.block_w2_reg[19]$_DFFE_PN0P_  (.D(_00776_),
    .RN(net84),
    .CK(clknet_leaf_354_clk),
    .Q(\core.enc_block.block_w2_reg[19] ),
    .QN(_21663_));
 DFFR_X1 \core.enc_block.block_w2_reg[1]$_DFFE_PN0P_  (.D(_00777_),
    .RN(net84),
    .CK(clknet_leaf_355_clk),
    .Q(\core.enc_block.block_w2_reg[1] ),
    .QN(_21662_));
 DFFR_X1 \core.enc_block.block_w2_reg[20]$_DFFE_PN0P_  (.D(_00778_),
    .RN(net84),
    .CK(clknet_leaf_359_clk),
    .Q(\core.enc_block.block_w2_reg[20] ),
    .QN(_21661_));
 DFFR_X1 \core.enc_block.block_w2_reg[21]$_DFFE_PN0P_  (.D(_00779_),
    .RN(net84),
    .CK(clknet_leaf_354_clk),
    .Q(\core.enc_block.block_w2_reg[21] ),
    .QN(_21660_));
 DFFR_X1 \core.enc_block.block_w2_reg[22]$_DFFE_PN0P_  (.D(_00780_),
    .RN(net83),
    .CK(clknet_leaf_335_clk),
    .Q(\core.enc_block.block_w2_reg[22] ),
    .QN(_21659_));
 DFFR_X1 \core.enc_block.block_w2_reg[23]$_DFFE_PN0P_  (.D(_00781_),
    .RN(net83),
    .CK(clknet_leaf_338_clk),
    .Q(\core.enc_block.block_w2_reg[23] ),
    .QN(_21658_));
 DFFR_X1 \core.enc_block.block_w2_reg[24]$_DFFE_PN0P_  (.D(_00782_),
    .RN(net84),
    .CK(clknet_leaf_341_clk),
    .Q(\core.enc_block.block_w2_reg[24] ),
    .QN(_21657_));
 DFFR_X1 \core.enc_block.block_w2_reg[25]$_DFFE_PN0P_  (.D(_00783_),
    .RN(net84),
    .CK(clknet_leaf_344_clk),
    .Q(\core.enc_block.block_w2_reg[25] ),
    .QN(_00309_));
 DFFR_X1 \core.enc_block.block_w2_reg[26]$_DFFE_PN0P_  (.D(_00784_),
    .RN(net83),
    .CK(clknet_leaf_330_clk),
    .Q(\core.enc_block.block_w2_reg[26] ),
    .QN(_21656_));
 DFFR_X1 \core.enc_block.block_w2_reg[27]$_DFFE_PN0P_  (.D(_00785_),
    .RN(net84),
    .CK(clknet_leaf_331_clk),
    .Q(\core.enc_block.block_w2_reg[27] ),
    .QN(_21655_));
 DFFR_X2 \core.enc_block.block_w2_reg[28]$_DFFE_PN0P_  (.D(_00786_),
    .RN(net83),
    .CK(clknet_leaf_335_clk),
    .Q(\core.enc_block.block_w2_reg[28] ),
    .QN(_00310_));
 DFFR_X1 \core.enc_block.block_w2_reg[29]$_DFFE_PN0P_  (.D(_00787_),
    .RN(net83),
    .CK(clknet_leaf_335_clk),
    .Q(\core.enc_block.block_w2_reg[29] ),
    .QN(_21654_));
 DFFR_X1 \core.enc_block.block_w2_reg[2]$_DFFE_PN0P_  (.D(_00788_),
    .RN(net84),
    .CK(clknet_leaf_355_clk),
    .Q(\core.enc_block.block_w2_reg[2] ),
    .QN(_21653_));
 DFFR_X1 \core.enc_block.block_w2_reg[30]$_DFFE_PN0P_  (.D(_00789_),
    .RN(net83),
    .CK(clknet_leaf_330_clk),
    .Q(\core.enc_block.block_w2_reg[30] ),
    .QN(_21652_));
 DFFR_X1 \core.enc_block.block_w2_reg[31]$_DFFE_PN0P_  (.D(_00790_),
    .RN(net83),
    .CK(clknet_leaf_331_clk),
    .Q(\core.enc_block.block_w2_reg[31] ),
    .QN(_21651_));
 DFFR_X1 \core.enc_block.block_w2_reg[3]$_DFFE_PN0P_  (.D(_00791_),
    .RN(net83),
    .CK(clknet_leaf_336_clk),
    .Q(\core.enc_block.block_w2_reg[3] ),
    .QN(_21650_));
 DFFR_X1 \core.enc_block.block_w2_reg[4]$_DFFE_PN0P_  (.D(_00792_),
    .RN(net84),
    .CK(clknet_leaf_354_clk),
    .Q(\core.enc_block.block_w2_reg[4] ),
    .QN(_21649_));
 DFFR_X1 \core.enc_block.block_w2_reg[5]$_DFFE_PN0P_  (.D(_00793_),
    .RN(net84),
    .CK(clknet_leaf_355_clk),
    .Q(\core.enc_block.block_w2_reg[5] ),
    .QN(_21648_));
 DFFR_X1 \core.enc_block.block_w2_reg[6]$_DFFE_PN0P_  (.D(_00794_),
    .RN(net83),
    .CK(clknet_leaf_335_clk),
    .Q(\core.enc_block.block_w2_reg[6] ),
    .QN(_21647_));
 DFFR_X1 \core.enc_block.block_w2_reg[7]$_DFFE_PN0P_  (.D(_00795_),
    .RN(net83),
    .CK(clknet_leaf_358_clk),
    .Q(\core.enc_block.block_w2_reg[7] ),
    .QN(_00302_));
 DFFR_X1 \core.enc_block.block_w2_reg[8]$_DFFE_PN0P_  (.D(_00796_),
    .RN(net83),
    .CK(clknet_leaf_338_clk),
    .Q(\core.enc_block.block_w2_reg[8] ),
    .QN(_21646_));
 DFFR_X2 \core.enc_block.block_w2_reg[9]$_DFFE_PN0P_  (.D(_00797_),
    .RN(net84),
    .CK(clknet_leaf_313_clk),
    .Q(\core.enc_block.block_w2_reg[9] ),
    .QN(_00312_));
 DFFR_X2 \core.enc_block.block_w3_reg[0]$_DFFE_PN0P_  (.D(_00798_),
    .RN(net83),
    .CK(clknet_leaf_338_clk),
    .Q(\core.enc_block.block_w3_reg[0] ),
    .QN(_00361_));
 DFFR_X2 \core.enc_block.block_w3_reg[10]$_DFFE_PN0P_  (.D(_00799_),
    .RN(net83),
    .CK(clknet_leaf_332_clk),
    .Q(\core.enc_block.block_w3_reg[10] ),
    .QN(_00400_));
 DFFR_X2 \core.enc_block.block_w3_reg[11]$_DFFE_PN0P_  (.D(_00800_),
    .RN(net83),
    .CK(clknet_leaf_334_clk),
    .Q(\core.enc_block.block_w3_reg[11] ),
    .QN(_00403_));
 DFFR_X1 \core.enc_block.block_w3_reg[12]$_DFFE_PN0P_  (.D(_00801_),
    .RN(net83),
    .CK(clknet_leaf_334_clk),
    .Q(\core.enc_block.block_w3_reg[12] ),
    .QN(_00383_));
 DFFR_X1 \core.enc_block.block_w3_reg[13]$_DFFE_PN0P_  (.D(_00802_),
    .RN(net84),
    .CK(clknet_leaf_357_clk),
    .Q(\core.enc_block.block_w3_reg[13] ),
    .QN(_00386_));
 DFFR_X1 \core.enc_block.block_w3_reg[14]$_DFFE_PN0P_  (.D(_00803_),
    .RN(net83),
    .CK(clknet_leaf_339_clk),
    .Q(\core.enc_block.block_w3_reg[14] ),
    .QN(_00389_));
 DFFR_X2 \core.enc_block.block_w3_reg[15]$_DFFE_PN0P_  (.D(_00804_),
    .RN(net84),
    .CK(clknet_leaf_343_clk),
    .Q(\core.enc_block.block_w3_reg[15] ),
    .QN(_00392_));
 DFFR_X1 \core.enc_block.block_w3_reg[16]$_DFFE_PN0P_  (.D(_00805_),
    .RN(net83),
    .CK(clknet_leaf_334_clk),
    .Q(\core.enc_block.block_w3_reg[16] ),
    .QN(_00424_));
 DFFR_X1 \core.enc_block.block_w3_reg[17]$_DFFE_PN0P_  (.D(_00806_),
    .RN(net84),
    .CK(clknet_leaf_344_clk),
    .Q(\core.enc_block.block_w3_reg[17] ),
    .QN(_00427_));
 DFFR_X1 \core.enc_block.block_w3_reg[18]$_DFFE_PN0P_  (.D(_00807_),
    .RN(net84),
    .CK(clknet_leaf_343_clk),
    .Q(\core.enc_block.block_w3_reg[18] ),
    .QN(_00430_));
 DFFR_X2 \core.enc_block.block_w3_reg[19]$_DFFE_PN0P_  (.D(_00808_),
    .RN(net84),
    .CK(clknet_leaf_344_clk),
    .Q(\core.enc_block.block_w3_reg[19] ),
    .QN(_00433_));
 DFFR_X2 \core.enc_block.block_w3_reg[1]$_DFFE_PN0P_  (.D(_00809_),
    .RN(net84),
    .CK(clknet_leaf_359_clk),
    .Q(\core.enc_block.block_w3_reg[1] ),
    .QN(_00364_));
 DFFR_X2 \core.enc_block.block_w3_reg[20]$_DFFE_PN0P_  (.D(_00810_),
    .RN(net84),
    .CK(clknet_leaf_340_clk),
    .Q(\core.enc_block.block_w3_reg[20] ),
    .QN(_00413_));
 DFFR_X1 \core.enc_block.block_w3_reg[21]$_DFFE_PN0P_  (.D(_00811_),
    .RN(net84),
    .CK(clknet_leaf_357_clk),
    .Q(\core.enc_block.block_w3_reg[21] ),
    .QN(_00416_));
 DFFR_X2 \core.enc_block.block_w3_reg[22]$_DFFE_PN0P_  (.D(_00812_),
    .RN(net83),
    .CK(clknet_leaf_334_clk),
    .Q(\core.enc_block.block_w3_reg[22] ),
    .QN(_00419_));
 DFFR_X1 \core.enc_block.block_w3_reg[23]$_DFFE_PN0P_  (.D(_00813_),
    .RN(net84),
    .CK(clknet_leaf_344_clk),
    .Q(\core.enc_block.block_w3_reg[23] ),
    .QN(_00422_));
 DFFR_X1 \core.enc_block.block_w3_reg[24]$_DFFE_PN0P_  (.D(_00814_),
    .RN(net83),
    .CK(clknet_leaf_339_clk),
    .Q(\core.enc_block.block_w3_reg[24] ),
    .QN(_00341_));
 DFFR_X1 \core.enc_block.block_w3_reg[25]$_DFFE_PN0P_  (.D(_00815_),
    .RN(net83),
    .CK(clknet_leaf_357_clk),
    .Q(\core.enc_block.block_w3_reg[25] ),
    .QN(_00344_));
 DFFR_X2 \core.enc_block.block_w3_reg[26]$_DFFE_PN0P_  (.D(_00816_),
    .RN(net83),
    .CK(clknet_leaf_314_clk),
    .Q(\core.enc_block.block_w3_reg[26] ),
    .QN(_21645_));
 DFFR_X2 \core.enc_block.block_w3_reg[27]$_DFFE_PN0P_  (.D(_00817_),
    .RN(net83),
    .CK(clknet_leaf_336_clk),
    .Q(\core.enc_block.block_w3_reg[27] ),
    .QN(_00348_));
 DFFR_X2 \core.enc_block.block_w3_reg[28]$_DFFE_PN0P_  (.D(_00818_),
    .RN(net84),
    .CK(clknet_leaf_313_clk),
    .Q(\core.enc_block.block_w3_reg[28] ),
    .QN(_00331_));
 DFFR_X1 \core.enc_block.block_w3_reg[29]$_DFFE_PN0P_  (.D(_00819_),
    .RN(net83),
    .CK(clknet_leaf_359_clk),
    .Q(\core.enc_block.block_w3_reg[29] ),
    .QN(_00334_));
 DFFR_X2 \core.enc_block.block_w3_reg[2]$_DFFE_PN0P_  (.D(_00820_),
    .RN(net83),
    .CK(clknet_leaf_358_clk),
    .Q(\core.enc_block.block_w3_reg[2] ),
    .QN(_00367_));
 DFFR_X1 \core.enc_block.block_w3_reg[30]$_DFFE_PN0P_  (.D(_00821_),
    .RN(net83),
    .CK(clknet_leaf_337_clk),
    .Q(\core.enc_block.block_w3_reg[30] ),
    .QN(_00337_));
 DFFR_X2 \core.enc_block.block_w3_reg[31]$_DFFE_PN0P_  (.D(_00822_),
    .RN(net83),
    .CK(clknet_leaf_337_clk),
    .Q(\core.enc_block.block_w3_reg[31] ),
    .QN(_00340_));
 DFFR_X2 \core.enc_block.block_w3_reg[3]$_DFFE_PN0P_  (.D(_00823_),
    .RN(net83),
    .CK(clknet_leaf_358_clk),
    .Q(\core.enc_block.block_w3_reg[3] ),
    .QN(_00370_));
 DFFR_X2 \core.enc_block.block_w3_reg[4]$_DFFE_PN0P_  (.D(_00824_),
    .RN(net84),
    .CK(clknet_leaf_358_clk),
    .Q(\core.enc_block.block_w3_reg[4] ),
    .QN(_00350_));
 DFFR_X2 \core.enc_block.block_w3_reg[5]$_DFFE_PN0P_  (.D(_00825_),
    .RN(net84),
    .CK(clknet_leaf_360_clk),
    .Q(\core.enc_block.block_w3_reg[5] ),
    .QN(_00353_));
 DFFR_X2 \core.enc_block.block_w3_reg[6]$_DFFE_PN0P_  (.D(_00826_),
    .RN(net84),
    .CK(clknet_leaf_312_clk),
    .Q(\core.enc_block.block_w3_reg[6] ),
    .QN(_00356_));
 DFFR_X1 \core.enc_block.block_w3_reg[7]$_DFFE_PN0P_  (.D(_00827_),
    .RN(net84),
    .CK(clknet_leaf_360_clk),
    .Q(\core.enc_block.block_w3_reg[7] ),
    .QN(_00359_));
 DFFR_X2 \core.enc_block.block_w3_reg[8]$_DFFE_PN0P_  (.D(_00828_),
    .RN(net83),
    .CK(clknet_leaf_332_clk),
    .Q(\core.enc_block.block_w3_reg[8] ),
    .QN(_00394_));
 DFFR_X1 \core.enc_block.block_w3_reg[9]$_DFFE_PN0P_  (.D(_00829_),
    .RN(net83),
    .CK(clknet_leaf_332_clk),
    .Q(\core.enc_block.block_w3_reg[9] ),
    .QN(_00397_));
 DFFS_X1 \core.enc_block.enc_ctrl_reg[0]$_DFF_PN1_  (.D(_00011_),
    .SN(net84),
    .CK(clknet_leaf_349_clk),
    .Q(\core.enc_block.enc_ctrl_reg[0] ),
    .QN(_00322_));
 DFFR_X1 \core.enc_block.enc_ctrl_reg[1]$_DFF_PN0_  (.D(_00012_),
    .RN(net84),
    .CK(clknet_leaf_349_clk),
    .Q(\core.enc_block.enc_ctrl_reg[1] ),
    .QN(_00321_));
 DFFR_X1 \core.enc_block.enc_ctrl_reg[2]$_DFF_PN0_  (.D(_00002_),
    .RN(net84),
    .CK(clknet_leaf_349_clk),
    .Q(\core.enc_block.enc_ctrl_reg[2] ),
    .QN(_00329_));
 DFFR_X1 \core.enc_block.enc_ctrl_reg[3]$_DFF_PN0_  (.D(_00003_),
    .RN(net84),
    .CK(clknet_leaf_344_clk),
    .Q(\core.enc_block.enc_ctrl_reg[3] ),
    .QN(_21644_));
 DFFS_X1 \core.enc_block.ready_reg$_DFFE_PN1P_  (.D(_00830_),
    .SN(net84),
    .CK(clknet_leaf_356_clk),
    .Q(\core.enc_block.ready ),
    .QN(_21643_));
 DFFR_X2 \core.enc_block.round_ctr_reg[0]$_DFFE_PN0P_  (.D(_00831_),
    .RN(net94),
    .CK(clknet_leaf_213_clk),
    .Q(\core.enc_block.round[0] ),
    .QN(_21642_));
 DFFR_X1 \core.enc_block.round_ctr_reg[1]$_DFFE_PN0P_  (.D(_00832_),
    .RN(net91),
    .CK(clknet_leaf_284_clk),
    .Q(\core.enc_block.round[1] ),
    .QN(_21641_));
 DFFR_X2 \core.enc_block.round_ctr_reg[2]$_DFFE_PN0P_  (.D(_00833_),
    .RN(net91),
    .CK(clknet_leaf_284_clk),
    .Q(\core.enc_block.round[2] ),
    .QN(_21640_));
 DFFR_X2 \core.enc_block.round_ctr_reg[3]$_DFFE_PN0P_  (.D(_00834_),
    .RN(net94),
    .CK(clknet_leaf_213_clk),
    .Q(\core.enc_block.round[3] ),
    .QN(_00323_));
 DFFR_X2 \core.enc_block.sword_ctr_reg[0]$_DFFE_PN0P_  (.D(_00835_),
    .RN(net86),
    .CK(clknet_leaf_345_clk),
    .Q(\core.enc_block.sword_ctr_reg[0] ),
    .QN(_22116_));
 DFFR_X1 \core.enc_block.sword_ctr_reg[1]$_DFFE_PN0P_  (.D(_00836_),
    .RN(net86),
    .CK(clknet_leaf_344_clk),
    .Q(\core.enc_block.sword_ctr_reg[1] ),
    .QN(_22117_));
 DFFR_X1 \core.keymem.key_mem[0][0]$_DFFE_PN0P_  (.D(_00837_),
    .RN(net94),
    .CK(clknet_leaf_220_clk),
    .Q(\core.keymem.key_mem[0][0] ),
    .QN(_00173_));
 DFFR_X1 \core.keymem.key_mem[0][100]$_DFFE_PN0P_  (.D(_00838_),
    .RN(net94),
    .CK(clknet_leaf_208_clk),
    .Q(\core.keymem.key_mem[0][100] ),
    .QN(_00210_));
 DFFR_X2 \core.keymem.key_mem[0][101]$_DFFE_PN0P_  (.D(_00839_),
    .RN(net93),
    .CK(clknet_leaf_374_clk),
    .Q(\core.keymem.key_mem[0][101] ),
    .QN(_00183_));
 DFFR_X1 \core.keymem.key_mem[0][102]$_DFFE_PN0P_  (.D(_00840_),
    .RN(net94),
    .CK(clknet_leaf_212_clk),
    .Q(\core.keymem.key_mem[0][102] ),
    .QN(_00184_));
 DFFR_X1 \core.keymem.key_mem[0][103]$_DFFE_PN0P_  (.D(_00841_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[0][103] ),
    .QN(_00185_));
 DFFR_X1 \core.keymem.key_mem[0][104]$_DFFE_PN0P_  (.D(_00842_),
    .RN(net92),
    .CK(clknet_leaf_201_clk),
    .Q(\core.keymem.key_mem[0][104] ),
    .QN(_00182_));
 DFFR_X1 \core.keymem.key_mem[0][105]$_DFFE_PN0P_  (.D(_00843_),
    .RN(net92),
    .CK(clknet_leaf_267_clk),
    .Q(\core.keymem.key_mem[0][105] ),
    .QN(_00193_));
 DFFR_X1 \core.keymem.key_mem[0][106]$_DFFE_PN0P_  (.D(_00844_),
    .RN(net92),
    .CK(clknet_leaf_277_clk),
    .Q(\core.keymem.key_mem[0][106] ),
    .QN(_00199_));
 DFFR_X1 \core.keymem.key_mem[0][107]$_DFFE_PN0P_  (.D(_00845_),
    .RN(net92),
    .CK(clknet_leaf_272_clk),
    .Q(\core.keymem.key_mem[0][107] ),
    .QN(_00204_));
 DFFR_X1 \core.keymem.key_mem[0][108]$_DFFE_PN0P_  (.D(_00846_),
    .RN(net91),
    .CK(clknet_leaf_278_clk),
    .Q(\core.keymem.key_mem[0][108] ),
    .QN(_00209_));
 DFFR_X1 \core.keymem.key_mem[0][109]$_DFFE_PN0P_  (.D(_00847_),
    .RN(net92),
    .CK(clknet_leaf_268_clk),
    .Q(\core.keymem.key_mem[0][109] ),
    .QN(_00181_));
 DFFR_X1 \core.keymem.key_mem[0][10]$_DFFE_PN0P_  (.D(_00848_),
    .RN(net89),
    .CK(clknet_leaf_381_clk),
    .Q(\core.keymem.key_mem[0][10] ),
    .QN(_00235_));
 DFFR_X2 \core.keymem.key_mem[0][110]$_DFFE_PN0P_  (.D(_00849_),
    .RN(net96),
    .CK(clknet_leaf_213_clk),
    .Q(\core.keymem.key_mem[0][110] ),
    .QN(_00192_));
 DFFR_X1 \core.keymem.key_mem[0][111]$_DFFE_PN0P_  (.D(_00850_),
    .RN(net94),
    .CK(clknet_leaf_215_clk),
    .Q(\core.keymem.key_mem[0][111] ),
    .QN(_00198_));
 DFFR_X1 \core.keymem.key_mem[0][112]$_DFFE_PN0P_  (.D(_00851_),
    .RN(net94),
    .CK(clknet_leaf_263_clk),
    .Q(\core.keymem.key_mem[0][112] ),
    .QN(_00180_));
 DFFR_X1 \core.keymem.key_mem[0][113]$_DFFE_PN0P_  (.D(_00852_),
    .RN(net91),
    .CK(clknet_leaf_273_clk),
    .Q(\core.keymem.key_mem[0][113] ),
    .QN(_00191_));
 DFFR_X1 \core.keymem.key_mem[0][114]$_DFFE_PN0P_  (.D(_00853_),
    .RN(net91),
    .CK(clknet_leaf_284_clk),
    .Q(\core.keymem.key_mem[0][114] ),
    .QN(_00197_));
 DFFR_X1 \core.keymem.key_mem[0][115]$_DFFE_PN0P_  (.D(_00854_),
    .RN(net91),
    .CK(clknet_leaf_288_clk),
    .Q(\core.keymem.key_mem[0][115] ),
    .QN(_00203_));
 DFFR_X1 \core.keymem.key_mem[0][116]$_DFFE_PN0P_  (.D(_00855_),
    .RN(net92),
    .CK(clknet_leaf_267_clk),
    .Q(\core.keymem.key_mem[0][116] ),
    .QN(_00208_));
 DFFR_X1 \core.keymem.key_mem[0][117]$_DFFE_PN0P_  (.D(_00856_),
    .RN(net91),
    .CK(clknet_leaf_288_clk),
    .Q(\core.keymem.key_mem[0][117] ),
    .QN(_00178_));
 DFFR_X1 \core.keymem.key_mem[0][118]$_DFFE_PN0P_  (.D(_00857_),
    .RN(net93),
    .CK(clknet_leaf_373_clk),
    .Q(\core.keymem.key_mem[0][118] ),
    .QN(_00179_));
 DFFR_X1 \core.keymem.key_mem[0][119]$_DFFE_PN0P_  (.D(_00858_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[0][119] ),
    .QN(_00190_));
 DFFR_X1 \core.keymem.key_mem[0][11]$_DFFE_PN0P_  (.D(_00859_),
    .RN(net89),
    .CK(clknet_leaf_53_clk),
    .Q(\core.keymem.key_mem[0][11] ),
    .QN(_00241_));
 DFFR_X1 \core.keymem.key_mem[0][120]$_DFFE_PN0P_  (.D(_00860_),
    .RN(net94),
    .CK(clknet_leaf_204_clk),
    .Q(\core.keymem.key_mem[0][120] ),
    .QN(_00177_));
 DFFR_X1 \core.keymem.key_mem[0][121]$_DFFE_PN0P_  (.D(_00861_),
    .RN(net92),
    .CK(clknet_leaf_268_clk),
    .Q(\core.keymem.key_mem[0][121] ),
    .QN(_00189_));
 DFFR_X1 \core.keymem.key_mem[0][122]$_DFFE_PN0P_  (.D(_00862_),
    .RN(net89),
    .CK(clknet_leaf_375_clk),
    .Q(\core.keymem.key_mem[0][122] ),
    .QN(_00196_));
 DFFR_X1 \core.keymem.key_mem[0][123]$_DFFE_PN0P_  (.D(_00863_),
    .RN(net93),
    .CK(clknet_leaf_197_clk),
    .Q(\core.keymem.key_mem[0][123] ),
    .QN(_00202_));
 DFFR_X1 \core.keymem.key_mem[0][124]$_DFFE_PN0P_  (.D(_00864_),
    .RN(net89),
    .CK(clknet_leaf_378_clk),
    .Q(\core.keymem.key_mem[0][124] ),
    .QN(_00207_));
 DFFR_X1 \core.keymem.key_mem[0][125]$_DFFE_PN0P_  (.D(_00865_),
    .RN(net89),
    .CK(clknet_leaf_379_clk),
    .Q(\core.keymem.key_mem[0][125] ),
    .QN(_00175_));
 DFFR_X1 \core.keymem.key_mem[0][126]$_DFFE_PN0P_  (.D(_00866_),
    .RN(net94),
    .CK(clknet_leaf_188_clk),
    .Q(\core.keymem.key_mem[0][126] ),
    .QN(_00188_));
 DFFR_X1 \core.keymem.key_mem[0][127]$_DFFE_PN0P_  (.D(_00867_),
    .RN(net93),
    .CK(clknet_leaf_373_clk),
    .Q(\core.keymem.key_mem[0][127] ),
    .QN(_00176_));
 DFFR_X1 \core.keymem.key_mem[0][12]$_DFFE_PN0P_  (.D(_00868_),
    .RN(net89),
    .CK(clknet_leaf_375_clk),
    .Q(\core.keymem.key_mem[0][12] ),
    .QN(_00246_));
 DFFR_X1 \core.keymem.key_mem[0][13]$_DFFE_PN0P_  (.D(_00869_),
    .RN(net85),
    .CK(clknet_leaf_52_clk),
    .Q(\core.keymem.key_mem[0][13] ),
    .QN(_00251_));
 DFFR_X1 \core.keymem.key_mem[0][14]$_DFFE_PN0P_  (.D(_00870_),
    .RN(net89),
    .CK(clknet_leaf_374_clk),
    .Q(\core.keymem.key_mem[0][14] ),
    .QN(_00252_));
 DFFR_X1 \core.keymem.key_mem[0][15]$_DFFE_PN0P_  (.D(_00871_),
    .RN(net89),
    .CK(clknet_leaf_380_clk),
    .Q(\core.keymem.key_mem[0][15] ),
    .QN(_00253_));
 DFFR_X1 \core.keymem.key_mem[0][16]$_DFFE_PN0P_  (.D(_00872_),
    .RN(net89),
    .CK(clknet_leaf_375_clk),
    .Q(\core.keymem.key_mem[0][16] ),
    .QN(_00254_));
 DFFR_X1 \core.keymem.key_mem[0][17]$_DFFE_PN0P_  (.D(_00873_),
    .RN(net89),
    .CK(clknet_leaf_375_clk),
    .Q(\core.keymem.key_mem[0][17] ),
    .QN(_00267_));
 DFFR_X1 \core.keymem.key_mem[0][18]$_DFFE_PN0P_  (.D(_00874_),
    .RN(net85),
    .CK(clknet_leaf_52_clk),
    .Q(\core.keymem.key_mem[0][18] ),
    .QN(_00275_));
 DFFR_X1 \core.keymem.key_mem[0][19]$_DFFE_PN0P_  (.D(_00875_),
    .RN(net85),
    .CK(clknet_leaf_52_clk),
    .Q(\core.keymem.key_mem[0][19] ),
    .QN(_00281_));
 DFFR_X2 \core.keymem.key_mem[0][1]$_DFFE_PN0P_  (.D(_00876_),
    .RN(net88),
    .CK(clknet_leaf_43_clk),
    .Q(\core.keymem.key_mem[0][1] ),
    .QN(_00187_));
 DFFR_X1 \core.keymem.key_mem[0][20]$_DFFE_PN0P_  (.D(_00877_),
    .RN(net89),
    .CK(clknet_leaf_381_clk),
    .Q(\core.keymem.key_mem[0][20] ),
    .QN(_00286_));
 DFFR_X1 \core.keymem.key_mem[0][21]$_DFFE_PN0P_  (.D(_00878_),
    .RN(net85),
    .CK(clknet_leaf_380_clk),
    .Q(\core.keymem.key_mem[0][21] ),
    .QN(_00291_));
 DFFR_X1 \core.keymem.key_mem[0][22]$_DFFE_PN0P_  (.D(_00879_),
    .RN(net93),
    .CK(clknet_leaf_373_clk),
    .Q(\core.keymem.key_mem[0][22] ),
    .QN(_00292_));
 DFFR_X1 \core.keymem.key_mem[0][23]$_DFFE_PN0P_  (.D(_00880_),
    .RN(net89),
    .CK(clknet_leaf_381_clk),
    .Q(\core.keymem.key_mem[0][23] ),
    .QN(_00293_));
 DFFR_X1 \core.keymem.key_mem[0][24]$_DFFE_PN0P_  (.D(_00881_),
    .RN(net85),
    .CK(clknet_leaf_51_clk),
    .Q(\core.keymem.key_mem[0][24] ),
    .QN(_00294_));
 DFFR_X1 \core.keymem.key_mem[0][25]$_DFFE_PN0P_  (.D(_00882_),
    .RN(net85),
    .CK(clknet_leaf_51_clk),
    .Q(\core.keymem.key_mem[0][25] ),
    .QN(_00298_));
 DFFR_X1 \core.keymem.key_mem[0][26]$_DFFE_PN0P_  (.D(_00883_),
    .RN(net88),
    .CK(clknet_leaf_44_clk),
    .Q(\core.keymem.key_mem[0][26] ),
    .QN(_00299_));
 DFFR_X1 \core.keymem.key_mem[0][27]$_DFFE_PN0P_  (.D(_00884_),
    .RN(net88),
    .CK(clknet_leaf_44_clk),
    .Q(\core.keymem.key_mem[0][27] ),
    .QN(_00300_));
 DFFR_X1 \core.keymem.key_mem[0][28]$_DFFE_PN0P_  (.D(_00885_),
    .RN(net87),
    .CK(clknet_leaf_32_clk),
    .Q(\core.keymem.key_mem[0][28] ),
    .QN(_00301_));
 DFFR_X1 \core.keymem.key_mem[0][29]$_DFFE_PN0P_  (.D(_00886_),
    .RN(net85),
    .CK(clknet_leaf_51_clk),
    .Q(\core.keymem.key_mem[0][29] ),
    .QN(_00295_));
 DFFR_X1 \core.keymem.key_mem[0][2]$_DFFE_PN0P_  (.D(_00887_),
    .RN(net85),
    .CK(clknet_leaf_51_clk),
    .Q(\core.keymem.key_mem[0][2] ),
    .QN(_00195_));
 DFFR_X1 \core.keymem.key_mem[0][30]$_DFFE_PN0P_  (.D(_00888_),
    .RN(net87),
    .CK(clknet_leaf_45_clk),
    .Q(\core.keymem.key_mem[0][30] ),
    .QN(_00296_));
 DFFR_X1 \core.keymem.key_mem[0][31]$_DFFE_PN0P_  (.D(_00889_),
    .RN(net87),
    .CK(clknet_leaf_32_clk),
    .Q(\core.keymem.key_mem[0][31] ),
    .QN(_00297_));
 DFFR_X2 \core.keymem.key_mem[0][32]$_DFFE_PN0P_  (.D(_00890_),
    .RN(net88),
    .CK(clknet_leaf_28_clk),
    .Q(\core.keymem.key_mem[0][32] ),
    .QN(_00265_));
 DFFR_X1 \core.keymem.key_mem[0][33]$_DFFE_PN0P_  (.D(_00891_),
    .RN(net88),
    .CK(clknet_leaf_31_clk),
    .Q(\core.keymem.key_mem[0][33] ),
    .QN(_00273_));
 DFFR_X1 \core.keymem.key_mem[0][34]$_DFFE_PN0P_  (.D(_00892_),
    .RN(net99),
    .CK(clknet_leaf_117_clk),
    .Q(\core.keymem.key_mem[0][34] ),
    .QN(_00279_));
 DFFR_X1 \core.keymem.key_mem[0][35]$_DFFE_PN0P_  (.D(_00893_),
    .RN(net89),
    .CK(clknet_leaf_25_clk),
    .Q(\core.keymem.key_mem[0][35] ),
    .QN(_00284_));
 DFFR_X1 \core.keymem.key_mem[0][36]$_DFFE_PN0P_  (.D(_00894_),
    .RN(net88),
    .CK(clknet_leaf_31_clk),
    .Q(\core.keymem.key_mem[0][36] ),
    .QN(_00289_));
 DFFR_X1 \core.keymem.key_mem[0][37]$_DFFE_PN0P_  (.D(_00895_),
    .RN(net88),
    .CK(clknet_leaf_90_clk),
    .Q(\core.keymem.key_mem[0][37] ),
    .QN(_00263_));
 DFFR_X1 \core.keymem.key_mem[0][38]$_DFFE_PN0P_  (.D(_00896_),
    .RN(net88),
    .CK(clknet_leaf_28_clk),
    .Q(\core.keymem.key_mem[0][38] ),
    .QN(_00264_));
 DFFR_X1 \core.keymem.key_mem[0][39]$_DFFE_PN0P_  (.D(_00897_),
    .RN(net88),
    .CK(clknet_leaf_45_clk),
    .Q(\core.keymem.key_mem[0][39] ),
    .QN(_00272_));
 DFFR_X1 \core.keymem.key_mem[0][3]$_DFFE_PN0P_  (.D(_00898_),
    .RN(net89),
    .CK(clknet_leaf_374_clk),
    .Q(\core.keymem.key_mem[0][3] ),
    .QN(_00201_));
 DFFR_X1 \core.keymem.key_mem[0][40]$_DFFE_PN0P_  (.D(_00899_),
    .RN(net88),
    .CK(clknet_leaf_46_clk),
    .Q(\core.keymem.key_mem[0][40] ),
    .QN(_00262_));
 DFFR_X1 \core.keymem.key_mem[0][41]$_DFFE_PN0P_  (.D(_00900_),
    .RN(net87),
    .CK(clknet_leaf_45_clk),
    .Q(\core.keymem.key_mem[0][41] ),
    .QN(_00271_));
 DFFR_X1 \core.keymem.key_mem[0][42]$_DFFE_PN0P_  (.D(_00901_),
    .RN(net88),
    .CK(clknet_leaf_45_clk),
    .Q(\core.keymem.key_mem[0][42] ),
    .QN(_00278_));
 DFFR_X1 \core.keymem.key_mem[0][43]$_DFFE_PN0P_  (.D(_00902_),
    .RN(net88),
    .CK(clknet_leaf_46_clk),
    .Q(\core.keymem.key_mem[0][43] ),
    .QN(_00283_));
 DFFR_X1 \core.keymem.key_mem[0][44]$_DFFE_PN0P_  (.D(_00903_),
    .RN(net99),
    .CK(clknet_leaf_115_clk),
    .Q(\core.keymem.key_mem[0][44] ),
    .QN(_00288_));
 DFFR_X1 \core.keymem.key_mem[0][45]$_DFFE_PN0P_  (.D(_00904_),
    .RN(net85),
    .CK(clknet_leaf_48_clk),
    .Q(\core.keymem.key_mem[0][45] ),
    .QN(_00260_));
 DFFR_X1 \core.keymem.key_mem[0][46]$_DFFE_PN0P_  (.D(_00905_),
    .RN(net88),
    .CK(clknet_leaf_30_clk),
    .Q(\core.keymem.key_mem[0][46] ),
    .QN(_00270_));
 DFFR_X1 \core.keymem.key_mem[0][47]$_DFFE_PN0P_  (.D(_00906_),
    .RN(net98),
    .CK(clknet_leaf_180_clk),
    .Q(\core.keymem.key_mem[0][47] ),
    .QN(_00261_));
 DFFR_X1 \core.keymem.key_mem[0][48]$_DFFE_PN0P_  (.D(_00907_),
    .RN(net95),
    .CK(clknet_leaf_119_clk),
    .Q(\core.keymem.key_mem[0][48] ),
    .QN(_00266_));
 DFFR_X1 \core.keymem.key_mem[0][49]$_DFFE_PN0P_  (.D(_00908_),
    .RN(net88),
    .CK(clknet_leaf_46_clk),
    .Q(\core.keymem.key_mem[0][49] ),
    .QN(_00274_));
 DFFR_X1 \core.keymem.key_mem[0][4]$_DFFE_PN0P_  (.D(_00909_),
    .RN(net87),
    .CK(clknet_leaf_36_clk),
    .Q(\core.keymem.key_mem[0][4] ),
    .QN(_00206_));
 DFFR_X1 \core.keymem.key_mem[0][50]$_DFFE_PN0P_  (.D(_00910_),
    .RN(net88),
    .CK(clknet_leaf_45_clk),
    .Q(\core.keymem.key_mem[0][50] ),
    .QN(_00280_));
 DFFR_X1 \core.keymem.key_mem[0][51]$_DFFE_PN0P_  (.D(_00911_),
    .RN(net87),
    .CK(clknet_leaf_37_clk),
    .Q(\core.keymem.key_mem[0][51] ),
    .QN(_00285_));
 DFFR_X1 \core.keymem.key_mem[0][52]$_DFFE_PN0P_  (.D(_00912_),
    .RN(net99),
    .CK(clknet_leaf_70_clk),
    .Q(\core.keymem.key_mem[0][52] ),
    .QN(_00290_));
 DFFR_X1 \core.keymem.key_mem[0][53]$_DFFE_PN0P_  (.D(_00913_),
    .RN(net85),
    .CK(clknet_leaf_50_clk),
    .Q(\core.keymem.key_mem[0][53] ),
    .QN(_00257_));
 DFFR_X1 \core.keymem.key_mem[0][54]$_DFFE_PN0P_  (.D(_00914_),
    .RN(net88),
    .CK(clknet_leaf_46_clk),
    .Q(\core.keymem.key_mem[0][54] ),
    .QN(_00258_));
 DFFR_X1 \core.keymem.key_mem[0][55]$_DFFE_PN0P_  (.D(_00915_),
    .RN(net85),
    .CK(clknet_leaf_51_clk),
    .Q(\core.keymem.key_mem[0][55] ),
    .QN(_00259_));
 DFFR_X1 \core.keymem.key_mem[0][56]$_DFFE_PN0P_  (.D(_00916_),
    .RN(net88),
    .CK(clknet_leaf_44_clk),
    .Q(\core.keymem.key_mem[0][56] ),
    .QN(_00256_));
 DFFR_X1 \core.keymem.key_mem[0][57]$_DFFE_PN0P_  (.D(_00917_),
    .RN(net85),
    .CK(clknet_leaf_44_clk),
    .Q(\core.keymem.key_mem[0][57] ),
    .QN(_00269_));
 DFFR_X1 \core.keymem.key_mem[0][58]$_DFFE_PN0P_  (.D(_00918_),
    .RN(net87),
    .CK(clknet_leaf_45_clk),
    .Q(\core.keymem.key_mem[0][58] ),
    .QN(_00277_));
 DFFR_X1 \core.keymem.key_mem[0][59]$_DFFE_PN0P_  (.D(_00919_),
    .RN(net87),
    .CK(clknet_leaf_32_clk),
    .Q(\core.keymem.key_mem[0][59] ),
    .QN(_00282_));
 DFFR_X1 \core.keymem.key_mem[0][5]$_DFFE_PN0P_  (.D(_00920_),
    .RN(net100),
    .CK(clknet_leaf_21_clk),
    .Q(\core.keymem.key_mem[0][5] ),
    .QN(_00211_));
 DFFR_X1 \core.keymem.key_mem[0][60]$_DFFE_PN0P_  (.D(_00921_),
    .RN(net82),
    .CK(clknet_leaf_10_clk),
    .Q(\core.keymem.key_mem[0][60] ),
    .QN(_00287_));
 DFFR_X2 \core.keymem.key_mem[0][61]$_DFFE_PN0P_  (.D(_00922_),
    .RN(net82),
    .CK(clknet_leaf_35_clk),
    .Q(\core.keymem.key_mem[0][61] ),
    .QN(_00255_));
 DFFR_X1 \core.keymem.key_mem[0][62]$_DFFE_PN0P_  (.D(_00923_),
    .RN(net88),
    .CK(clknet_leaf_45_clk),
    .Q(\core.keymem.key_mem[0][62] ),
    .QN(_00268_));
 DFFR_X1 \core.keymem.key_mem[0][63]$_DFFE_PN0P_  (.D(_00924_),
    .RN(net82),
    .CK(clknet_leaf_10_clk),
    .Q(\core.keymem.key_mem[0][63] ),
    .QN(_00276_));
 DFFR_X1 \core.keymem.key_mem[0][64]$_DFFE_PN0P_  (.D(_00925_),
    .RN(net82),
    .CK(clknet_leaf_23_clk),
    .Q(\core.keymem.key_mem[0][64] ),
    .QN(_00225_));
 DFFR_X1 \core.keymem.key_mem[0][65]$_DFFE_PN0P_  (.D(_00926_),
    .RN(net87),
    .CK(clknet_leaf_36_clk),
    .Q(\core.keymem.key_mem[0][65] ),
    .QN(_00233_));
 DFFR_X1 \core.keymem.key_mem[0][66]$_DFFE_PN0P_  (.D(_00927_),
    .RN(net82),
    .CK(clknet_leaf_10_clk),
    .Q(\core.keymem.key_mem[0][66] ),
    .QN(_00239_));
 DFFR_X1 \core.keymem.key_mem[0][67]$_DFFE_PN0P_  (.D(_00928_),
    .RN(net82),
    .CK(clknet_leaf_35_clk),
    .Q(\core.keymem.key_mem[0][67] ),
    .QN(_00244_));
 DFFR_X1 \core.keymem.key_mem[0][68]$_DFFE_PN0P_  (.D(_00929_),
    .RN(net95),
    .CK(clknet_leaf_77_clk),
    .Q(\core.keymem.key_mem[0][68] ),
    .QN(_00249_));
 DFFR_X1 \core.keymem.key_mem[0][69]$_DFFE_PN0P_  (.D(_00930_),
    .RN(net88),
    .CK(clknet_leaf_44_clk),
    .Q(\core.keymem.key_mem[0][69] ),
    .QN(_00223_));
 DFFR_X1 \core.keymem.key_mem[0][6]$_DFFE_PN0P_  (.D(_00931_),
    .RN(net85),
    .CK(clknet_leaf_52_clk),
    .Q(\core.keymem.key_mem[0][6] ),
    .QN(_00212_));
 DFFR_X1 \core.keymem.key_mem[0][70]$_DFFE_PN0P_  (.D(_00932_),
    .RN(net88),
    .CK(clknet_leaf_30_clk),
    .Q(\core.keymem.key_mem[0][70] ),
    .QN(_00232_));
 DFFR_X1 \core.keymem.key_mem[0][71]$_DFFE_PN0P_  (.D(_00933_),
    .RN(net99),
    .CK(clknet_leaf_70_clk),
    .Q(\core.keymem.key_mem[0][71] ),
    .QN(_00224_));
 DFFR_X1 \core.keymem.key_mem[0][72]$_DFFE_PN0P_  (.D(_00934_),
    .RN(net95),
    .CK(clknet_leaf_76_clk),
    .Q(\core.keymem.key_mem[0][72] ),
    .QN(_00226_));
 DFFR_X1 \core.keymem.key_mem[0][73]$_DFFE_PN0P_  (.D(_00935_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[0][73] ),
    .QN(_00234_));
 DFFR_X1 \core.keymem.key_mem[0][74]$_DFFE_PN0P_  (.D(_00936_),
    .RN(net93),
    .CK(clknet_leaf_373_clk),
    .Q(\core.keymem.key_mem[0][74] ),
    .QN(_00240_));
 DFFR_X1 \core.keymem.key_mem[0][75]$_DFFE_PN0P_  (.D(_00937_),
    .RN(net85),
    .CK(clknet_leaf_382_clk),
    .Q(\core.keymem.key_mem[0][75] ),
    .QN(_00245_));
 DFFR_X1 \core.keymem.key_mem[0][76]$_DFFE_PN0P_  (.D(_00938_),
    .RN(net89),
    .CK(clknet_leaf_374_clk),
    .Q(\core.keymem.key_mem[0][76] ),
    .QN(_00250_));
 DFFR_X2 \core.keymem.key_mem[0][77]$_DFFE_PN0P_  (.D(_00939_),
    .RN(net89),
    .CK(clknet_leaf_381_clk),
    .Q(\core.keymem.key_mem[0][77] ),
    .QN(_00220_));
 DFFR_X1 \core.keymem.key_mem[0][78]$_DFFE_PN0P_  (.D(_00940_),
    .RN(net98),
    .CK(clknet_leaf_170_clk),
    .Q(\core.keymem.key_mem[0][78] ),
    .QN(_00221_));
 DFFR_X2 \core.keymem.key_mem[0][79]$_DFFE_PN0P_  (.D(_00941_),
    .RN(net93),
    .CK(clknet_leaf_376_clk),
    .Q(\core.keymem.key_mem[0][79] ),
    .QN(_00222_));
 DFFR_X1 \core.keymem.key_mem[0][7]$_DFFE_PN0P_  (.D(_00942_),
    .RN(net88),
    .CK(clknet_leaf_42_clk),
    .Q(\core.keymem.key_mem[0][7] ),
    .QN(_00213_));
 DFFR_X1 \core.keymem.key_mem[0][80]$_DFFE_PN0P_  (.D(_00943_),
    .RN(net85),
    .CK(clknet_leaf_53_clk),
    .Q(\core.keymem.key_mem[0][80] ),
    .QN(_00219_));
 DFFR_X1 \core.keymem.key_mem[0][81]$_DFFE_PN0P_  (.D(_00944_),
    .RN(net89),
    .CK(clknet_leaf_374_clk),
    .Q(\core.keymem.key_mem[0][81] ),
    .QN(_00231_));
 DFFR_X1 \core.keymem.key_mem[0][82]$_DFFE_PN0P_  (.D(_00945_),
    .RN(net85),
    .CK(clknet_leaf_52_clk),
    .Q(\core.keymem.key_mem[0][82] ),
    .QN(_00238_));
 DFFR_X1 \core.keymem.key_mem[0][83]$_DFFE_PN0P_  (.D(_00946_),
    .RN(net85),
    .CK(clknet_leaf_43_clk),
    .Q(\core.keymem.key_mem[0][83] ),
    .QN(_00243_));
 DFFR_X1 \core.keymem.key_mem[0][84]$_DFFE_PN0P_  (.D(_00947_),
    .RN(net95),
    .CK(clknet_leaf_72_clk),
    .Q(\core.keymem.key_mem[0][84] ),
    .QN(_00248_));
 DFFR_X1 \core.keymem.key_mem[0][85]$_DFFE_PN0P_  (.D(_00948_),
    .RN(net89),
    .CK(clknet_leaf_371_clk),
    .Q(\core.keymem.key_mem[0][85] ),
    .QN(_00218_));
 DFFR_X1 \core.keymem.key_mem[0][86]$_DFFE_PN0P_  (.D(_00949_),
    .RN(net95),
    .CK(clknet_leaf_208_clk),
    .Q(\core.keymem.key_mem[0][86] ),
    .QN(_00230_));
 DFFR_X1 \core.keymem.key_mem[0][87]$_DFFE_PN0P_  (.D(_00950_),
    .RN(net89),
    .CK(clknet_leaf_379_clk),
    .Q(\core.keymem.key_mem[0][87] ),
    .QN(_00237_));
 DFFR_X1 \core.keymem.key_mem[0][88]$_DFFE_PN0P_  (.D(_00951_),
    .RN(net93),
    .CK(clknet_leaf_376_clk),
    .Q(\core.keymem.key_mem[0][88] ),
    .QN(_00217_));
 DFFR_X1 \core.keymem.key_mem[0][89]$_DFFE_PN0P_  (.D(_00952_),
    .RN(net93),
    .CK(clknet_leaf_376_clk),
    .Q(\core.keymem.key_mem[0][89] ),
    .QN(_00229_));
 DFFR_X1 \core.keymem.key_mem[0][8]$_DFFE_PN0P_  (.D(_00953_),
    .RN(net89),
    .CK(clknet_leaf_375_clk),
    .Q(\core.keymem.key_mem[0][8] ),
    .QN(_00214_));
 DFFR_X1 \core.keymem.key_mem[0][90]$_DFFE_PN0P_  (.D(_00954_),
    .RN(net89),
    .CK(clknet_leaf_53_clk),
    .Q(\core.keymem.key_mem[0][90] ),
    .QN(_00236_));
 DFFR_X1 \core.keymem.key_mem[0][91]$_DFFE_PN0P_  (.D(_00955_),
    .RN(net85),
    .CK(clknet_leaf_52_clk),
    .Q(\core.keymem.key_mem[0][91] ),
    .QN(_00242_));
 DFFR_X1 \core.keymem.key_mem[0][92]$_DFFE_PN0P_  (.D(_00956_),
    .RN(net85),
    .CK(clknet_leaf_51_clk),
    .Q(\core.keymem.key_mem[0][92] ),
    .QN(_00247_));
 DFFR_X1 \core.keymem.key_mem[0][93]$_DFFE_PN0P_  (.D(_00957_),
    .RN(net89),
    .CK(clknet_leaf_379_clk),
    .Q(\core.keymem.key_mem[0][93] ),
    .QN(_00215_));
 DFFR_X1 \core.keymem.key_mem[0][94]$_DFFE_PN0P_  (.D(_00958_),
    .RN(net91),
    .CK(clknet_leaf_285_clk),
    .Q(\core.keymem.key_mem[0][94] ),
    .QN(_00216_));
 DFFR_X1 \core.keymem.key_mem[0][95]$_DFFE_PN0P_  (.D(_00959_),
    .RN(net91),
    .CK(clknet_leaf_285_clk),
    .Q(\core.keymem.key_mem[0][95] ),
    .QN(_00228_));
 DFFR_X2 \core.keymem.key_mem[0][96]$_DFFE_PN0P_  (.D(_00960_),
    .RN(net93),
    .CK(clknet_leaf_374_clk),
    .Q(\core.keymem.key_mem[0][96] ),
    .QN(_00186_));
 DFFR_X1 \core.keymem.key_mem[0][97]$_DFFE_PN0P_  (.D(_00961_),
    .RN(net93),
    .CK(clknet_leaf_192_clk),
    .Q(\core.keymem.key_mem[0][97] ),
    .QN(_00194_));
 DFFR_X1 \core.keymem.key_mem[0][98]$_DFFE_PN0P_  (.D(_00962_),
    .RN(net91),
    .CK(clknet_leaf_284_clk),
    .Q(\core.keymem.key_mem[0][98] ),
    .QN(_00200_));
 DFFR_X1 \core.keymem.key_mem[0][99]$_DFFE_PN0P_  (.D(_00963_),
    .RN(net93),
    .CK(clknet_leaf_376_clk),
    .Q(\core.keymem.key_mem[0][99] ),
    .QN(_00205_));
 DFFR_X1 \core.keymem.key_mem[0][9]$_DFFE_PN0P_  (.D(_00964_),
    .RN(net89),
    .CK(clknet_leaf_379_clk),
    .Q(\core.keymem.key_mem[0][9] ),
    .QN(_00227_));
 DFFR_X1 \core.keymem.key_mem[10][0]$_DFFE_PN0P_  (.D(_00965_),
    .RN(net96),
    .CK(clknet_leaf_221_clk),
    .Q(\core.keymem.key_mem[10][0] ),
    .QN(_21639_));
 DFFR_X1 \core.keymem.key_mem[10][100]$_DFFE_PN0P_  (.D(_00966_),
    .RN(net94),
    .CK(clknet_leaf_210_clk),
    .Q(\core.keymem.key_mem[10][100] ),
    .QN(_21638_));
 DFFR_X1 \core.keymem.key_mem[10][101]$_DFFE_PN0P_  (.D(_00967_),
    .RN(net96),
    .CK(clknet_leaf_223_clk),
    .Q(\core.keymem.key_mem[10][101] ),
    .QN(_21637_));
 DFFR_X1 \core.keymem.key_mem[10][102]$_DFFE_PN0P_  (.D(_00968_),
    .RN(net96),
    .CK(clknet_leaf_232_clk),
    .Q(\core.keymem.key_mem[10][102] ),
    .QN(_21636_));
 DFFR_X1 \core.keymem.key_mem[10][103]$_DFFE_PN0P_  (.D(_00969_),
    .RN(net96),
    .CK(clknet_leaf_246_clk),
    .Q(\core.keymem.key_mem[10][103] ),
    .QN(_21635_));
 DFFR_X1 \core.keymem.key_mem[10][104]$_DFFE_PN0P_  (.D(_00970_),
    .RN(net93),
    .CK(clknet_leaf_193_clk),
    .Q(\core.keymem.key_mem[10][104] ),
    .QN(_21634_));
 DFFR_X1 \core.keymem.key_mem[10][105]$_DFFE_PN0P_  (.D(_00971_),
    .RN(net96),
    .CK(clknet_leaf_247_clk),
    .Q(\core.keymem.key_mem[10][105] ),
    .QN(_21633_));
 DFFR_X1 \core.keymem.key_mem[10][106]$_DFFE_PN0P_  (.D(_00972_),
    .RN(net92),
    .CK(clknet_leaf_258_clk),
    .Q(\core.keymem.key_mem[10][106] ),
    .QN(_21632_));
 DFFR_X1 \core.keymem.key_mem[10][107]$_DFFE_PN0P_  (.D(_00973_),
    .RN(net92),
    .CK(clknet_leaf_270_clk),
    .Q(\core.keymem.key_mem[10][107] ),
    .QN(_21631_));
 DFFR_X1 \core.keymem.key_mem[10][108]$_DFFE_PN0P_  (.D(_00974_),
    .RN(net91),
    .CK(clknet_leaf_280_clk),
    .Q(\core.keymem.key_mem[10][108] ),
    .QN(_21630_));
 DFFR_X1 \core.keymem.key_mem[10][109]$_DFFE_PN0P_  (.D(_00975_),
    .RN(net94),
    .CK(clknet_leaf_259_clk),
    .Q(\core.keymem.key_mem[10][109] ),
    .QN(_21629_));
 DFFR_X1 \core.keymem.key_mem[10][10]$_DFFE_PN0P_  (.D(_00976_),
    .RN(net94),
    .CK(clknet_leaf_187_clk),
    .Q(\core.keymem.key_mem[10][10] ),
    .QN(_21628_));
 DFFR_X1 \core.keymem.key_mem[10][110]$_DFFE_PN0P_  (.D(_00977_),
    .RN(net96),
    .CK(clknet_leaf_250_clk),
    .Q(\core.keymem.key_mem[10][110] ),
    .QN(_21627_));
 DFFR_X1 \core.keymem.key_mem[10][111]$_DFFE_PN0P_  (.D(_00978_),
    .RN(net96),
    .CK(clknet_leaf_227_clk),
    .Q(\core.keymem.key_mem[10][111] ),
    .QN(_21626_));
 DFFR_X1 \core.keymem.key_mem[10][112]$_DFFE_PN0P_  (.D(_00979_),
    .RN(net94),
    .CK(clknet_leaf_260_clk),
    .Q(\core.keymem.key_mem[10][112] ),
    .QN(_21625_));
 DFFR_X1 \core.keymem.key_mem[10][113]$_DFFE_PN0P_  (.D(_00980_),
    .RN(net91),
    .CK(clknet_leaf_273_clk),
    .Q(\core.keymem.key_mem[10][113] ),
    .QN(_21624_));
 DFFR_X1 \core.keymem.key_mem[10][114]$_DFFE_PN0P_  (.D(_00981_),
    .RN(net91),
    .CK(clknet_leaf_274_clk),
    .Q(\core.keymem.key_mem[10][114] ),
    .QN(_21623_));
 DFFR_X1 \core.keymem.key_mem[10][115]$_DFFE_PN0P_  (.D(_00982_),
    .RN(net92),
    .CK(clknet_leaf_275_clk),
    .Q(\core.keymem.key_mem[10][115] ),
    .QN(_21622_));
 DFFR_X1 \core.keymem.key_mem[10][116]$_DFFE_PN0P_  (.D(_00983_),
    .RN(net94),
    .CK(clknet_leaf_263_clk),
    .Q(\core.keymem.key_mem[10][116] ),
    .QN(_21621_));
 DFFR_X1 \core.keymem.key_mem[10][117]$_DFFE_PN0P_  (.D(_00984_),
    .RN(net96),
    .CK(clknet_leaf_226_clk),
    .Q(\core.keymem.key_mem[10][117] ),
    .QN(_21620_));
 DFFR_X1 \core.keymem.key_mem[10][118]$_DFFE_PN0P_  (.D(_00985_),
    .RN(net97),
    .CK(clknet_leaf_242_clk),
    .Q(\core.keymem.key_mem[10][118] ),
    .QN(_21619_));
 DFFR_X1 \core.keymem.key_mem[10][119]$_DFFE_PN0P_  (.D(_00986_),
    .RN(net94),
    .CK(clknet_leaf_262_clk),
    .Q(\core.keymem.key_mem[10][119] ),
    .QN(_21618_));
 DFFR_X1 \core.keymem.key_mem[10][11]$_DFFE_PN0P_  (.D(_00987_),
    .RN(net95),
    .CK(clknet_leaf_60_clk),
    .Q(\core.keymem.key_mem[10][11] ),
    .QN(_21617_));
 DFFR_X1 \core.keymem.key_mem[10][120]$_DFFE_PN0P_  (.D(_00988_),
    .RN(net94),
    .CK(clknet_leaf_205_clk),
    .Q(\core.keymem.key_mem[10][120] ),
    .QN(_21616_));
 DFFR_X1 \core.keymem.key_mem[10][121]$_DFFE_PN0P_  (.D(_00989_),
    .RN(net94),
    .CK(clknet_leaf_264_clk),
    .Q(\core.keymem.key_mem[10][121] ),
    .QN(_21615_));
 DFFR_X1 \core.keymem.key_mem[10][122]$_DFFE_PN0P_  (.D(_00990_),
    .RN(net97),
    .CK(clknet_leaf_237_clk),
    .Q(\core.keymem.key_mem[10][122] ),
    .QN(_21614_));
 DFFR_X1 \core.keymem.key_mem[10][123]$_DFFE_PN0P_  (.D(_00991_),
    .RN(net93),
    .CK(clknet_leaf_197_clk),
    .Q(\core.keymem.key_mem[10][123] ),
    .QN(_21613_));
 DFFR_X1 \core.keymem.key_mem[10][124]$_DFFE_PN0P_  (.D(_00992_),
    .RN(net93),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[10][124] ),
    .QN(_21612_));
 DFFR_X1 \core.keymem.key_mem[10][125]$_DFFE_PN0P_  (.D(_00993_),
    .RN(net97),
    .CK(clknet_leaf_236_clk),
    .Q(\core.keymem.key_mem[10][125] ),
    .QN(_21611_));
 DFFR_X1 \core.keymem.key_mem[10][126]$_DFFE_PN0P_  (.D(_00994_),
    .RN(net98),
    .CK(clknet_leaf_166_clk),
    .Q(\core.keymem.key_mem[10][126] ),
    .QN(_21610_));
 DFFR_X1 \core.keymem.key_mem[10][127]$_DFFE_PN0P_  (.D(_00995_),
    .RN(net97),
    .CK(clknet_leaf_241_clk),
    .Q(\core.keymem.key_mem[10][127] ),
    .QN(_21609_));
 DFFR_X1 \core.keymem.key_mem[10][12]$_DFFE_PN0P_  (.D(_00996_),
    .RN(net93),
    .CK(clknet_leaf_208_clk),
    .Q(\core.keymem.key_mem[10][12] ),
    .QN(_21608_));
 DFFR_X1 \core.keymem.key_mem[10][13]$_DFFE_PN0P_  (.D(_00997_),
    .RN(net87),
    .CK(clknet_leaf_32_clk),
    .Q(\core.keymem.key_mem[10][13] ),
    .QN(_21607_));
 DFFR_X1 \core.keymem.key_mem[10][14]$_DFFE_PN0P_  (.D(_00998_),
    .RN(net94),
    .CK(clknet_leaf_211_clk),
    .Q(\core.keymem.key_mem[10][14] ),
    .QN(_21606_));
 DFFR_X1 \core.keymem.key_mem[10][15]$_DFFE_PN0P_  (.D(_00999_),
    .RN(net96),
    .CK(clknet_leaf_165_clk),
    .Q(\core.keymem.key_mem[10][15] ),
    .QN(_21605_));
 DFFR_X1 \core.keymem.key_mem[10][16]$_DFFE_PN0P_  (.D(_01000_),
    .RN(net89),
    .CK(clknet_leaf_34_clk),
    .Q(\core.keymem.key_mem[10][16] ),
    .QN(_21604_));
 DFFR_X1 \core.keymem.key_mem[10][17]$_DFFE_PN0P_  (.D(_01001_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[10][17] ),
    .QN(_21603_));
 DFFR_X1 \core.keymem.key_mem[10][18]$_DFFE_PN0P_  (.D(_01002_),
    .RN(net89),
    .CK(clknet_leaf_26_clk),
    .Q(\core.keymem.key_mem[10][18] ),
    .QN(_21602_));
 DFFR_X1 \core.keymem.key_mem[10][19]$_DFFE_PN0P_  (.D(_01003_),
    .RN(net85),
    .CK(clknet_leaf_54_clk),
    .Q(\core.keymem.key_mem[10][19] ),
    .QN(_21601_));
 DFFR_X1 \core.keymem.key_mem[10][1]$_DFFE_PN0P_  (.D(_01004_),
    .RN(net89),
    .CK(clknet_leaf_21_clk),
    .Q(\core.keymem.key_mem[10][1] ),
    .QN(_21600_));
 DFFR_X1 \core.keymem.key_mem[10][20]$_DFFE_PN0P_  (.D(_01005_),
    .RN(net89),
    .CK(clknet_leaf_96_clk),
    .Q(\core.keymem.key_mem[10][20] ),
    .QN(_21599_));
 DFFR_X1 \core.keymem.key_mem[10][21]$_DFFE_PN0P_  (.D(_01006_),
    .RN(net85),
    .CK(clknet_leaf_66_clk),
    .Q(\core.keymem.key_mem[10][21] ),
    .QN(_21598_));
 DFFR_X1 \core.keymem.key_mem[10][22]$_DFFE_PN0P_  (.D(_01007_),
    .RN(net96),
    .CK(clknet_leaf_222_clk),
    .Q(\core.keymem.key_mem[10][22] ),
    .QN(_21597_));
 DFFR_X1 \core.keymem.key_mem[10][23]$_DFFE_PN0P_  (.D(_01008_),
    .RN(net89),
    .CK(clknet_leaf_55_clk),
    .Q(\core.keymem.key_mem[10][23] ),
    .QN(_21596_));
 DFFR_X1 \core.keymem.key_mem[10][24]$_DFFE_PN0P_  (.D(_01009_),
    .RN(net85),
    .CK(clknet_leaf_49_clk),
    .Q(\core.keymem.key_mem[10][24] ),
    .QN(_21595_));
 DFFR_X1 \core.keymem.key_mem[10][25]$_DFFE_PN0P_  (.D(_01010_),
    .RN(net85),
    .CK(clknet_leaf_48_clk),
    .Q(\core.keymem.key_mem[10][25] ),
    .QN(_21594_));
 DFFR_X1 \core.keymem.key_mem[10][26]$_DFFE_PN0P_  (.D(_01011_),
    .RN(net100),
    .CK(clknet_leaf_97_clk),
    .Q(\core.keymem.key_mem[10][26] ),
    .QN(_21593_));
 DFFR_X1 \core.keymem.key_mem[10][27]$_DFFE_PN0P_  (.D(_01012_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[10][27] ),
    .QN(_21592_));
 DFFR_X1 \core.keymem.key_mem[10][28]$_DFFE_PN0P_  (.D(_01013_),
    .RN(net16),
    .CK(clknet_leaf_131_clk),
    .Q(\core.keymem.key_mem[10][28] ),
    .QN(_21591_));
 DFFR_X1 \core.keymem.key_mem[10][29]$_DFFE_PN0P_  (.D(_01014_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[10][29] ),
    .QN(_21590_));
 DFFR_X1 \core.keymem.key_mem[10][2]$_DFFE_PN0P_  (.D(_01015_),
    .RN(net95),
    .CK(clknet_leaf_60_clk),
    .Q(\core.keymem.key_mem[10][2] ),
    .QN(_21589_));
 DFFR_X1 \core.keymem.key_mem[10][30]$_DFFE_PN0P_  (.D(_01016_),
    .RN(net98),
    .CK(clknet_leaf_149_clk),
    .Q(\core.keymem.key_mem[10][30] ),
    .QN(_21588_));
 DFFR_X1 \core.keymem.key_mem[10][31]$_DFFE_PN0P_  (.D(_01017_),
    .RN(net98),
    .CK(clknet_leaf_143_clk),
    .Q(\core.keymem.key_mem[10][31] ),
    .QN(_21587_));
 DFFR_X1 \core.keymem.key_mem[10][32]$_DFFE_PN0P_  (.D(_01018_),
    .RN(net100),
    .CK(clknet_leaf_113_clk),
    .Q(\core.keymem.key_mem[10][32] ),
    .QN(_21586_));
 DFFR_X1 \core.keymem.key_mem[10][33]$_DFFE_PN0P_  (.D(_01019_),
    .RN(net16),
    .CK(clknet_leaf_126_clk),
    .Q(\core.keymem.key_mem[10][33] ),
    .QN(_21585_));
 DFFR_X1 \core.keymem.key_mem[10][34]$_DFFE_PN0P_  (.D(_01020_),
    .RN(net16),
    .CK(clknet_leaf_136_clk),
    .Q(\core.keymem.key_mem[10][34] ),
    .QN(_21584_));
 DFFR_X1 \core.keymem.key_mem[10][35]$_DFFE_PN0P_  (.D(_01021_),
    .RN(net99),
    .CK(clknet_leaf_128_clk),
    .Q(\core.keymem.key_mem[10][35] ),
    .QN(_21583_));
 DFFR_X1 \core.keymem.key_mem[10][36]$_DFFE_PN0P_  (.D(_01022_),
    .RN(net88),
    .CK(clknet_leaf_89_clk),
    .Q(\core.keymem.key_mem[10][36] ),
    .QN(_21582_));
 DFFR_X1 \core.keymem.key_mem[10][37]$_DFFE_PN0P_  (.D(_01023_),
    .RN(net88),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[10][37] ),
    .QN(_21581_));
 DFFR_X1 \core.keymem.key_mem[10][38]$_DFFE_PN0P_  (.D(_01024_),
    .RN(net16),
    .CK(clknet_leaf_124_clk),
    .Q(\core.keymem.key_mem[10][38] ),
    .QN(_21580_));
 DFFR_X1 \core.keymem.key_mem[10][39]$_DFFE_PN0P_  (.D(_01025_),
    .RN(net85),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[10][39] ),
    .QN(_21579_));
 DFFR_X1 \core.keymem.key_mem[10][3]$_DFFE_PN0P_  (.D(_01026_),
    .RN(net88),
    .CK(clknet_leaf_27_clk),
    .Q(\core.keymem.key_mem[10][3] ),
    .QN(_21578_));
 DFFR_X1 \core.keymem.key_mem[10][40]$_DFFE_PN0P_  (.D(_01027_),
    .RN(net88),
    .CK(clknet_leaf_90_clk),
    .Q(\core.keymem.key_mem[10][40] ),
    .QN(_21577_));
 DFFR_X1 \core.keymem.key_mem[10][41]$_DFFE_PN0P_  (.D(_01028_),
    .RN(net99),
    .CK(clknet_leaf_115_clk),
    .Q(\core.keymem.key_mem[10][41] ),
    .QN(_21576_));
 DFFR_X1 \core.keymem.key_mem[10][42]$_DFFE_PN0P_  (.D(_01029_),
    .RN(net100),
    .CK(clknet_leaf_129_clk),
    .Q(\core.keymem.key_mem[10][42] ),
    .QN(_21575_));
 DFFR_X1 \core.keymem.key_mem[10][43]$_DFFE_PN0P_  (.D(_01030_),
    .RN(net85),
    .CK(clknet_leaf_88_clk),
    .Q(\core.keymem.key_mem[10][43] ),
    .QN(_21574_));
 DFFR_X1 \core.keymem.key_mem[10][44]$_DFFE_PN0P_  (.D(_01031_),
    .RN(net100),
    .CK(clknet_leaf_113_clk),
    .Q(\core.keymem.key_mem[10][44] ),
    .QN(_21573_));
 DFFR_X1 \core.keymem.key_mem[10][45]$_DFFE_PN0P_  (.D(_01032_),
    .RN(net99),
    .CK(clknet_leaf_69_clk),
    .Q(\core.keymem.key_mem[10][45] ),
    .QN(_21572_));
 DFFR_X1 \core.keymem.key_mem[10][46]$_DFFE_PN0P_  (.D(_01033_),
    .RN(net99),
    .CK(clknet_leaf_85_clk),
    .Q(\core.keymem.key_mem[10][46] ),
    .QN(_21571_));
 DFFR_X1 \core.keymem.key_mem[10][47]$_DFFE_PN0P_  (.D(_01034_),
    .RN(net98),
    .CK(clknet_leaf_146_clk),
    .Q(\core.keymem.key_mem[10][47] ),
    .QN(_21570_));
 DFFR_X1 \core.keymem.key_mem[10][48]$_DFFE_PN0P_  (.D(_01035_),
    .RN(net95),
    .CK(clknet_leaf_119_clk),
    .Q(\core.keymem.key_mem[10][48] ),
    .QN(_21569_));
 DFFR_X1 \core.keymem.key_mem[10][49]$_DFFE_PN0P_  (.D(_01036_),
    .RN(net99),
    .CK(clknet_leaf_78_clk),
    .Q(\core.keymem.key_mem[10][49] ),
    .QN(_21568_));
 DFFR_X1 \core.keymem.key_mem[10][4]$_DFFE_PN0P_  (.D(_01037_),
    .RN(net100),
    .CK(clknet_leaf_106_clk),
    .Q(\core.keymem.key_mem[10][4] ),
    .QN(_21567_));
 DFFR_X1 \core.keymem.key_mem[10][50]$_DFFE_PN0P_  (.D(_01038_),
    .RN(net98),
    .CK(clknet_leaf_137_clk),
    .Q(\core.keymem.key_mem[10][50] ),
    .QN(_21566_));
 DFFR_X1 \core.keymem.key_mem[10][51]$_DFFE_PN0P_  (.D(_01039_),
    .RN(net99),
    .CK(clknet_leaf_128_clk),
    .Q(\core.keymem.key_mem[10][51] ),
    .QN(_21565_));
 DFFR_X1 \core.keymem.key_mem[10][52]$_DFFE_PN0P_  (.D(_01040_),
    .RN(net99),
    .CK(clknet_leaf_80_clk),
    .Q(\core.keymem.key_mem[10][52] ),
    .QN(_21564_));
 DFFR_X1 \core.keymem.key_mem[10][53]$_DFFE_PN0P_  (.D(_01041_),
    .RN(net98),
    .CK(clknet_leaf_172_clk),
    .Q(\core.keymem.key_mem[10][53] ),
    .QN(_21563_));
 DFFR_X1 \core.keymem.key_mem[10][54]$_DFFE_PN0P_  (.D(_01042_),
    .RN(net98),
    .CK(clknet_leaf_143_clk),
    .Q(\core.keymem.key_mem[10][54] ),
    .QN(_21562_));
 DFFR_X1 \core.keymem.key_mem[10][55]$_DFFE_PN0P_  (.D(_01043_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[10][55] ),
    .QN(_21561_));
 DFFR_X1 \core.keymem.key_mem[10][56]$_DFFE_PN0P_  (.D(_01044_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[10][56] ),
    .QN(_21560_));
 DFFR_X1 \core.keymem.key_mem[10][57]$_DFFE_PN0P_  (.D(_01045_),
    .RN(net100),
    .CK(clknet_leaf_108_clk),
    .Q(\core.keymem.key_mem[10][57] ),
    .QN(_21559_));
 DFFR_X1 \core.keymem.key_mem[10][58]$_DFFE_PN0P_  (.D(_01046_),
    .RN(net100),
    .CK(clknet_leaf_106_clk),
    .Q(\core.keymem.key_mem[10][58] ),
    .QN(_21558_));
 DFFR_X1 \core.keymem.key_mem[10][59]$_DFFE_PN0P_  (.D(_01047_),
    .RN(net100),
    .CK(clknet_leaf_18_clk),
    .Q(\core.keymem.key_mem[10][59] ),
    .QN(_21557_));
 DFFR_X1 \core.keymem.key_mem[10][5]$_DFFE_PN0P_  (.D(_01048_),
    .RN(net100),
    .CK(clknet_leaf_19_clk),
    .Q(\core.keymem.key_mem[10][5] ),
    .QN(_21556_));
 DFFR_X1 \core.keymem.key_mem[10][60]$_DFFE_PN0P_  (.D(_01049_),
    .RN(net82),
    .CK(clknet_leaf_24_clk),
    .Q(\core.keymem.key_mem[10][60] ),
    .QN(_21555_));
 DFFR_X1 \core.keymem.key_mem[10][61]$_DFFE_PN0P_  (.D(_01050_),
    .RN(net89),
    .CK(clknet_leaf_94_clk),
    .Q(\core.keymem.key_mem[10][61] ),
    .QN(_21554_));
 DFFR_X1 \core.keymem.key_mem[10][62]$_DFFE_PN0P_  (.D(_01051_),
    .RN(net100),
    .CK(clknet_leaf_99_clk),
    .Q(\core.keymem.key_mem[10][62] ),
    .QN(_21553_));
 DFFR_X1 \core.keymem.key_mem[10][63]$_DFFE_PN0P_  (.D(_01052_),
    .RN(net100),
    .CK(clknet_leaf_20_clk),
    .Q(\core.keymem.key_mem[10][63] ),
    .QN(_21552_));
 DFFR_X1 \core.keymem.key_mem[10][64]$_DFFE_PN0P_  (.D(_01053_),
    .RN(net100),
    .CK(clknet_leaf_15_clk),
    .Q(\core.keymem.key_mem[10][64] ),
    .QN(_21551_));
 DFFR_X1 \core.keymem.key_mem[10][65]$_DFFE_PN0P_  (.D(_01054_),
    .RN(net98),
    .CK(clknet_leaf_140_clk),
    .Q(\core.keymem.key_mem[10][65] ),
    .QN(_21550_));
 DFFR_X1 \core.keymem.key_mem[10][66]$_DFFE_PN0P_  (.D(_01055_),
    .RN(net100),
    .CK(clknet_leaf_15_clk),
    .Q(\core.keymem.key_mem[10][66] ),
    .QN(_21549_));
 DFFR_X1 \core.keymem.key_mem[10][67]$_DFFE_PN0P_  (.D(_01056_),
    .RN(net95),
    .CK(clknet_leaf_78_clk),
    .Q(\core.keymem.key_mem[10][67] ),
    .QN(_21548_));
 DFFR_X1 \core.keymem.key_mem[10][68]$_DFFE_PN0P_  (.D(_01057_),
    .RN(net95),
    .CK(clknet_leaf_76_clk),
    .Q(\core.keymem.key_mem[10][68] ),
    .QN(_21547_));
 DFFR_X1 \core.keymem.key_mem[10][69]$_DFFE_PN0P_  (.D(_01058_),
    .RN(net95),
    .CK(clknet_leaf_178_clk),
    .Q(\core.keymem.key_mem[10][69] ),
    .QN(_21546_));
 DFFR_X1 \core.keymem.key_mem[10][6]$_DFFE_PN0P_  (.D(_01059_),
    .RN(net100),
    .CK(clknet_leaf_103_clk),
    .Q(\core.keymem.key_mem[10][6] ),
    .QN(_21545_));
 DFFR_X1 \core.keymem.key_mem[10][70]$_DFFE_PN0P_  (.D(_01060_),
    .RN(net100),
    .CK(clknet_leaf_100_clk),
    .Q(\core.keymem.key_mem[10][70] ),
    .QN(_21544_));
 DFFR_X1 \core.keymem.key_mem[10][71]$_DFFE_PN0P_  (.D(_01061_),
    .RN(net99),
    .CK(clknet_leaf_74_clk),
    .Q(\core.keymem.key_mem[10][71] ),
    .QN(_21543_));
 DFFR_X1 \core.keymem.key_mem[10][72]$_DFFE_PN0P_  (.D(_01062_),
    .RN(net95),
    .CK(clknet_leaf_178_clk),
    .Q(\core.keymem.key_mem[10][72] ),
    .QN(_21542_));
 DFFR_X1 \core.keymem.key_mem[10][73]$_DFFE_PN0P_  (.D(_01063_),
    .RN(net97),
    .CK(clknet_leaf_147_clk),
    .Q(\core.keymem.key_mem[10][73] ),
    .QN(_21541_));
 DFFR_X1 \core.keymem.key_mem[10][74]$_DFFE_PN0P_  (.D(_01064_),
    .RN(net97),
    .CK(clknet_leaf_153_clk),
    .Q(\core.keymem.key_mem[10][74] ),
    .QN(_21540_));
 DFFR_X1 \core.keymem.key_mem[10][75]$_DFFE_PN0P_  (.D(_01065_),
    .RN(net97),
    .CK(clknet_leaf_154_clk),
    .Q(\core.keymem.key_mem[10][75] ),
    .QN(_21539_));
 DFFR_X1 \core.keymem.key_mem[10][76]$_DFFE_PN0P_  (.D(_01066_),
    .RN(net93),
    .CK(clknet_leaf_283_clk),
    .Q(\core.keymem.key_mem[10][76] ),
    .QN(_21538_));
 DFFR_X1 \core.keymem.key_mem[10][77]$_DFFE_PN0P_  (.D(_01067_),
    .RN(net97),
    .CK(clknet_leaf_160_clk),
    .Q(\core.keymem.key_mem[10][77] ),
    .QN(_21537_));
 DFFR_X1 \core.keymem.key_mem[10][78]$_DFFE_PN0P_  (.D(_01068_),
    .RN(net98),
    .CK(clknet_leaf_174_clk),
    .Q(\core.keymem.key_mem[10][78] ),
    .QN(_21536_));
 DFFR_X1 \core.keymem.key_mem[10][79]$_DFFE_PN0P_  (.D(_01069_),
    .RN(net96),
    .CK(clknet_leaf_229_clk),
    .Q(\core.keymem.key_mem[10][79] ),
    .QN(_21535_));
 DFFR_X1 \core.keymem.key_mem[10][7]$_DFFE_PN0P_  (.D(_01070_),
    .RN(net98),
    .CK(clknet_leaf_172_clk),
    .Q(\core.keymem.key_mem[10][7] ),
    .QN(_21534_));
 DFFR_X1 \core.keymem.key_mem[10][80]$_DFFE_PN0P_  (.D(_01071_),
    .RN(net97),
    .CK(clknet_leaf_158_clk),
    .Q(\core.keymem.key_mem[10][80] ),
    .QN(_21533_));
 DFFR_X1 \core.keymem.key_mem[10][81]$_DFFE_PN0P_  (.D(_01072_),
    .RN(net97),
    .CK(clknet_leaf_155_clk),
    .Q(\core.keymem.key_mem[10][81] ),
    .QN(_21532_));
 DFFR_X1 \core.keymem.key_mem[10][82]$_DFFE_PN0P_  (.D(_01073_),
    .RN(net98),
    .CK(clknet_leaf_180_clk),
    .Q(\core.keymem.key_mem[10][82] ),
    .QN(_21531_));
 DFFR_X1 \core.keymem.key_mem[10][83]$_DFFE_PN0P_  (.D(_01074_),
    .RN(net94),
    .CK(clknet_leaf_186_clk),
    .Q(\core.keymem.key_mem[10][83] ),
    .QN(_21530_));
 DFFR_X1 \core.keymem.key_mem[10][84]$_DFFE_PN0P_  (.D(_01075_),
    .RN(net95),
    .CK(clknet_leaf_179_clk),
    .Q(\core.keymem.key_mem[10][84] ),
    .QN(_21529_));
 DFFR_X1 \core.keymem.key_mem[10][85]$_DFFE_PN0P_  (.D(_01076_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[10][85] ),
    .QN(_21528_));
 DFFR_X1 \core.keymem.key_mem[10][86]$_DFFE_PN0P_  (.D(_01077_),
    .RN(net94),
    .CK(clknet_leaf_189_clk),
    .Q(\core.keymem.key_mem[10][86] ),
    .QN(_21527_));
 DFFR_X1 \core.keymem.key_mem[10][87]$_DFFE_PN0P_  (.D(_01078_),
    .RN(net93),
    .CK(clknet_leaf_57_clk),
    .Q(\core.keymem.key_mem[10][87] ),
    .QN(_21526_));
 DFFR_X1 \core.keymem.key_mem[10][88]$_DFFE_PN0P_  (.D(_01079_),
    .RN(net91),
    .CK(clknet_leaf_279_clk),
    .Q(\core.keymem.key_mem[10][88] ),
    .QN(_21525_));
 DFFR_X1 \core.keymem.key_mem[10][89]$_DFFE_PN0P_  (.D(_01080_),
    .RN(net93),
    .CK(clknet_leaf_281_clk),
    .Q(\core.keymem.key_mem[10][89] ),
    .QN(_21524_));
 DFFR_X1 \core.keymem.key_mem[10][8]$_DFFE_PN0P_  (.D(_01081_),
    .RN(net93),
    .CK(clknet_leaf_377_clk),
    .Q(\core.keymem.key_mem[10][8] ),
    .QN(_21523_));
 DFFR_X1 \core.keymem.key_mem[10][90]$_DFFE_PN0P_  (.D(_01082_),
    .RN(net97),
    .CK(clknet_leaf_161_clk),
    .Q(\core.keymem.key_mem[10][90] ),
    .QN(_21522_));
 DFFR_X1 \core.keymem.key_mem[10][91]$_DFFE_PN0P_  (.D(_01083_),
    .RN(net93),
    .CK(clknet_leaf_184_clk),
    .Q(\core.keymem.key_mem[10][91] ),
    .QN(_21521_));
 DFFR_X1 \core.keymem.key_mem[10][92]$_DFFE_PN0P_  (.D(_01084_),
    .RN(net95),
    .CK(clknet_leaf_63_clk),
    .Q(\core.keymem.key_mem[10][92] ),
    .QN(_21520_));
 DFFR_X1 \core.keymem.key_mem[10][93]$_DFFE_PN0P_  (.D(_01085_),
    .RN(net96),
    .CK(clknet_leaf_231_clk),
    .Q(\core.keymem.key_mem[10][93] ),
    .QN(_21519_));
 DFFR_X1 \core.keymem.key_mem[10][94]$_DFFE_PN0P_  (.D(_01086_),
    .RN(net94),
    .CK(clknet_leaf_214_clk),
    .Q(\core.keymem.key_mem[10][94] ),
    .QN(_21518_));
 DFFR_X1 \core.keymem.key_mem[10][95]$_DFFE_PN0P_  (.D(_01087_),
    .RN(net96),
    .CK(clknet_leaf_242_clk),
    .Q(\core.keymem.key_mem[10][95] ),
    .QN(_21517_));
 DFFR_X1 \core.keymem.key_mem[10][96]$_DFFE_PN0P_  (.D(_01088_),
    .RN(net92),
    .CK(clknet_leaf_266_clk),
    .Q(\core.keymem.key_mem[10][96] ),
    .QN(_21516_));
 DFFR_X1 \core.keymem.key_mem[10][97]$_DFFE_PN0P_  (.D(_01089_),
    .RN(net95),
    .CK(clknet_leaf_183_clk),
    .Q(\core.keymem.key_mem[10][97] ),
    .QN(_21515_));
 DFFR_X1 \core.keymem.key_mem[10][98]$_DFFE_PN0P_  (.D(_01090_),
    .RN(net93),
    .CK(clknet_leaf_195_clk),
    .Q(\core.keymem.key_mem[10][98] ),
    .QN(_21514_));
 DFFR_X1 \core.keymem.key_mem[10][99]$_DFFE_PN0P_  (.D(_01091_),
    .RN(net91),
    .CK(clknet_leaf_200_clk),
    .Q(\core.keymem.key_mem[10][99] ),
    .QN(_21513_));
 DFFR_X1 \core.keymem.key_mem[10][9]$_DFFE_PN0P_  (.D(_01092_),
    .RN(net91),
    .CK(clknet_leaf_203_clk),
    .Q(\core.keymem.key_mem[10][9] ),
    .QN(_21512_));
 DFFR_X1 \core.keymem.key_mem[11][0]$_DFFE_PN0P_  (.D(_01093_),
    .RN(net96),
    .CK(clknet_leaf_244_clk),
    .Q(\core.keymem.key_mem[11][0] ),
    .QN(_21511_));
 DFFR_X1 \core.keymem.key_mem[11][100]$_DFFE_PN0P_  (.D(_01094_),
    .RN(net98),
    .CK(clknet_leaf_212_clk),
    .Q(\core.keymem.key_mem[11][100] ),
    .QN(_21510_));
 DFFR_X1 \core.keymem.key_mem[11][101]$_DFFE_PN0P_  (.D(_01095_),
    .RN(net94),
    .CK(clknet_leaf_218_clk),
    .Q(\core.keymem.key_mem[11][101] ),
    .QN(_21509_));
 DFFR_X1 \core.keymem.key_mem[11][102]$_DFFE_PN0P_  (.D(_01096_),
    .RN(net96),
    .CK(clknet_leaf_234_clk),
    .Q(\core.keymem.key_mem[11][102] ),
    .QN(_21508_));
 DFFR_X1 \core.keymem.key_mem[11][103]$_DFFE_PN0P_  (.D(_01097_),
    .RN(net96),
    .CK(clknet_leaf_245_clk),
    .Q(\core.keymem.key_mem[11][103] ),
    .QN(_21507_));
 DFFR_X1 \core.keymem.key_mem[11][104]$_DFFE_PN0P_  (.D(_01098_),
    .RN(net93),
    .CK(clknet_leaf_192_clk),
    .Q(\core.keymem.key_mem[11][104] ),
    .QN(_21506_));
 DFFR_X1 \core.keymem.key_mem[11][105]$_DFFE_PN0P_  (.D(_01099_),
    .RN(net96),
    .CK(clknet_leaf_248_clk),
    .Q(\core.keymem.key_mem[11][105] ),
    .QN(_21505_));
 DFFR_X1 \core.keymem.key_mem[11][106]$_DFFE_PN0P_  (.D(_01100_),
    .RN(net92),
    .CK(clknet_leaf_269_clk),
    .Q(\core.keymem.key_mem[11][106] ),
    .QN(_21504_));
 DFFR_X1 \core.keymem.key_mem[11][107]$_DFFE_PN0P_  (.D(_01101_),
    .RN(net92),
    .CK(clknet_leaf_270_clk),
    .Q(\core.keymem.key_mem[11][107] ),
    .QN(_21503_));
 DFFR_X1 \core.keymem.key_mem[11][108]$_DFFE_PN0P_  (.D(_01102_),
    .RN(net92),
    .CK(clknet_leaf_277_clk),
    .Q(\core.keymem.key_mem[11][108] ),
    .QN(_21502_));
 DFFR_X1 \core.keymem.key_mem[11][109]$_DFFE_PN0P_  (.D(_01103_),
    .RN(net94),
    .CK(clknet_leaf_260_clk),
    .Q(\core.keymem.key_mem[11][109] ),
    .QN(_21501_));
 DFFR_X1 \core.keymem.key_mem[11][10]$_DFFE_PN0P_  (.D(_01104_),
    .RN(net95),
    .CK(clknet_leaf_187_clk),
    .Q(\core.keymem.key_mem[11][10] ),
    .QN(_21500_));
 DFFR_X1 \core.keymem.key_mem[11][110]$_DFFE_PN0P_  (.D(_01105_),
    .RN(net96),
    .CK(clknet_leaf_250_clk),
    .Q(\core.keymem.key_mem[11][110] ),
    .QN(_21499_));
 DFFR_X1 \core.keymem.key_mem[11][111]$_DFFE_PN0P_  (.D(_01106_),
    .RN(net96),
    .CK(clknet_leaf_224_clk),
    .Q(\core.keymem.key_mem[11][111] ),
    .QN(_21498_));
 DFFR_X1 \core.keymem.key_mem[11][112]$_DFFE_PN0P_  (.D(_01107_),
    .RN(net94),
    .CK(clknet_leaf_260_clk),
    .Q(\core.keymem.key_mem[11][112] ),
    .QN(_21497_));
 DFFR_X1 \core.keymem.key_mem[11][113]$_DFFE_PN0P_  (.D(_01108_),
    .RN(net92),
    .CK(clknet_leaf_273_clk),
    .Q(\core.keymem.key_mem[11][113] ),
    .QN(_21496_));
 DFFR_X1 \core.keymem.key_mem[11][114]$_DFFE_PN0P_  (.D(_01109_),
    .RN(net91),
    .CK(clknet_leaf_279_clk),
    .Q(\core.keymem.key_mem[11][114] ),
    .QN(_21495_));
 DFFR_X1 \core.keymem.key_mem[11][115]$_DFFE_PN0P_  (.D(_01110_),
    .RN(net92),
    .CK(clknet_leaf_276_clk),
    .Q(\core.keymem.key_mem[11][115] ),
    .QN(_21494_));
 DFFR_X1 \core.keymem.key_mem[11][116]$_DFFE_PN0P_  (.D(_01111_),
    .RN(net94),
    .CK(clknet_leaf_263_clk),
    .Q(\core.keymem.key_mem[11][116] ),
    .QN(_21493_));
 DFFR_X1 \core.keymem.key_mem[11][117]$_DFFE_PN0P_  (.D(_01112_),
    .RN(net96),
    .CK(clknet_leaf_222_clk),
    .Q(\core.keymem.key_mem[11][117] ),
    .QN(_21492_));
 DFFR_X1 \core.keymem.key_mem[11][118]$_DFFE_PN0P_  (.D(_01113_),
    .RN(net97),
    .CK(clknet_leaf_241_clk),
    .Q(\core.keymem.key_mem[11][118] ),
    .QN(_21491_));
 DFFR_X1 \core.keymem.key_mem[11][119]$_DFFE_PN0P_  (.D(_01114_),
    .RN(net94),
    .CK(clknet_leaf_262_clk),
    .Q(\core.keymem.key_mem[11][119] ),
    .QN(_21490_));
 DFFR_X1 \core.keymem.key_mem[11][11]$_DFFE_PN0P_  (.D(_01115_),
    .RN(net95),
    .CK(clknet_leaf_60_clk),
    .Q(\core.keymem.key_mem[11][11] ),
    .QN(_21489_));
 DFFR_X1 \core.keymem.key_mem[11][120]$_DFFE_PN0P_  (.D(_01116_),
    .RN(net94),
    .CK(clknet_leaf_216_clk),
    .Q(\core.keymem.key_mem[11][120] ),
    .QN(_21488_));
 DFFR_X1 \core.keymem.key_mem[11][121]$_DFFE_PN0P_  (.D(_01117_),
    .RN(net94),
    .CK(clknet_leaf_264_clk),
    .Q(\core.keymem.key_mem[11][121] ),
    .QN(_21487_));
 DFFR_X1 \core.keymem.key_mem[11][122]$_DFFE_PN0P_  (.D(_01118_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[11][122] ),
    .QN(_21486_));
 DFFR_X1 \core.keymem.key_mem[11][123]$_DFFE_PN0P_  (.D(_01119_),
    .RN(net93),
    .CK(clknet_leaf_196_clk),
    .Q(\core.keymem.key_mem[11][123] ),
    .QN(_21485_));
 DFFR_X1 \core.keymem.key_mem[11][124]$_DFFE_PN0P_  (.D(_01120_),
    .RN(net93),
    .CK(clknet_leaf_57_clk),
    .Q(\core.keymem.key_mem[11][124] ),
    .QN(_21484_));
 DFFR_X1 \core.keymem.key_mem[11][125]$_DFFE_PN0P_  (.D(_01121_),
    .RN(net97),
    .CK(clknet_leaf_236_clk),
    .Q(\core.keymem.key_mem[11][125] ),
    .QN(_21483_));
 DFFR_X1 \core.keymem.key_mem[11][126]$_DFFE_PN0P_  (.D(_01122_),
    .RN(net98),
    .CK(clknet_leaf_167_clk),
    .Q(\core.keymem.key_mem[11][126] ),
    .QN(_21482_));
 DFFR_X1 \core.keymem.key_mem[11][127]$_DFFE_PN0P_  (.D(_01123_),
    .RN(net97),
    .CK(clknet_leaf_243_clk),
    .Q(\core.keymem.key_mem[11][127] ),
    .QN(_21481_));
 DFFR_X1 \core.keymem.key_mem[11][12]$_DFFE_PN0P_  (.D(_01124_),
    .RN(net93),
    .CK(clknet_leaf_205_clk),
    .Q(\core.keymem.key_mem[11][12] ),
    .QN(_21480_));
 DFFR_X1 \core.keymem.key_mem[11][13]$_DFFE_PN0P_  (.D(_01125_),
    .RN(net87),
    .CK(clknet_leaf_31_clk),
    .Q(\core.keymem.key_mem[11][13] ),
    .QN(_21479_));
 DFFR_X1 \core.keymem.key_mem[11][14]$_DFFE_PN0P_  (.D(_01126_),
    .RN(net94),
    .CK(clknet_leaf_209_clk),
    .Q(\core.keymem.key_mem[11][14] ),
    .QN(_21478_));
 DFFR_X1 \core.keymem.key_mem[11][15]$_DFFE_PN0P_  (.D(_01127_),
    .RN(net96),
    .CK(clknet_leaf_165_clk),
    .Q(\core.keymem.key_mem[11][15] ),
    .QN(_21477_));
 DFFR_X1 \core.keymem.key_mem[11][16]$_DFFE_PN0P_  (.D(_01128_),
    .RN(net87),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[11][16] ),
    .QN(_21476_));
 DFFR_X1 \core.keymem.key_mem[11][17]$_DFFE_PN0P_  (.D(_01129_),
    .RN(net98),
    .CK(clknet_leaf_168_clk),
    .Q(\core.keymem.key_mem[11][17] ),
    .QN(_21475_));
 DFFR_X1 \core.keymem.key_mem[11][18]$_DFFE_PN0P_  (.D(_01130_),
    .RN(net89),
    .CK(clknet_leaf_34_clk),
    .Q(\core.keymem.key_mem[11][18] ),
    .QN(_21474_));
 DFFR_X1 \core.keymem.key_mem[11][19]$_DFFE_PN0P_  (.D(_01131_),
    .RN(net85),
    .CK(clknet_leaf_49_clk),
    .Q(\core.keymem.key_mem[11][19] ),
    .QN(_21473_));
 DFFR_X1 \core.keymem.key_mem[11][1]$_DFFE_PN0P_  (.D(_01132_),
    .RN(net89),
    .CK(clknet_leaf_22_clk),
    .Q(\core.keymem.key_mem[11][1] ),
    .QN(_21472_));
 DFFR_X1 \core.keymem.key_mem[11][20]$_DFFE_PN0P_  (.D(_01133_),
    .RN(net100),
    .CK(clknet_leaf_22_clk),
    .Q(\core.keymem.key_mem[11][20] ),
    .QN(_21471_));
 DFFR_X1 \core.keymem.key_mem[11][21]$_DFFE_PN0P_  (.D(_01134_),
    .RN(net85),
    .CK(clknet_leaf_67_clk),
    .Q(\core.keymem.key_mem[11][21] ),
    .QN(_21470_));
 DFFR_X1 \core.keymem.key_mem[11][22]$_DFFE_PN0P_  (.D(_01135_),
    .RN(net94),
    .CK(clknet_leaf_219_clk),
    .Q(\core.keymem.key_mem[11][22] ),
    .QN(_21469_));
 DFFR_X1 \core.keymem.key_mem[11][23]$_DFFE_PN0P_  (.D(_01136_),
    .RN(net89),
    .CK(clknet_leaf_379_clk),
    .Q(\core.keymem.key_mem[11][23] ),
    .QN(_21468_));
 DFFR_X1 \core.keymem.key_mem[11][24]$_DFFE_PN0P_  (.D(_01137_),
    .RN(net85),
    .CK(clknet_leaf_49_clk),
    .Q(\core.keymem.key_mem[11][24] ),
    .QN(_21467_));
 DFFR_X1 \core.keymem.key_mem[11][25]$_DFFE_PN0P_  (.D(_01138_),
    .RN(net85),
    .CK(clknet_leaf_48_clk),
    .Q(\core.keymem.key_mem[11][25] ),
    .QN(_21466_));
 DFFR_X1 \core.keymem.key_mem[11][26]$_DFFE_PN0P_  (.D(_01139_),
    .RN(net100),
    .CK(clknet_leaf_97_clk),
    .Q(\core.keymem.key_mem[11][26] ),
    .QN(_21465_));
 DFFR_X1 \core.keymem.key_mem[11][27]$_DFFE_PN0P_  (.D(_01140_),
    .RN(net16),
    .CK(clknet_leaf_151_clk),
    .Q(\core.keymem.key_mem[11][27] ),
    .QN(_21464_));
 DFFR_X1 \core.keymem.key_mem[11][28]$_DFFE_PN0P_  (.D(_01141_),
    .RN(net16),
    .CK(clknet_leaf_131_clk),
    .Q(\core.keymem.key_mem[11][28] ),
    .QN(_21463_));
 DFFR_X1 \core.keymem.key_mem[11][29]$_DFFE_PN0P_  (.D(_01142_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[11][29] ),
    .QN(_21462_));
 DFFR_X1 \core.keymem.key_mem[11][2]$_DFFE_PN0P_  (.D(_01143_),
    .RN(net89),
    .CK(clknet_leaf_63_clk),
    .Q(\core.keymem.key_mem[11][2] ),
    .QN(_21461_));
 DFFR_X1 \core.keymem.key_mem[11][30]$_DFFE_PN0P_  (.D(_01144_),
    .RN(net16),
    .CK(clknet_leaf_139_clk),
    .Q(\core.keymem.key_mem[11][30] ),
    .QN(_21460_));
 DFFR_X1 \core.keymem.key_mem[11][31]$_DFFE_PN0P_  (.D(_01145_),
    .RN(net16),
    .CK(clknet_leaf_138_clk),
    .Q(\core.keymem.key_mem[11][31] ),
    .QN(_21459_));
 DFFR_X1 \core.keymem.key_mem[11][32]$_DFFE_PN0P_  (.D(_01146_),
    .RN(net100),
    .CK(clknet_leaf_111_clk),
    .Q(\core.keymem.key_mem[11][32] ),
    .QN(_21458_));
 DFFR_X1 \core.keymem.key_mem[11][33]$_DFFE_PN0P_  (.D(_01147_),
    .RN(net99),
    .CK(clknet_leaf_127_clk),
    .Q(\core.keymem.key_mem[11][33] ),
    .QN(_21457_));
 DFFR_X1 \core.keymem.key_mem[11][34]$_DFFE_PN0P_  (.D(_01148_),
    .RN(net16),
    .CK(clknet_leaf_125_clk),
    .Q(\core.keymem.key_mem[11][34] ),
    .QN(_21456_));
 DFFR_X1 \core.keymem.key_mem[11][35]$_DFFE_PN0P_  (.D(_01149_),
    .RN(net99),
    .CK(clknet_leaf_122_clk),
    .Q(\core.keymem.key_mem[11][35] ),
    .QN(_21455_));
 DFFR_X1 \core.keymem.key_mem[11][36]$_DFFE_PN0P_  (.D(_01150_),
    .RN(net87),
    .CK(clknet_leaf_28_clk),
    .Q(\core.keymem.key_mem[11][36] ),
    .QN(_21454_));
 DFFR_X1 \core.keymem.key_mem[11][37]$_DFFE_PN0P_  (.D(_01151_),
    .RN(net88),
    .CK(clknet_leaf_90_clk),
    .Q(\core.keymem.key_mem[11][37] ),
    .QN(_21453_));
 DFFR_X1 \core.keymem.key_mem[11][38]$_DFFE_PN0P_  (.D(_01152_),
    .RN(net99),
    .CK(clknet_leaf_127_clk),
    .Q(\core.keymem.key_mem[11][38] ),
    .QN(_21452_));
 DFFR_X1 \core.keymem.key_mem[11][39]$_DFFE_PN0P_  (.D(_01153_),
    .RN(net85),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[11][39] ),
    .QN(_21451_));
 DFFR_X1 \core.keymem.key_mem[11][3]$_DFFE_PN0P_  (.D(_01154_),
    .RN(net85),
    .CK(clknet_leaf_46_clk),
    .Q(\core.keymem.key_mem[11][3] ),
    .QN(_21450_));
 DFFR_X1 \core.keymem.key_mem[11][40]$_DFFE_PN0P_  (.D(_01155_),
    .RN(net88),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[11][40] ),
    .QN(_21449_));
 DFFR_X1 \core.keymem.key_mem[11][41]$_DFFE_PN0P_  (.D(_01156_),
    .RN(net100),
    .CK(clknet_leaf_114_clk),
    .Q(\core.keymem.key_mem[11][41] ),
    .QN(_21448_));
 DFFR_X1 \core.keymem.key_mem[11][42]$_DFFE_PN0P_  (.D(_01157_),
    .RN(net100),
    .CK(clknet_leaf_128_clk),
    .Q(\core.keymem.key_mem[11][42] ),
    .QN(_21447_));
 DFFR_X1 \core.keymem.key_mem[11][43]$_DFFE_PN0P_  (.D(_01158_),
    .RN(net85),
    .CK(clknet_leaf_88_clk),
    .Q(\core.keymem.key_mem[11][43] ),
    .QN(_21446_));
 DFFR_X1 \core.keymem.key_mem[11][44]$_DFFE_PN0P_  (.D(_01159_),
    .RN(net100),
    .CK(clknet_leaf_113_clk),
    .Q(\core.keymem.key_mem[11][44] ),
    .QN(_21445_));
 DFFR_X1 \core.keymem.key_mem[11][45]$_DFFE_PN0P_  (.D(_01160_),
    .RN(net89),
    .CK(clknet_leaf_70_clk),
    .Q(\core.keymem.key_mem[11][45] ),
    .QN(_21444_));
 DFFR_X1 \core.keymem.key_mem[11][46]$_DFFE_PN0P_  (.D(_01161_),
    .RN(net99),
    .CK(clknet_leaf_82_clk),
    .Q(\core.keymem.key_mem[11][46] ),
    .QN(_21443_));
 DFFR_X1 \core.keymem.key_mem[11][47]$_DFFE_PN0P_  (.D(_01162_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[11][47] ),
    .QN(_21442_));
 DFFR_X1 \core.keymem.key_mem[11][48]$_DFFE_PN0P_  (.D(_01163_),
    .RN(net95),
    .CK(clknet_leaf_121_clk),
    .Q(\core.keymem.key_mem[11][48] ),
    .QN(_21441_));
 DFFR_X1 \core.keymem.key_mem[11][49]$_DFFE_PN0P_  (.D(_01164_),
    .RN(net99),
    .CK(clknet_leaf_81_clk),
    .Q(\core.keymem.key_mem[11][49] ),
    .QN(_21440_));
 DFFR_X1 \core.keymem.key_mem[11][4]$_DFFE_PN0P_  (.D(_01165_),
    .RN(net100),
    .CK(clknet_leaf_104_clk),
    .Q(\core.keymem.key_mem[11][4] ),
    .QN(_21439_));
 DFFR_X1 \core.keymem.key_mem[11][50]$_DFFE_PN0P_  (.D(_01166_),
    .RN(net98),
    .CK(clknet_leaf_140_clk),
    .Q(\core.keymem.key_mem[11][50] ),
    .QN(_21438_));
 DFFR_X1 \core.keymem.key_mem[11][51]$_DFFE_PN0P_  (.D(_01167_),
    .RN(net100),
    .CK(clknet_leaf_130_clk),
    .Q(\core.keymem.key_mem[11][51] ),
    .QN(_21437_));
 DFFR_X1 \core.keymem.key_mem[11][52]$_DFFE_PN0P_  (.D(_01168_),
    .RN(net99),
    .CK(clknet_leaf_80_clk),
    .Q(\core.keymem.key_mem[11][52] ),
    .QN(_21436_));
 DFFR_X1 \core.keymem.key_mem[11][53]$_DFFE_PN0P_  (.D(_01169_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[11][53] ),
    .QN(_21435_));
 DFFR_X1 \core.keymem.key_mem[11][54]$_DFFE_PN0P_  (.D(_01170_),
    .RN(net98),
    .CK(clknet_leaf_142_clk),
    .Q(\core.keymem.key_mem[11][54] ),
    .QN(_21434_));
 DFFR_X1 \core.keymem.key_mem[11][55]$_DFFE_PN0P_  (.D(_01171_),
    .RN(net16),
    .CK(clknet_leaf_138_clk),
    .Q(\core.keymem.key_mem[11][55] ),
    .QN(_21433_));
 DFFR_X1 \core.keymem.key_mem[11][56]$_DFFE_PN0P_  (.D(_01172_),
    .RN(net16),
    .CK(clknet_leaf_138_clk),
    .Q(\core.keymem.key_mem[11][56] ),
    .QN(_21432_));
 DFFR_X1 \core.keymem.key_mem[11][57]$_DFFE_PN0P_  (.D(_01173_),
    .RN(net100),
    .CK(clknet_leaf_109_clk),
    .Q(\core.keymem.key_mem[11][57] ),
    .QN(_21431_));
 DFFR_X1 \core.keymem.key_mem[11][58]$_DFFE_PN0P_  (.D(_01174_),
    .RN(net100),
    .CK(clknet_leaf_107_clk),
    .Q(\core.keymem.key_mem[11][58] ),
    .QN(_21430_));
 DFFR_X1 \core.keymem.key_mem[11][59]$_DFFE_PN0P_  (.D(_01175_),
    .RN(net100),
    .CK(clknet_leaf_17_clk),
    .Q(\core.keymem.key_mem[11][59] ),
    .QN(_21429_));
 DFFR_X1 \core.keymem.key_mem[11][5]$_DFFE_PN0P_  (.D(_01176_),
    .RN(net100),
    .CK(clknet_leaf_19_clk),
    .Q(\core.keymem.key_mem[11][5] ),
    .QN(_21428_));
 DFFR_X1 \core.keymem.key_mem[11][60]$_DFFE_PN0P_  (.D(_01177_),
    .RN(net82),
    .CK(clknet_leaf_24_clk),
    .Q(\core.keymem.key_mem[11][60] ),
    .QN(_21427_));
 DFFR_X1 \core.keymem.key_mem[11][61]$_DFFE_PN0P_  (.D(_01178_),
    .RN(net88),
    .CK(clknet_leaf_94_clk),
    .Q(\core.keymem.key_mem[11][61] ),
    .QN(_21426_));
 DFFR_X1 \core.keymem.key_mem[11][62]$_DFFE_PN0P_  (.D(_01179_),
    .RN(net100),
    .CK(clknet_leaf_98_clk),
    .Q(\core.keymem.key_mem[11][62] ),
    .QN(_21425_));
 DFFR_X1 \core.keymem.key_mem[11][63]$_DFFE_PN0P_  (.D(_01180_),
    .RN(net100),
    .CK(clknet_leaf_20_clk),
    .Q(\core.keymem.key_mem[11][63] ),
    .QN(_21424_));
 DFFR_X1 \core.keymem.key_mem[11][64]$_DFFE_PN0P_  (.D(_01181_),
    .RN(net100),
    .CK(clknet_leaf_15_clk),
    .Q(\core.keymem.key_mem[11][64] ),
    .QN(_21423_));
 DFFR_X1 \core.keymem.key_mem[11][65]$_DFFE_PN0P_  (.D(_01182_),
    .RN(net98),
    .CK(clknet_leaf_140_clk),
    .Q(\core.keymem.key_mem[11][65] ),
    .QN(_21422_));
 DFFR_X1 \core.keymem.key_mem[11][66]$_DFFE_PN0P_  (.D(_01183_),
    .RN(net100),
    .CK(clknet_leaf_17_clk),
    .Q(\core.keymem.key_mem[11][66] ),
    .QN(_21421_));
 DFFR_X1 \core.keymem.key_mem[11][67]$_DFFE_PN0P_  (.D(_01184_),
    .RN(net95),
    .CK(clknet_leaf_75_clk),
    .Q(\core.keymem.key_mem[11][67] ),
    .QN(_21420_));
 DFFR_X1 \core.keymem.key_mem[11][68]$_DFFE_PN0P_  (.D(_01185_),
    .RN(net95),
    .CK(clknet_leaf_118_clk),
    .Q(\core.keymem.key_mem[11][68] ),
    .QN(_21419_));
 DFFR_X1 \core.keymem.key_mem[11][69]$_DFFE_PN0P_  (.D(_01186_),
    .RN(net98),
    .CK(clknet_leaf_177_clk),
    .Q(\core.keymem.key_mem[11][69] ),
    .QN(_21418_));
 DFFR_X1 \core.keymem.key_mem[11][6]$_DFFE_PN0P_  (.D(_01187_),
    .RN(net100),
    .CK(clknet_leaf_101_clk),
    .Q(\core.keymem.key_mem[11][6] ),
    .QN(_21417_));
 DFFR_X1 \core.keymem.key_mem[11][70]$_DFFE_PN0P_  (.D(_01188_),
    .RN(net100),
    .CK(clknet_leaf_101_clk),
    .Q(\core.keymem.key_mem[11][70] ),
    .QN(_21416_));
 DFFR_X1 \core.keymem.key_mem[11][71]$_DFFE_PN0P_  (.D(_01189_),
    .RN(net99),
    .CK(clknet_leaf_73_clk),
    .Q(\core.keymem.key_mem[11][71] ),
    .QN(_21415_));
 DFFR_X1 \core.keymem.key_mem[11][72]$_DFFE_PN0P_  (.D(_01190_),
    .RN(net95),
    .CK(clknet_leaf_179_clk),
    .Q(\core.keymem.key_mem[11][72] ),
    .QN(_21414_));
 DFFR_X1 \core.keymem.key_mem[11][73]$_DFFE_PN0P_  (.D(_01191_),
    .RN(net97),
    .CK(clknet_leaf_152_clk),
    .Q(\core.keymem.key_mem[11][73] ),
    .QN(_21413_));
 DFFR_X1 \core.keymem.key_mem[11][74]$_DFFE_PN0P_  (.D(_01192_),
    .RN(net97),
    .CK(clknet_leaf_157_clk),
    .Q(\core.keymem.key_mem[11][74] ),
    .QN(_21412_));
 DFFR_X1 \core.keymem.key_mem[11][75]$_DFFE_PN0P_  (.D(_01193_),
    .RN(net97),
    .CK(clknet_leaf_152_clk),
    .Q(\core.keymem.key_mem[11][75] ),
    .QN(_21411_));
 DFFR_X1 \core.keymem.key_mem[11][76]$_DFFE_PN0P_  (.D(_01194_),
    .RN(net91),
    .CK(clknet_leaf_284_clk),
    .Q(\core.keymem.key_mem[11][76] ),
    .QN(_21410_));
 DFFR_X1 \core.keymem.key_mem[11][77]$_DFFE_PN0P_  (.D(_01195_),
    .RN(net97),
    .CK(clknet_leaf_160_clk),
    .Q(\core.keymem.key_mem[11][77] ),
    .QN(_21409_));
 DFFR_X1 \core.keymem.key_mem[11][78]$_DFFE_PN0P_  (.D(_01196_),
    .RN(net97),
    .CK(clknet_leaf_164_clk),
    .Q(\core.keymem.key_mem[11][78] ),
    .QN(_21408_));
 DFFR_X1 \core.keymem.key_mem[11][79]$_DFFE_PN0P_  (.D(_01197_),
    .RN(net98),
    .CK(clknet_leaf_228_clk),
    .Q(\core.keymem.key_mem[11][79] ),
    .QN(_21407_));
 DFFR_X1 \core.keymem.key_mem[11][7]$_DFFE_PN0P_  (.D(_01198_),
    .RN(net98),
    .CK(clknet_leaf_174_clk),
    .Q(\core.keymem.key_mem[11][7] ),
    .QN(_21406_));
 DFFR_X1 \core.keymem.key_mem[11][80]$_DFFE_PN0P_  (.D(_01199_),
    .RN(net97),
    .CK(clknet_leaf_157_clk),
    .Q(\core.keymem.key_mem[11][80] ),
    .QN(_21405_));
 DFFR_X1 \core.keymem.key_mem[11][81]$_DFFE_PN0P_  (.D(_01200_),
    .RN(net97),
    .CK(clknet_leaf_153_clk),
    .Q(\core.keymem.key_mem[11][81] ),
    .QN(_21404_));
 DFFR_X1 \core.keymem.key_mem[11][82]$_DFFE_PN0P_  (.D(_01201_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[11][82] ),
    .QN(_21403_));
 DFFR_X1 \core.keymem.key_mem[11][83]$_DFFE_PN0P_  (.D(_01202_),
    .RN(net95),
    .CK(clknet_leaf_185_clk),
    .Q(\core.keymem.key_mem[11][83] ),
    .QN(_21402_));
 DFFR_X1 \core.keymem.key_mem[11][84]$_DFFE_PN0P_  (.D(_01203_),
    .RN(net95),
    .CK(clknet_leaf_179_clk),
    .Q(\core.keymem.key_mem[11][84] ),
    .QN(_21401_));
 DFFR_X1 \core.keymem.key_mem[11][85]$_DFFE_PN0P_  (.D(_01204_),
    .RN(net97),
    .CK(clknet_leaf_237_clk),
    .Q(\core.keymem.key_mem[11][85] ),
    .QN(_21400_));
 DFFR_X1 \core.keymem.key_mem[11][86]$_DFFE_PN0P_  (.D(_01205_),
    .RN(net94),
    .CK(clknet_leaf_209_clk),
    .Q(\core.keymem.key_mem[11][86] ),
    .QN(_21399_));
 DFFR_X1 \core.keymem.key_mem[11][87]$_DFFE_PN0P_  (.D(_01206_),
    .RN(net93),
    .CK(clknet_leaf_57_clk),
    .Q(\core.keymem.key_mem[11][87] ),
    .QN(_21398_));
 DFFR_X1 \core.keymem.key_mem[11][88]$_DFFE_PN0P_  (.D(_01207_),
    .RN(net91),
    .CK(clknet_leaf_283_clk),
    .Q(\core.keymem.key_mem[11][88] ),
    .QN(_21397_));
 DFFR_X1 \core.keymem.key_mem[11][89]$_DFFE_PN0P_  (.D(_01208_),
    .RN(net93),
    .CK(clknet_leaf_199_clk),
    .Q(\core.keymem.key_mem[11][89] ),
    .QN(_21396_));
 DFFR_X1 \core.keymem.key_mem[11][8]$_DFFE_PN0P_  (.D(_01209_),
    .RN(net89),
    .CK(clknet_leaf_377_clk),
    .Q(\core.keymem.key_mem[11][8] ),
    .QN(_21395_));
 DFFR_X1 \core.keymem.key_mem[11][90]$_DFFE_PN0P_  (.D(_01210_),
    .RN(net97),
    .CK(clknet_leaf_156_clk),
    .Q(\core.keymem.key_mem[11][90] ),
    .QN(_21394_));
 DFFR_X1 \core.keymem.key_mem[11][91]$_DFFE_PN0P_  (.D(_01211_),
    .RN(net95),
    .CK(clknet_leaf_185_clk),
    .Q(\core.keymem.key_mem[11][91] ),
    .QN(_21393_));
 DFFR_X1 \core.keymem.key_mem[11][92]$_DFFE_PN0P_  (.D(_01212_),
    .RN(net95),
    .CK(clknet_leaf_72_clk),
    .Q(\core.keymem.key_mem[11][92] ),
    .QN(_21392_));
 DFFR_X1 \core.keymem.key_mem[11][93]$_DFFE_PN0P_  (.D(_01213_),
    .RN(net94),
    .CK(clknet_leaf_189_clk),
    .Q(\core.keymem.key_mem[11][93] ),
    .QN(_21391_));
 DFFR_X1 \core.keymem.key_mem[11][94]$_DFFE_PN0P_  (.D(_01214_),
    .RN(net94),
    .CK(clknet_leaf_218_clk),
    .Q(\core.keymem.key_mem[11][94] ),
    .QN(_21390_));
 DFFR_X1 \core.keymem.key_mem[11][95]$_DFFE_PN0P_  (.D(_01215_),
    .RN(net96),
    .CK(clknet_leaf_244_clk),
    .Q(\core.keymem.key_mem[11][95] ),
    .QN(_21389_));
 DFFR_X1 \core.keymem.key_mem[11][96]$_DFFE_PN0P_  (.D(_01216_),
    .RN(net92),
    .CK(clknet_leaf_204_clk),
    .Q(\core.keymem.key_mem[11][96] ),
    .QN(_21388_));
 DFFR_X1 \core.keymem.key_mem[11][97]$_DFFE_PN0P_  (.D(_01217_),
    .RN(net93),
    .CK(clknet_leaf_194_clk),
    .Q(\core.keymem.key_mem[11][97] ),
    .QN(_21387_));
 DFFR_X1 \core.keymem.key_mem[11][98]$_DFFE_PN0P_  (.D(_01218_),
    .RN(net95),
    .CK(clknet_leaf_194_clk),
    .Q(\core.keymem.key_mem[11][98] ),
    .QN(_21386_));
 DFFR_X1 \core.keymem.key_mem[11][99]$_DFFE_PN0P_  (.D(_01219_),
    .RN(net92),
    .CK(clknet_leaf_207_clk),
    .Q(\core.keymem.key_mem[11][99] ),
    .QN(_21385_));
 DFFR_X1 \core.keymem.key_mem[11][9]$_DFFE_PN0P_  (.D(_01220_),
    .RN(net92),
    .CK(clknet_leaf_205_clk),
    .Q(\core.keymem.key_mem[11][9] ),
    .QN(_21384_));
 DFFR_X1 \core.keymem.key_mem[12][0]$_DFFE_PN0P_  (.D(_01221_),
    .RN(net96),
    .CK(clknet_leaf_247_clk),
    .Q(\core.keymem.key_mem[12][0] ),
    .QN(_21383_));
 DFFR_X1 \core.keymem.key_mem[12][100]$_DFFE_PN0P_  (.D(_01222_),
    .RN(net94),
    .CK(clknet_leaf_211_clk),
    .Q(\core.keymem.key_mem[12][100] ),
    .QN(_21382_));
 DFFR_X1 \core.keymem.key_mem[12][101]$_DFFE_PN0P_  (.D(_01223_),
    .RN(net94),
    .CK(clknet_leaf_218_clk),
    .Q(\core.keymem.key_mem[12][101] ),
    .QN(_21381_));
 DFFR_X1 \core.keymem.key_mem[12][102]$_DFFE_PN0P_  (.D(_01224_),
    .RN(net96),
    .CK(clknet_leaf_232_clk),
    .Q(\core.keymem.key_mem[12][102] ),
    .QN(_21380_));
 DFFR_X1 \core.keymem.key_mem[12][103]$_DFFE_PN0P_  (.D(_01225_),
    .RN(net96),
    .CK(clknet_leaf_246_clk),
    .Q(\core.keymem.key_mem[12][103] ),
    .QN(_21379_));
 DFFR_X1 \core.keymem.key_mem[12][104]$_DFFE_PN0P_  (.D(_01226_),
    .RN(net93),
    .CK(clknet_leaf_192_clk),
    .Q(\core.keymem.key_mem[12][104] ),
    .QN(_21378_));
 DFFR_X1 \core.keymem.key_mem[12][105]$_DFFE_PN0P_  (.D(_01227_),
    .RN(net96),
    .CK(clknet_leaf_246_clk),
    .Q(\core.keymem.key_mem[12][105] ),
    .QN(_21377_));
 DFFR_X1 \core.keymem.key_mem[12][106]$_DFFE_PN0P_  (.D(_01228_),
    .RN(net92),
    .CK(clknet_leaf_269_clk),
    .Q(\core.keymem.key_mem[12][106] ),
    .QN(_21376_));
 DFFR_X1 \core.keymem.key_mem[12][107]$_DFFE_PN0P_  (.D(_01229_),
    .RN(net92),
    .CK(clknet_leaf_267_clk),
    .Q(\core.keymem.key_mem[12][107] ),
    .QN(_21375_));
 DFFR_X1 \core.keymem.key_mem[12][108]$_DFFE_PN0P_  (.D(_01230_),
    .RN(net92),
    .CK(clknet_leaf_277_clk),
    .Q(\core.keymem.key_mem[12][108] ),
    .QN(_21374_));
 DFFR_X1 \core.keymem.key_mem[12][109]$_DFFE_PN0P_  (.D(_01231_),
    .RN(net94),
    .CK(clknet_leaf_263_clk),
    .Q(\core.keymem.key_mem[12][109] ),
    .QN(_21373_));
 DFFR_X1 \core.keymem.key_mem[12][10]$_DFFE_PN0P_  (.D(_01232_),
    .RN(net98),
    .CK(clknet_leaf_167_clk),
    .Q(\core.keymem.key_mem[12][10] ),
    .QN(_21372_));
 DFFR_X1 \core.keymem.key_mem[12][110]$_DFFE_PN0P_  (.D(_01233_),
    .RN(net96),
    .CK(clknet_leaf_249_clk),
    .Q(\core.keymem.key_mem[12][110] ),
    .QN(_21371_));
 DFFR_X1 \core.keymem.key_mem[12][111]$_DFFE_PN0P_  (.D(_01234_),
    .RN(net96),
    .CK(clknet_leaf_224_clk),
    .Q(\core.keymem.key_mem[12][111] ),
    .QN(_21370_));
 DFFR_X1 \core.keymem.key_mem[12][112]$_DFFE_PN0P_  (.D(_01235_),
    .RN(net94),
    .CK(clknet_leaf_261_clk),
    .Q(\core.keymem.key_mem[12][112] ),
    .QN(_21369_));
 DFFR_X1 \core.keymem.key_mem[12][113]$_DFFE_PN0P_  (.D(_01236_),
    .RN(net91),
    .CK(clknet_leaf_274_clk),
    .Q(\core.keymem.key_mem[12][113] ),
    .QN(_21368_));
 DFFR_X1 \core.keymem.key_mem[12][114]$_DFFE_PN0P_  (.D(_01237_),
    .RN(net91),
    .CK(clknet_leaf_278_clk),
    .Q(\core.keymem.key_mem[12][114] ),
    .QN(_21367_));
 DFFR_X1 \core.keymem.key_mem[12][115]$_DFFE_PN0P_  (.D(_01238_),
    .RN(net92),
    .CK(clknet_leaf_275_clk),
    .Q(\core.keymem.key_mem[12][115] ),
    .QN(_21366_));
 DFFR_X1 \core.keymem.key_mem[12][116]$_DFFE_PN0P_  (.D(_01239_),
    .RN(net94),
    .CK(clknet_leaf_265_clk),
    .Q(\core.keymem.key_mem[12][116] ),
    .QN(_21365_));
 DFFR_X1 \core.keymem.key_mem[12][117]$_DFFE_PN0P_  (.D(_01240_),
    .RN(net96),
    .CK(clknet_leaf_223_clk),
    .Q(\core.keymem.key_mem[12][117] ),
    .QN(_21364_));
 DFFR_X1 \core.keymem.key_mem[12][118]$_DFFE_PN0P_  (.D(_01241_),
    .RN(net97),
    .CK(clknet_leaf_244_clk),
    .Q(\core.keymem.key_mem[12][118] ),
    .QN(_21363_));
 DFFR_X1 \core.keymem.key_mem[12][119]$_DFFE_PN0P_  (.D(_01242_),
    .RN(net94),
    .CK(clknet_leaf_220_clk),
    .Q(\core.keymem.key_mem[12][119] ),
    .QN(_21362_));
 DFFR_X1 \core.keymem.key_mem[12][11]$_DFFE_PN0P_  (.D(_01243_),
    .RN(net95),
    .CK(clknet_leaf_60_clk),
    .Q(\core.keymem.key_mem[12][11] ),
    .QN(_21361_));
 DFFR_X1 \core.keymem.key_mem[12][120]$_DFFE_PN0P_  (.D(_01244_),
    .RN(net94),
    .CK(clknet_leaf_215_clk),
    .Q(\core.keymem.key_mem[12][120] ),
    .QN(_21360_));
 DFFR_X1 \core.keymem.key_mem[12][121]$_DFFE_PN0P_  (.D(_01245_),
    .RN(net94),
    .CK(clknet_leaf_216_clk),
    .Q(\core.keymem.key_mem[12][121] ),
    .QN(_21359_));
 DFFR_X1 \core.keymem.key_mem[12][122]$_DFFE_PN0P_  (.D(_01246_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[12][122] ),
    .QN(_21358_));
 DFFR_X1 \core.keymem.key_mem[12][123]$_DFFE_PN0P_  (.D(_01247_),
    .RN(net93),
    .CK(clknet_leaf_196_clk),
    .Q(\core.keymem.key_mem[12][123] ),
    .QN(_21357_));
 DFFR_X1 \core.keymem.key_mem[12][124]$_DFFE_PN0P_  (.D(_01248_),
    .RN(net93),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[12][124] ),
    .QN(_21356_));
 DFFR_X1 \core.keymem.key_mem[12][125]$_DFFE_PN0P_  (.D(_01249_),
    .RN(net97),
    .CK(clknet_leaf_235_clk),
    .Q(\core.keymem.key_mem[12][125] ),
    .QN(_21355_));
 DFFR_X1 \core.keymem.key_mem[12][126]$_DFFE_PN0P_  (.D(_01250_),
    .RN(net98),
    .CK(clknet_leaf_167_clk),
    .Q(\core.keymem.key_mem[12][126] ),
    .QN(_21354_));
 DFFR_X1 \core.keymem.key_mem[12][127]$_DFFE_PN0P_  (.D(_01251_),
    .RN(net97),
    .CK(clknet_leaf_241_clk),
    .Q(\core.keymem.key_mem[12][127] ),
    .QN(_21353_));
 DFFR_X1 \core.keymem.key_mem[12][12]$_DFFE_PN0P_  (.D(_01252_),
    .RN(net93),
    .CK(clknet_leaf_206_clk),
    .Q(\core.keymem.key_mem[12][12] ),
    .QN(_21352_));
 DFFR_X1 \core.keymem.key_mem[12][13]$_DFFE_PN0P_  (.D(_01253_),
    .RN(net87),
    .CK(clknet_leaf_32_clk),
    .Q(\core.keymem.key_mem[12][13] ),
    .QN(_21351_));
 DFFR_X2 \core.keymem.key_mem[12][14]$_DFFE_PN0P_  (.D(_01254_),
    .RN(net94),
    .CK(clknet_leaf_209_clk),
    .Q(\core.keymem.key_mem[12][14] ),
    .QN(_21350_));
 DFFR_X1 \core.keymem.key_mem[12][15]$_DFFE_PN0P_  (.D(_01255_),
    .RN(net96),
    .CK(clknet_leaf_165_clk),
    .Q(\core.keymem.key_mem[12][15] ),
    .QN(_21349_));
 DFFR_X1 \core.keymem.key_mem[12][16]$_DFFE_PN0P_  (.D(_01256_),
    .RN(net89),
    .CK(clknet_leaf_34_clk),
    .Q(\core.keymem.key_mem[12][16] ),
    .QN(_21348_));
 DFFR_X1 \core.keymem.key_mem[12][17]$_DFFE_PN0P_  (.D(_01257_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[12][17] ),
    .QN(_21347_));
 DFFR_X1 \core.keymem.key_mem[12][18]$_DFFE_PN0P_  (.D(_01258_),
    .RN(net82),
    .CK(clknet_leaf_34_clk),
    .Q(\core.keymem.key_mem[12][18] ),
    .QN(_21346_));
 DFFR_X1 \core.keymem.key_mem[12][19]$_DFFE_PN0P_  (.D(_01259_),
    .RN(net89),
    .CK(clknet_leaf_65_clk),
    .Q(\core.keymem.key_mem[12][19] ),
    .QN(_21345_));
 DFFR_X1 \core.keymem.key_mem[12][1]$_DFFE_PN0P_  (.D(_01260_),
    .RN(net100),
    .CK(clknet_leaf_22_clk),
    .Q(\core.keymem.key_mem[12][1] ),
    .QN(_21344_));
 DFFR_X1 \core.keymem.key_mem[12][20]$_DFFE_PN0P_  (.D(_01261_),
    .RN(net82),
    .CK(clknet_leaf_23_clk),
    .Q(\core.keymem.key_mem[12][20] ),
    .QN(_21343_));
 DFFR_X1 \core.keymem.key_mem[12][21]$_DFFE_PN0P_  (.D(_01262_),
    .RN(net85),
    .CK(clknet_leaf_66_clk),
    .Q(\core.keymem.key_mem[12][21] ),
    .QN(_21342_));
 DFFR_X1 \core.keymem.key_mem[12][22]$_DFFE_PN0P_  (.D(_01263_),
    .RN(net94),
    .CK(clknet_leaf_220_clk),
    .Q(\core.keymem.key_mem[12][22] ),
    .QN(_21341_));
 DFFR_X1 \core.keymem.key_mem[12][23]$_DFFE_PN0P_  (.D(_01264_),
    .RN(net89),
    .CK(clknet_leaf_55_clk),
    .Q(\core.keymem.key_mem[12][23] ),
    .QN(_21340_));
 DFFR_X1 \core.keymem.key_mem[12][24]$_DFFE_PN0P_  (.D(_01265_),
    .RN(net89),
    .CK(clknet_leaf_65_clk),
    .Q(\core.keymem.key_mem[12][24] ),
    .QN(_21339_));
 DFFR_X1 \core.keymem.key_mem[12][25]$_DFFE_PN0P_  (.D(_01266_),
    .RN(net85),
    .CK(clknet_leaf_48_clk),
    .Q(\core.keymem.key_mem[12][25] ),
    .QN(_21338_));
 DFFR_X1 \core.keymem.key_mem[12][26]$_DFFE_PN0P_  (.D(_01267_),
    .RN(net89),
    .CK(clknet_leaf_21_clk),
    .Q(\core.keymem.key_mem[12][26] ),
    .QN(_21337_));
 DFFR_X1 \core.keymem.key_mem[12][27]$_DFFE_PN0P_  (.D(_01268_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[12][27] ),
    .QN(_21336_));
 DFFR_X1 \core.keymem.key_mem[12][28]$_DFFE_PN0P_  (.D(_01269_),
    .RN(net16),
    .CK(clknet_leaf_131_clk),
    .Q(\core.keymem.key_mem[12][28] ),
    .QN(_21335_));
 DFFR_X1 \core.keymem.key_mem[12][29]$_DFFE_PN0P_  (.D(_01270_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[12][29] ),
    .QN(_21334_));
 DFFR_X1 \core.keymem.key_mem[12][2]$_DFFE_PN0P_  (.D(_01271_),
    .RN(net89),
    .CK(clknet_leaf_64_clk),
    .Q(\core.keymem.key_mem[12][2] ),
    .QN(_21333_));
 DFFR_X1 \core.keymem.key_mem[12][30]$_DFFE_PN0P_  (.D(_01272_),
    .RN(net98),
    .CK(clknet_leaf_149_clk),
    .Q(\core.keymem.key_mem[12][30] ),
    .QN(_21332_));
 DFFR_X1 \core.keymem.key_mem[12][31]$_DFFE_PN0P_  (.D(_01273_),
    .RN(net16),
    .CK(clknet_leaf_138_clk),
    .Q(\core.keymem.key_mem[12][31] ),
    .QN(_21331_));
 DFFR_X1 \core.keymem.key_mem[12][32]$_DFFE_PN0P_  (.D(_01274_),
    .RN(net100),
    .CK(clknet_leaf_113_clk),
    .Q(\core.keymem.key_mem[12][32] ),
    .QN(_21330_));
 DFFR_X1 \core.keymem.key_mem[12][33]$_DFFE_PN0P_  (.D(_01275_),
    .RN(net99),
    .CK(clknet_leaf_112_clk),
    .Q(\core.keymem.key_mem[12][33] ),
    .QN(_21329_));
 DFFR_X1 \core.keymem.key_mem[12][34]$_DFFE_PN0P_  (.D(_01276_),
    .RN(net16),
    .CK(clknet_leaf_124_clk),
    .Q(\core.keymem.key_mem[12][34] ),
    .QN(_21328_));
 DFFR_X1 \core.keymem.key_mem[12][35]$_DFFE_PN0P_  (.D(_01277_),
    .RN(net99),
    .CK(clknet_leaf_128_clk),
    .Q(\core.keymem.key_mem[12][35] ),
    .QN(_21327_));
 DFFR_X1 \core.keymem.key_mem[12][36]$_DFFE_PN0P_  (.D(_01278_),
    .RN(net88),
    .CK(clknet_leaf_91_clk),
    .Q(\core.keymem.key_mem[12][36] ),
    .QN(_21326_));
 DFFR_X1 \core.keymem.key_mem[12][37]$_DFFE_PN0P_  (.D(_01279_),
    .RN(net88),
    .CK(clknet_leaf_93_clk),
    .Q(\core.keymem.key_mem[12][37] ),
    .QN(_21325_));
 DFFR_X1 \core.keymem.key_mem[12][38]$_DFFE_PN0P_  (.D(_01280_),
    .RN(net99),
    .CK(clknet_leaf_123_clk),
    .Q(\core.keymem.key_mem[12][38] ),
    .QN(_21324_));
 DFFR_X1 \core.keymem.key_mem[12][39]$_DFFE_PN0P_  (.D(_01281_),
    .RN(net89),
    .CK(clknet_leaf_86_clk),
    .Q(\core.keymem.key_mem[12][39] ),
    .QN(_21323_));
 DFFR_X1 \core.keymem.key_mem[12][3]$_DFFE_PN0P_  (.D(_01282_),
    .RN(net88),
    .CK(clknet_leaf_91_clk),
    .Q(\core.keymem.key_mem[12][3] ),
    .QN(_21322_));
 DFFR_X1 \core.keymem.key_mem[12][40]$_DFFE_PN0P_  (.D(_01283_),
    .RN(net88),
    .CK(clknet_leaf_90_clk),
    .Q(\core.keymem.key_mem[12][40] ),
    .QN(_21321_));
 DFFR_X1 \core.keymem.key_mem[12][41]$_DFFE_PN0P_  (.D(_01284_),
    .RN(net100),
    .CK(clknet_leaf_114_clk),
    .Q(\core.keymem.key_mem[12][41] ),
    .QN(_21320_));
 DFFR_X1 \core.keymem.key_mem[12][42]$_DFFE_PN0P_  (.D(_01285_),
    .RN(net100),
    .CK(clknet_leaf_128_clk),
    .Q(\core.keymem.key_mem[12][42] ),
    .QN(_21319_));
 DFFR_X1 \core.keymem.key_mem[12][43]$_DFFE_PN0P_  (.D(_01286_),
    .RN(net85),
    .CK(clknet_leaf_68_clk),
    .Q(\core.keymem.key_mem[12][43] ),
    .QN(_21318_));
 DFFR_X1 \core.keymem.key_mem[12][44]$_DFFE_PN0P_  (.D(_01287_),
    .RN(net100),
    .CK(clknet_leaf_108_clk),
    .Q(\core.keymem.key_mem[12][44] ),
    .QN(_21317_));
 DFFR_X1 \core.keymem.key_mem[12][45]$_DFFE_PN0P_  (.D(_01288_),
    .RN(net89),
    .CK(clknet_leaf_68_clk),
    .Q(\core.keymem.key_mem[12][45] ),
    .QN(_21316_));
 DFFR_X1 \core.keymem.key_mem[12][46]$_DFFE_PN0P_  (.D(_01289_),
    .RN(net89),
    .CK(clknet_leaf_83_clk),
    .Q(\core.keymem.key_mem[12][46] ),
    .QN(_21315_));
 DFFR_X1 \core.keymem.key_mem[12][47]$_DFFE_PN0P_  (.D(_01290_),
    .RN(net98),
    .CK(clknet_leaf_145_clk),
    .Q(\core.keymem.key_mem[12][47] ),
    .QN(_21314_));
 DFFR_X1 \core.keymem.key_mem[12][48]$_DFFE_PN0P_  (.D(_01291_),
    .RN(net95),
    .CK(clknet_leaf_117_clk),
    .Q(\core.keymem.key_mem[12][48] ),
    .QN(_21313_));
 DFFR_X1 \core.keymem.key_mem[12][49]$_DFFE_PN0P_  (.D(_01292_),
    .RN(net99),
    .CK(clknet_leaf_81_clk),
    .Q(\core.keymem.key_mem[12][49] ),
    .QN(_21312_));
 DFFR_X1 \core.keymem.key_mem[12][4]$_DFFE_PN0P_  (.D(_01293_),
    .RN(net100),
    .CK(clknet_leaf_106_clk),
    .Q(\core.keymem.key_mem[12][4] ),
    .QN(_21311_));
 DFFR_X1 \core.keymem.key_mem[12][50]$_DFFE_PN0P_  (.D(_01294_),
    .RN(net98),
    .CK(clknet_leaf_140_clk),
    .Q(\core.keymem.key_mem[12][50] ),
    .QN(_21310_));
 DFFR_X1 \core.keymem.key_mem[12][51]$_DFFE_PN0P_  (.D(_01295_),
    .RN(net100),
    .CK(clknet_leaf_130_clk),
    .Q(\core.keymem.key_mem[12][51] ),
    .QN(_21309_));
 DFFR_X1 \core.keymem.key_mem[12][52]$_DFFE_PN0P_  (.D(_01296_),
    .RN(net99),
    .CK(clknet_leaf_81_clk),
    .Q(\core.keymem.key_mem[12][52] ),
    .QN(_21308_));
 DFFR_X1 \core.keymem.key_mem[12][53]$_DFFE_PN0P_  (.D(_01297_),
    .RN(net98),
    .CK(clknet_leaf_145_clk),
    .Q(\core.keymem.key_mem[12][53] ),
    .QN(_21307_));
 DFFR_X1 \core.keymem.key_mem[12][54]$_DFFE_PN0P_  (.D(_01298_),
    .RN(net98),
    .CK(clknet_leaf_143_clk),
    .Q(\core.keymem.key_mem[12][54] ),
    .QN(_21306_));
 DFFR_X1 \core.keymem.key_mem[12][55]$_DFFE_PN0P_  (.D(_01299_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[12][55] ),
    .QN(_21305_));
 DFFR_X1 \core.keymem.key_mem[12][56]$_DFFE_PN0P_  (.D(_01300_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[12][56] ),
    .QN(_21304_));
 DFFR_X1 \core.keymem.key_mem[12][57]$_DFFE_PN0P_  (.D(_01301_),
    .RN(net100),
    .CK(clknet_leaf_109_clk),
    .Q(\core.keymem.key_mem[12][57] ),
    .QN(_21303_));
 DFFR_X1 \core.keymem.key_mem[12][58]$_DFFE_PN0P_  (.D(_01302_),
    .RN(net100),
    .CK(clknet_leaf_107_clk),
    .Q(\core.keymem.key_mem[12][58] ),
    .QN(_21302_));
 DFFR_X1 \core.keymem.key_mem[12][59]$_DFFE_PN0P_  (.D(_01303_),
    .RN(net100),
    .CK(clknet_leaf_17_clk),
    .Q(\core.keymem.key_mem[12][59] ),
    .QN(_21301_));
 DFFR_X1 \core.keymem.key_mem[12][5]$_DFFE_PN0P_  (.D(_01304_),
    .RN(net100),
    .CK(clknet_leaf_19_clk),
    .Q(\core.keymem.key_mem[12][5] ),
    .QN(_21300_));
 DFFR_X1 \core.keymem.key_mem[12][60]$_DFFE_PN0P_  (.D(_01305_),
    .RN(net82),
    .CK(clknet_leaf_13_clk),
    .Q(\core.keymem.key_mem[12][60] ),
    .QN(_21299_));
 DFFR_X1 \core.keymem.key_mem[12][61]$_DFFE_PN0P_  (.D(_01306_),
    .RN(net89),
    .CK(clknet_leaf_94_clk),
    .Q(\core.keymem.key_mem[12][61] ),
    .QN(_21298_));
 DFFR_X1 \core.keymem.key_mem[12][62]$_DFFE_PN0P_  (.D(_01307_),
    .RN(net100),
    .CK(clknet_leaf_98_clk),
    .Q(\core.keymem.key_mem[12][62] ),
    .QN(_21297_));
 DFFR_X1 \core.keymem.key_mem[12][63]$_DFFE_PN0P_  (.D(_01308_),
    .RN(net100),
    .CK(clknet_leaf_97_clk),
    .Q(\core.keymem.key_mem[12][63] ),
    .QN(_21296_));
 DFFR_X1 \core.keymem.key_mem[12][64]$_DFFE_PN0P_  (.D(_01309_),
    .RN(net100),
    .CK(clknet_leaf_14_clk),
    .Q(\core.keymem.key_mem[12][64] ),
    .QN(_21295_));
 DFFR_X1 \core.keymem.key_mem[12][65]$_DFFE_PN0P_  (.D(_01310_),
    .RN(net98),
    .CK(clknet_leaf_123_clk),
    .Q(\core.keymem.key_mem[12][65] ),
    .QN(_21294_));
 DFFR_X1 \core.keymem.key_mem[12][66]$_DFFE_PN0P_  (.D(_01311_),
    .RN(net100),
    .CK(clknet_leaf_16_clk),
    .Q(\core.keymem.key_mem[12][66] ),
    .QN(_21293_));
 DFFR_X1 \core.keymem.key_mem[12][67]$_DFFE_PN0P_  (.D(_01312_),
    .RN(net95),
    .CK(clknet_leaf_76_clk),
    .Q(\core.keymem.key_mem[12][67] ),
    .QN(_21292_));
 DFFR_X1 \core.keymem.key_mem[12][68]$_DFFE_PN0P_  (.D(_01313_),
    .RN(net99),
    .CK(clknet_leaf_117_clk),
    .Q(\core.keymem.key_mem[12][68] ),
    .QN(_21291_));
 DFFR_X1 \core.keymem.key_mem[12][69]$_DFFE_PN0P_  (.D(_01314_),
    .RN(net98),
    .CK(clknet_leaf_142_clk),
    .Q(\core.keymem.key_mem[12][69] ),
    .QN(_21290_));
 DFFR_X1 \core.keymem.key_mem[12][6]$_DFFE_PN0P_  (.D(_01315_),
    .RN(net100),
    .CK(clknet_leaf_102_clk),
    .Q(\core.keymem.key_mem[12][6] ),
    .QN(_21289_));
 DFFR_X1 \core.keymem.key_mem[12][70]$_DFFE_PN0P_  (.D(_01316_),
    .RN(net100),
    .CK(clknet_leaf_101_clk),
    .Q(\core.keymem.key_mem[12][70] ),
    .QN(_21288_));
 DFFR_X1 \core.keymem.key_mem[12][71]$_DFFE_PN0P_  (.D(_01317_),
    .RN(net99),
    .CK(clknet_leaf_74_clk),
    .Q(\core.keymem.key_mem[12][71] ),
    .QN(_21287_));
 DFFR_X1 \core.keymem.key_mem[12][72]$_DFFE_PN0P_  (.D(_01318_),
    .RN(net95),
    .CK(clknet_leaf_178_clk),
    .Q(\core.keymem.key_mem[12][72] ),
    .QN(_21286_));
 DFFR_X1 \core.keymem.key_mem[12][73]$_DFFE_PN0P_  (.D(_01319_),
    .RN(net97),
    .CK(clknet_leaf_147_clk),
    .Q(\core.keymem.key_mem[12][73] ),
    .QN(_21285_));
 DFFR_X1 \core.keymem.key_mem[12][74]$_DFFE_PN0P_  (.D(_01320_),
    .RN(net97),
    .CK(clknet_leaf_154_clk),
    .Q(\core.keymem.key_mem[12][74] ),
    .QN(_21284_));
 DFFR_X1 \core.keymem.key_mem[12][75]$_DFFE_PN0P_  (.D(_01321_),
    .RN(net97),
    .CK(clknet_leaf_148_clk),
    .Q(\core.keymem.key_mem[12][75] ),
    .QN(_21283_));
 DFFR_X1 \core.keymem.key_mem[12][76]$_DFFE_PN0P_  (.D(_01322_),
    .RN(net93),
    .CK(clknet_leaf_285_clk),
    .Q(\core.keymem.key_mem[12][76] ),
    .QN(_21282_));
 DFFR_X1 \core.keymem.key_mem[12][77]$_DFFE_PN0P_  (.D(_01323_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[12][77] ),
    .QN(_21281_));
 DFFR_X1 \core.keymem.key_mem[12][78]$_DFFE_PN0P_  (.D(_01324_),
    .RN(net98),
    .CK(clknet_leaf_174_clk),
    .Q(\core.keymem.key_mem[12][78] ),
    .QN(_21280_));
 DFFR_X1 \core.keymem.key_mem[12][79]$_DFFE_PN0P_  (.D(_01325_),
    .RN(net96),
    .CK(clknet_leaf_228_clk),
    .Q(\core.keymem.key_mem[12][79] ),
    .QN(_21279_));
 DFFR_X1 \core.keymem.key_mem[12][7]$_DFFE_PN0P_  (.D(_01326_),
    .RN(net98),
    .CK(clknet_leaf_172_clk),
    .Q(\core.keymem.key_mem[12][7] ),
    .QN(_21278_));
 DFFR_X1 \core.keymem.key_mem[12][80]$_DFFE_PN0P_  (.D(_01327_),
    .RN(net97),
    .CK(clknet_leaf_159_clk),
    .Q(\core.keymem.key_mem[12][80] ),
    .QN(_21277_));
 DFFR_X1 \core.keymem.key_mem[12][81]$_DFFE_PN0P_  (.D(_01328_),
    .RN(net97),
    .CK(clknet_leaf_155_clk),
    .Q(\core.keymem.key_mem[12][81] ),
    .QN(_21276_));
 DFFR_X1 \core.keymem.key_mem[12][82]$_DFFE_PN0P_  (.D(_01329_),
    .RN(net98),
    .CK(clknet_leaf_175_clk),
    .Q(\core.keymem.key_mem[12][82] ),
    .QN(_21275_));
 DFFR_X1 \core.keymem.key_mem[12][83]$_DFFE_PN0P_  (.D(_01330_),
    .RN(net95),
    .CK(clknet_leaf_183_clk),
    .Q(\core.keymem.key_mem[12][83] ),
    .QN(_21274_));
 DFFR_X1 \core.keymem.key_mem[12][84]$_DFFE_PN0P_  (.D(_01331_),
    .RN(net95),
    .CK(clknet_leaf_72_clk),
    .Q(\core.keymem.key_mem[12][84] ),
    .QN(_21273_));
 DFFR_X1 \core.keymem.key_mem[12][85]$_DFFE_PN0P_  (.D(_01332_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[12][85] ),
    .QN(_21272_));
 DFFR_X1 \core.keymem.key_mem[12][86]$_DFFE_PN0P_  (.D(_01333_),
    .RN(net95),
    .CK(clknet_leaf_208_clk),
    .Q(\core.keymem.key_mem[12][86] ),
    .QN(_21271_));
 DFFR_X1 \core.keymem.key_mem[12][87]$_DFFE_PN0P_  (.D(_01334_),
    .RN(net89),
    .CK(clknet_leaf_378_clk),
    .Q(\core.keymem.key_mem[12][87] ),
    .QN(_21270_));
 DFFR_X1 \core.keymem.key_mem[12][88]$_DFFE_PN0P_  (.D(_01335_),
    .RN(net91),
    .CK(clknet_leaf_283_clk),
    .Q(\core.keymem.key_mem[12][88] ),
    .QN(_21269_));
 DFFR_X1 \core.keymem.key_mem[12][89]$_DFFE_PN0P_  (.D(_01336_),
    .RN(net93),
    .CK(clknet_leaf_199_clk),
    .Q(\core.keymem.key_mem[12][89] ),
    .QN(_21268_));
 DFFR_X1 \core.keymem.key_mem[12][8]$_DFFE_PN0P_  (.D(_01337_),
    .RN(net93),
    .CK(clknet_leaf_377_clk),
    .Q(\core.keymem.key_mem[12][8] ),
    .QN(_21267_));
 DFFR_X1 \core.keymem.key_mem[12][90]$_DFFE_PN0P_  (.D(_01338_),
    .RN(net97),
    .CK(clknet_leaf_162_clk),
    .Q(\core.keymem.key_mem[12][90] ),
    .QN(_21266_));
 DFFR_X1 \core.keymem.key_mem[12][91]$_DFFE_PN0P_  (.D(_01339_),
    .RN(net95),
    .CK(clknet_leaf_183_clk),
    .Q(\core.keymem.key_mem[12][91] ),
    .QN(_21265_));
 DFFR_X1 \core.keymem.key_mem[12][92]$_DFFE_PN0P_  (.D(_01340_),
    .RN(net95),
    .CK(clknet_leaf_62_clk),
    .Q(\core.keymem.key_mem[12][92] ),
    .QN(_21264_));
 DFFR_X1 \core.keymem.key_mem[12][93]$_DFFE_PN0P_  (.D(_01341_),
    .RN(net98),
    .CK(clknet_leaf_166_clk),
    .Q(\core.keymem.key_mem[12][93] ),
    .QN(_21263_));
 DFFR_X1 \core.keymem.key_mem[12][94]$_DFFE_PN0P_  (.D(_01342_),
    .RN(net94),
    .CK(clknet_leaf_218_clk),
    .Q(\core.keymem.key_mem[12][94] ),
    .QN(_21262_));
 DFFR_X1 \core.keymem.key_mem[12][95]$_DFFE_PN0P_  (.D(_01343_),
    .RN(net96),
    .CK(clknet_leaf_244_clk),
    .Q(\core.keymem.key_mem[12][95] ),
    .QN(_21261_));
 DFFR_X1 \core.keymem.key_mem[12][96]$_DFFE_PN0P_  (.D(_01344_),
    .RN(net92),
    .CK(clknet_leaf_204_clk),
    .Q(\core.keymem.key_mem[12][96] ),
    .QN(_21260_));
 DFFR_X1 \core.keymem.key_mem[12][97]$_DFFE_PN0P_  (.D(_01345_),
    .RN(net93),
    .CK(clknet_leaf_193_clk),
    .Q(\core.keymem.key_mem[12][97] ),
    .QN(_21259_));
 DFFR_X1 \core.keymem.key_mem[12][98]$_DFFE_PN0P_  (.D(_01346_),
    .RN(net93),
    .CK(clknet_leaf_195_clk),
    .Q(\core.keymem.key_mem[12][98] ),
    .QN(_21258_));
 DFFR_X1 \core.keymem.key_mem[12][99]$_DFFE_PN0P_  (.D(_01347_),
    .RN(net91),
    .CK(clknet_leaf_201_clk),
    .Q(\core.keymem.key_mem[12][99] ),
    .QN(_21257_));
 DFFR_X1 \core.keymem.key_mem[12][9]$_DFFE_PN0P_  (.D(_01348_),
    .RN(net92),
    .CK(clknet_leaf_202_clk),
    .Q(\core.keymem.key_mem[12][9] ),
    .QN(_21256_));
 DFFR_X1 \core.keymem.key_mem[13][0]$_DFFE_PN0P_  (.D(_01349_),
    .RN(net96),
    .CK(clknet_leaf_247_clk),
    .Q(\core.keymem.key_mem[13][0] ),
    .QN(_21255_));
 DFFR_X1 \core.keymem.key_mem[13][100]$_DFFE_PN0P_  (.D(_01350_),
    .RN(net98),
    .CK(clknet_leaf_210_clk),
    .Q(\core.keymem.key_mem[13][100] ),
    .QN(_21254_));
 DFFR_X1 \core.keymem.key_mem[13][101]$_DFFE_PN0P_  (.D(_01351_),
    .RN(net94),
    .CK(clknet_leaf_218_clk),
    .Q(\core.keymem.key_mem[13][101] ),
    .QN(_21253_));
 DFFR_X1 \core.keymem.key_mem[13][102]$_DFFE_PN0P_  (.D(_01352_),
    .RN(net96),
    .CK(clknet_leaf_232_clk),
    .Q(\core.keymem.key_mem[13][102] ),
    .QN(_21252_));
 DFFR_X1 \core.keymem.key_mem[13][103]$_DFFE_PN0P_  (.D(_01353_),
    .RN(net96),
    .CK(clknet_leaf_234_clk),
    .Q(\core.keymem.key_mem[13][103] ),
    .QN(_21251_));
 DFFR_X1 \core.keymem.key_mem[13][104]$_DFFE_PN0P_  (.D(_01354_),
    .RN(net93),
    .CK(clknet_leaf_192_clk),
    .Q(\core.keymem.key_mem[13][104] ),
    .QN(_21250_));
 DFFR_X1 \core.keymem.key_mem[13][105]$_DFFE_PN0P_  (.D(_01355_),
    .RN(net96),
    .CK(clknet_leaf_245_clk),
    .Q(\core.keymem.key_mem[13][105] ),
    .QN(_21249_));
 DFFR_X1 \core.keymem.key_mem[13][106]$_DFFE_PN0P_  (.D(_01356_),
    .RN(net92),
    .CK(clknet_leaf_269_clk),
    .Q(\core.keymem.key_mem[13][106] ),
    .QN(_21248_));
 DFFR_X1 \core.keymem.key_mem[13][107]$_DFFE_PN0P_  (.D(_01357_),
    .RN(net92),
    .CK(clknet_leaf_276_clk),
    .Q(\core.keymem.key_mem[13][107] ),
    .QN(_21247_));
 DFFR_X1 \core.keymem.key_mem[13][108]$_DFFE_PN0P_  (.D(_01358_),
    .RN(net91),
    .CK(clknet_leaf_277_clk),
    .Q(\core.keymem.key_mem[13][108] ),
    .QN(_21246_));
 DFFR_X1 \core.keymem.key_mem[13][109]$_DFFE_PN0P_  (.D(_01359_),
    .RN(net94),
    .CK(clknet_leaf_259_clk),
    .Q(\core.keymem.key_mem[13][109] ),
    .QN(_21245_));
 DFFR_X1 \core.keymem.key_mem[13][10]$_DFFE_PN0P_  (.D(_01360_),
    .RN(net94),
    .CK(clknet_leaf_187_clk),
    .Q(\core.keymem.key_mem[13][10] ),
    .QN(_21244_));
 DFFR_X1 \core.keymem.key_mem[13][110]$_DFFE_PN0P_  (.D(_01361_),
    .RN(net96),
    .CK(clknet_leaf_250_clk),
    .Q(\core.keymem.key_mem[13][110] ),
    .QN(_21243_));
 DFFR_X1 \core.keymem.key_mem[13][111]$_DFFE_PN0P_  (.D(_01362_),
    .RN(net96),
    .CK(clknet_leaf_227_clk),
    .Q(\core.keymem.key_mem[13][111] ),
    .QN(_21242_));
 DFFR_X1 \core.keymem.key_mem[13][112]$_DFFE_PN0P_  (.D(_01363_),
    .RN(net94),
    .CK(clknet_leaf_260_clk),
    .Q(\core.keymem.key_mem[13][112] ),
    .QN(_21241_));
 DFFR_X1 \core.keymem.key_mem[13][113]$_DFFE_PN0P_  (.D(_01364_),
    .RN(net92),
    .CK(clknet_leaf_272_clk),
    .Q(\core.keymem.key_mem[13][113] ),
    .QN(_21240_));
 DFFR_X1 \core.keymem.key_mem[13][114]$_DFFE_PN0P_  (.D(_01365_),
    .RN(net91),
    .CK(clknet_leaf_274_clk),
    .Q(\core.keymem.key_mem[13][114] ),
    .QN(_21239_));
 DFFR_X1 \core.keymem.key_mem[13][115]$_DFFE_PN0P_  (.D(_01366_),
    .RN(net92),
    .CK(clknet_leaf_274_clk),
    .Q(\core.keymem.key_mem[13][115] ),
    .QN(_21238_));
 DFFR_X1 \core.keymem.key_mem[13][116]$_DFFE_PN0P_  (.D(_01367_),
    .RN(net94),
    .CK(clknet_leaf_265_clk),
    .Q(\core.keymem.key_mem[13][116] ),
    .QN(_21237_));
 DFFR_X1 \core.keymem.key_mem[13][117]$_DFFE_PN0P_  (.D(_01368_),
    .RN(net96),
    .CK(clknet_leaf_222_clk),
    .Q(\core.keymem.key_mem[13][117] ),
    .QN(_21236_));
 DFFR_X1 \core.keymem.key_mem[13][118]$_DFFE_PN0P_  (.D(_01369_),
    .RN(net97),
    .CK(clknet_leaf_240_clk),
    .Q(\core.keymem.key_mem[13][118] ),
    .QN(_21235_));
 DFFR_X1 \core.keymem.key_mem[13][119]$_DFFE_PN0P_  (.D(_01370_),
    .RN(net94),
    .CK(clknet_leaf_262_clk),
    .Q(\core.keymem.key_mem[13][119] ),
    .QN(_21234_));
 DFFR_X1 \core.keymem.key_mem[13][11]$_DFFE_PN0P_  (.D(_01371_),
    .RN(net95),
    .CK(clknet_leaf_61_clk),
    .Q(\core.keymem.key_mem[13][11] ),
    .QN(_21233_));
 DFFR_X1 \core.keymem.key_mem[13][120]$_DFFE_PN0P_  (.D(_01372_),
    .RN(net94),
    .CK(clknet_leaf_216_clk),
    .Q(\core.keymem.key_mem[13][120] ),
    .QN(_21232_));
 DFFR_X1 \core.keymem.key_mem[13][121]$_DFFE_PN0P_  (.D(_01373_),
    .RN(net92),
    .CK(clknet_leaf_265_clk),
    .Q(\core.keymem.key_mem[13][121] ),
    .QN(_21231_));
 DFFR_X1 \core.keymem.key_mem[13][122]$_DFFE_PN0P_  (.D(_01374_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[13][122] ),
    .QN(_21230_));
 DFFR_X1 \core.keymem.key_mem[13][123]$_DFFE_PN0P_  (.D(_01375_),
    .RN(net93),
    .CK(clknet_leaf_196_clk),
    .Q(\core.keymem.key_mem[13][123] ),
    .QN(_21229_));
 DFFR_X1 \core.keymem.key_mem[13][124]$_DFFE_PN0P_  (.D(_01376_),
    .RN(net93),
    .CK(clknet_leaf_198_clk),
    .Q(\core.keymem.key_mem[13][124] ),
    .QN(_21228_));
 DFFR_X1 \core.keymem.key_mem[13][125]$_DFFE_PN0P_  (.D(_01377_),
    .RN(net97),
    .CK(clknet_leaf_236_clk),
    .Q(\core.keymem.key_mem[13][125] ),
    .QN(_21227_));
 DFFR_X1 \core.keymem.key_mem[13][126]$_DFFE_PN0P_  (.D(_01378_),
    .RN(net98),
    .CK(clknet_leaf_188_clk),
    .Q(\core.keymem.key_mem[13][126] ),
    .QN(_21226_));
 DFFR_X1 \core.keymem.key_mem[13][127]$_DFFE_PN0P_  (.D(_01379_),
    .RN(net97),
    .CK(clknet_leaf_240_clk),
    .Q(\core.keymem.key_mem[13][127] ),
    .QN(_21225_));
 DFFR_X1 \core.keymem.key_mem[13][12]$_DFFE_PN0P_  (.D(_01380_),
    .RN(net93),
    .CK(clknet_leaf_208_clk),
    .Q(\core.keymem.key_mem[13][12] ),
    .QN(_21224_));
 DFFR_X1 \core.keymem.key_mem[13][13]$_DFFE_PN0P_  (.D(_01381_),
    .RN(net88),
    .CK(clknet_leaf_31_clk),
    .Q(\core.keymem.key_mem[13][13] ),
    .QN(_21223_));
 DFFR_X1 \core.keymem.key_mem[13][14]$_DFFE_PN0P_  (.D(_01382_),
    .RN(net98),
    .CK(clknet_leaf_229_clk),
    .Q(\core.keymem.key_mem[13][14] ),
    .QN(_21222_));
 DFFR_X1 \core.keymem.key_mem[13][15]$_DFFE_PN0P_  (.D(_01383_),
    .RN(net96),
    .CK(clknet_leaf_171_clk),
    .Q(\core.keymem.key_mem[13][15] ),
    .QN(_21221_));
 DFFR_X1 \core.keymem.key_mem[13][16]$_DFFE_PN0P_  (.D(_01384_),
    .RN(net89),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[13][16] ),
    .QN(_21220_));
 DFFR_X1 \core.keymem.key_mem[13][17]$_DFFE_PN0P_  (.D(_01385_),
    .RN(net98),
    .CK(clknet_leaf_186_clk),
    .Q(\core.keymem.key_mem[13][17] ),
    .QN(_21219_));
 DFFR_X1 \core.keymem.key_mem[13][18]$_DFFE_PN0P_  (.D(_01386_),
    .RN(net88),
    .CK(clknet_leaf_26_clk),
    .Q(\core.keymem.key_mem[13][18] ),
    .QN(_21218_));
 DFFR_X1 \core.keymem.key_mem[13][19]$_DFFE_PN0P_  (.D(_01387_),
    .RN(net85),
    .CK(clknet_leaf_54_clk),
    .Q(\core.keymem.key_mem[13][19] ),
    .QN(_21217_));
 DFFR_X1 \core.keymem.key_mem[13][1]$_DFFE_PN0P_  (.D(_01388_),
    .RN(net89),
    .CK(clknet_leaf_22_clk),
    .Q(\core.keymem.key_mem[13][1] ),
    .QN(_21216_));
 DFFR_X1 \core.keymem.key_mem[13][20]$_DFFE_PN0P_  (.D(_01389_),
    .RN(net100),
    .CK(clknet_leaf_21_clk),
    .Q(\core.keymem.key_mem[13][20] ),
    .QN(_21215_));
 DFFR_X1 \core.keymem.key_mem[13][21]$_DFFE_PN0P_  (.D(_01390_),
    .RN(net89),
    .CK(clknet_leaf_66_clk),
    .Q(\core.keymem.key_mem[13][21] ),
    .QN(_21214_));
 DFFR_X1 \core.keymem.key_mem[13][22]$_DFFE_PN0P_  (.D(_01391_),
    .RN(net96),
    .CK(clknet_leaf_222_clk),
    .Q(\core.keymem.key_mem[13][22] ),
    .QN(_21213_));
 DFFR_X1 \core.keymem.key_mem[13][23]$_DFFE_PN0P_  (.D(_01392_),
    .RN(net89),
    .CK(clknet_leaf_55_clk),
    .Q(\core.keymem.key_mem[13][23] ),
    .QN(_21212_));
 DFFR_X1 \core.keymem.key_mem[13][24]$_DFFE_PN0P_  (.D(_01393_),
    .RN(net89),
    .CK(clknet_leaf_59_clk),
    .Q(\core.keymem.key_mem[13][24] ),
    .QN(_21211_));
 DFFR_X1 \core.keymem.key_mem[13][25]$_DFFE_PN0P_  (.D(_01394_),
    .RN(net85),
    .CK(clknet_leaf_48_clk),
    .Q(\core.keymem.key_mem[13][25] ),
    .QN(_21210_));
 DFFR_X1 \core.keymem.key_mem[13][26]$_DFFE_PN0P_  (.D(_01395_),
    .RN(net89),
    .CK(clknet_leaf_96_clk),
    .Q(\core.keymem.key_mem[13][26] ),
    .QN(_21209_));
 DFFR_X1 \core.keymem.key_mem[13][27]$_DFFE_PN0P_  (.D(_01396_),
    .RN(net16),
    .CK(clknet_leaf_132_clk),
    .Q(\core.keymem.key_mem[13][27] ),
    .QN(_21208_));
 DFFR_X1 \core.keymem.key_mem[13][28]$_DFFE_PN0P_  (.D(_01397_),
    .RN(net16),
    .CK(clknet_leaf_126_clk),
    .Q(\core.keymem.key_mem[13][28] ),
    .QN(_21207_));
 DFFR_X1 \core.keymem.key_mem[13][29]$_DFFE_PN0P_  (.D(_01398_),
    .RN(net16),
    .CK(clknet_leaf_132_clk),
    .Q(\core.keymem.key_mem[13][29] ),
    .QN(_21206_));
 DFFR_X1 \core.keymem.key_mem[13][2]$_DFFE_PN0P_  (.D(_01399_),
    .RN(net89),
    .CK(clknet_leaf_60_clk),
    .Q(\core.keymem.key_mem[13][2] ),
    .QN(_21205_));
 DFFR_X1 \core.keymem.key_mem[13][30]$_DFFE_PN0P_  (.D(_01400_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[13][30] ),
    .QN(_21204_));
 DFFR_X1 \core.keymem.key_mem[13][31]$_DFFE_PN0P_  (.D(_01401_),
    .RN(net16),
    .CK(clknet_leaf_138_clk),
    .Q(\core.keymem.key_mem[13][31] ),
    .QN(_21203_));
 DFFR_X1 \core.keymem.key_mem[13][32]$_DFFE_PN0P_  (.D(_01402_),
    .RN(net100),
    .CK(clknet_leaf_113_clk),
    .Q(\core.keymem.key_mem[13][32] ),
    .QN(_21202_));
 DFFR_X1 \core.keymem.key_mem[13][33]$_DFFE_PN0P_  (.D(_01403_),
    .RN(net99),
    .CK(clknet_leaf_126_clk),
    .Q(\core.keymem.key_mem[13][33] ),
    .QN(_21201_));
 DFFR_X1 \core.keymem.key_mem[13][34]$_DFFE_PN0P_  (.D(_01404_),
    .RN(net16),
    .CK(clknet_leaf_123_clk),
    .Q(\core.keymem.key_mem[13][34] ),
    .QN(_21200_));
 DFFR_X1 \core.keymem.key_mem[13][35]$_DFFE_PN0P_  (.D(_01405_),
    .RN(net99),
    .CK(clknet_leaf_111_clk),
    .Q(\core.keymem.key_mem[13][35] ),
    .QN(_21199_));
 DFFR_X1 \core.keymem.key_mem[13][36]$_DFFE_PN0P_  (.D(_01406_),
    .RN(net88),
    .CK(clknet_leaf_27_clk),
    .Q(\core.keymem.key_mem[13][36] ),
    .QN(_21198_));
 DFFR_X1 \core.keymem.key_mem[13][37]$_DFFE_PN0P_  (.D(_01407_),
    .RN(net89),
    .CK(clknet_leaf_93_clk),
    .Q(\core.keymem.key_mem[13][37] ),
    .QN(_21197_));
 DFFR_X1 \core.keymem.key_mem[13][38]$_DFFE_PN0P_  (.D(_01408_),
    .RN(net16),
    .CK(clknet_leaf_123_clk),
    .Q(\core.keymem.key_mem[13][38] ),
    .QN(_21196_));
 DFFR_X1 \core.keymem.key_mem[13][39]$_DFFE_PN0P_  (.D(_01409_),
    .RN(net99),
    .CK(clknet_leaf_70_clk),
    .Q(\core.keymem.key_mem[13][39] ),
    .QN(_21195_));
 DFFR_X1 \core.keymem.key_mem[13][3]$_DFFE_PN0P_  (.D(_01410_),
    .RN(net88),
    .CK(clknet_leaf_27_clk),
    .Q(\core.keymem.key_mem[13][3] ),
    .QN(_21194_));
 DFFR_X1 \core.keymem.key_mem[13][40]$_DFFE_PN0P_  (.D(_01411_),
    .RN(net85),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[13][40] ),
    .QN(_21193_));
 DFFR_X1 \core.keymem.key_mem[13][41]$_DFFE_PN0P_  (.D(_01412_),
    .RN(net89),
    .CK(clknet_leaf_83_clk),
    .Q(\core.keymem.key_mem[13][41] ),
    .QN(_21192_));
 DFFR_X1 \core.keymem.key_mem[13][42]$_DFFE_PN0P_  (.D(_01413_),
    .RN(net100),
    .CK(clknet_leaf_111_clk),
    .Q(\core.keymem.key_mem[13][42] ),
    .QN(_21191_));
 DFFR_X1 \core.keymem.key_mem[13][43]$_DFFE_PN0P_  (.D(_01414_),
    .RN(net85),
    .CK(clknet_leaf_88_clk),
    .Q(\core.keymem.key_mem[13][43] ),
    .QN(_21190_));
 DFFR_X1 \core.keymem.key_mem[13][44]$_DFFE_PN0P_  (.D(_01415_),
    .RN(net100),
    .CK(clknet_leaf_107_clk),
    .Q(\core.keymem.key_mem[13][44] ),
    .QN(_21189_));
 DFFR_X1 \core.keymem.key_mem[13][45]$_DFFE_PN0P_  (.D(_01416_),
    .RN(net89),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[13][45] ),
    .QN(_21188_));
 DFFR_X1 \core.keymem.key_mem[13][46]$_DFFE_PN0P_  (.D(_01417_),
    .RN(net99),
    .CK(clknet_leaf_82_clk),
    .Q(\core.keymem.key_mem[13][46] ),
    .QN(_21187_));
 DFFR_X1 \core.keymem.key_mem[13][47]$_DFFE_PN0P_  (.D(_01418_),
    .RN(net98),
    .CK(clknet_leaf_176_clk),
    .Q(\core.keymem.key_mem[13][47] ),
    .QN(_21186_));
 DFFR_X1 \core.keymem.key_mem[13][48]$_DFFE_PN0P_  (.D(_01419_),
    .RN(net99),
    .CK(clknet_leaf_119_clk),
    .Q(\core.keymem.key_mem[13][48] ),
    .QN(_21185_));
 DFFR_X1 \core.keymem.key_mem[13][49]$_DFFE_PN0P_  (.D(_01420_),
    .RN(net99),
    .CK(clknet_leaf_116_clk),
    .Q(\core.keymem.key_mem[13][49] ),
    .QN(_21184_));
 DFFR_X1 \core.keymem.key_mem[13][4]$_DFFE_PN0P_  (.D(_01421_),
    .RN(net100),
    .CK(clknet_leaf_105_clk),
    .Q(\core.keymem.key_mem[13][4] ),
    .QN(_21183_));
 DFFR_X1 \core.keymem.key_mem[13][50]$_DFFE_PN0P_  (.D(_01422_),
    .RN(net98),
    .CK(clknet_leaf_140_clk),
    .Q(\core.keymem.key_mem[13][50] ),
    .QN(_21182_));
 DFFR_X1 \core.keymem.key_mem[13][51]$_DFFE_PN0P_  (.D(_01423_),
    .RN(net100),
    .CK(clknet_leaf_129_clk),
    .Q(\core.keymem.key_mem[13][51] ),
    .QN(_21181_));
 DFFR_X1 \core.keymem.key_mem[13][52]$_DFFE_PN0P_  (.D(_01424_),
    .RN(net99),
    .CK(clknet_leaf_81_clk),
    .Q(\core.keymem.key_mem[13][52] ),
    .QN(_21180_));
 DFFR_X1 \core.keymem.key_mem[13][53]$_DFFE_PN0P_  (.D(_01425_),
    .RN(net98),
    .CK(clknet_leaf_176_clk),
    .Q(\core.keymem.key_mem[13][53] ),
    .QN(_21179_));
 DFFR_X1 \core.keymem.key_mem[13][54]$_DFFE_PN0P_  (.D(_01426_),
    .RN(net98),
    .CK(clknet_leaf_141_clk),
    .Q(\core.keymem.key_mem[13][54] ),
    .QN(_21178_));
 DFFR_X1 \core.keymem.key_mem[13][55]$_DFFE_PN0P_  (.D(_01427_),
    .RN(net16),
    .CK(clknet_leaf_135_clk),
    .Q(\core.keymem.key_mem[13][55] ),
    .QN(_21177_));
 DFFR_X1 \core.keymem.key_mem[13][56]$_DFFE_PN0P_  (.D(_01428_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[13][56] ),
    .QN(_21176_));
 DFFR_X1 \core.keymem.key_mem[13][57]$_DFFE_PN0P_  (.D(_01429_),
    .RN(net100),
    .CK(clknet_leaf_108_clk),
    .Q(\core.keymem.key_mem[13][57] ),
    .QN(_21175_));
 DFFR_X1 \core.keymem.key_mem[13][58]$_DFFE_PN0P_  (.D(_01430_),
    .RN(net100),
    .CK(clknet_leaf_106_clk),
    .Q(\core.keymem.key_mem[13][58] ),
    .QN(_21174_));
 DFFR_X1 \core.keymem.key_mem[13][59]$_DFFE_PN0P_  (.D(_01431_),
    .RN(net100),
    .CK(clknet_leaf_18_clk),
    .Q(\core.keymem.key_mem[13][59] ),
    .QN(_21173_));
 DFFR_X1 \core.keymem.key_mem[13][5]$_DFFE_PN0P_  (.D(_01432_),
    .RN(net100),
    .CK(clknet_leaf_18_clk),
    .Q(\core.keymem.key_mem[13][5] ),
    .QN(_21172_));
 DFFR_X1 \core.keymem.key_mem[13][60]$_DFFE_PN0P_  (.D(_01433_),
    .RN(net82),
    .CK(clknet_leaf_24_clk),
    .Q(\core.keymem.key_mem[13][60] ),
    .QN(_21171_));
 DFFR_X1 \core.keymem.key_mem[13][61]$_DFFE_PN0P_  (.D(_01434_),
    .RN(net88),
    .CK(clknet_leaf_93_clk),
    .Q(\core.keymem.key_mem[13][61] ),
    .QN(_21170_));
 DFFR_X1 \core.keymem.key_mem[13][62]$_DFFE_PN0P_  (.D(_01435_),
    .RN(net100),
    .CK(clknet_leaf_99_clk),
    .Q(\core.keymem.key_mem[13][62] ),
    .QN(_21169_));
 DFFR_X1 \core.keymem.key_mem[13][63]$_DFFE_PN0P_  (.D(_01436_),
    .RN(net100),
    .CK(clknet_leaf_97_clk),
    .Q(\core.keymem.key_mem[13][63] ),
    .QN(_21168_));
 DFFR_X1 \core.keymem.key_mem[13][64]$_DFFE_PN0P_  (.D(_01437_),
    .RN(net82),
    .CK(clknet_leaf_14_clk),
    .Q(\core.keymem.key_mem[13][64] ),
    .QN(_21167_));
 DFFR_X1 \core.keymem.key_mem[13][65]$_DFFE_PN0P_  (.D(_01438_),
    .RN(net99),
    .CK(clknet_leaf_120_clk),
    .Q(\core.keymem.key_mem[13][65] ),
    .QN(_21166_));
 DFFR_X1 \core.keymem.key_mem[13][66]$_DFFE_PN0P_  (.D(_01439_),
    .RN(net100),
    .CK(clknet_leaf_16_clk),
    .Q(\core.keymem.key_mem[13][66] ),
    .QN(_21165_));
 DFFR_X1 \core.keymem.key_mem[13][67]$_DFFE_PN0P_  (.D(_01440_),
    .RN(net95),
    .CK(clknet_leaf_77_clk),
    .Q(\core.keymem.key_mem[13][67] ),
    .QN(_21164_));
 DFFR_X1 \core.keymem.key_mem[13][68]$_DFFE_PN0P_  (.D(_01441_),
    .RN(net99),
    .CK(clknet_leaf_117_clk),
    .Q(\core.keymem.key_mem[13][68] ),
    .QN(_21163_));
 DFFR_X1 \core.keymem.key_mem[13][69]$_DFFE_PN0P_  (.D(_01442_),
    .RN(net95),
    .CK(clknet_leaf_178_clk),
    .Q(\core.keymem.key_mem[13][69] ),
    .QN(_21162_));
 DFFR_X1 \core.keymem.key_mem[13][6]$_DFFE_PN0P_  (.D(_01443_),
    .RN(net100),
    .CK(clknet_leaf_102_clk),
    .Q(\core.keymem.key_mem[13][6] ),
    .QN(_21161_));
 DFFR_X1 \core.keymem.key_mem[13][70]$_DFFE_PN0P_  (.D(_01444_),
    .RN(net100),
    .CK(clknet_leaf_100_clk),
    .Q(\core.keymem.key_mem[13][70] ),
    .QN(_21160_));
 DFFR_X1 \core.keymem.key_mem[13][71]$_DFFE_PN0P_  (.D(_01445_),
    .RN(net99),
    .CK(clknet_leaf_73_clk),
    .Q(\core.keymem.key_mem[13][71] ),
    .QN(_21159_));
 DFFR_X1 \core.keymem.key_mem[13][72]$_DFFE_PN0P_  (.D(_01446_),
    .RN(net95),
    .CK(clknet_leaf_178_clk),
    .Q(\core.keymem.key_mem[13][72] ),
    .QN(_21158_));
 DFFR_X1 \core.keymem.key_mem[13][73]$_DFFE_PN0P_  (.D(_01447_),
    .RN(net97),
    .CK(clknet_leaf_147_clk),
    .Q(\core.keymem.key_mem[13][73] ),
    .QN(_21157_));
 DFFR_X1 \core.keymem.key_mem[13][74]$_DFFE_PN0P_  (.D(_01448_),
    .RN(net97),
    .CK(clknet_leaf_157_clk),
    .Q(\core.keymem.key_mem[13][74] ),
    .QN(_21156_));
 DFFR_X1 \core.keymem.key_mem[13][75]$_DFFE_PN0P_  (.D(_01449_),
    .RN(net97),
    .CK(clknet_leaf_152_clk),
    .Q(\core.keymem.key_mem[13][75] ),
    .QN(_21155_));
 DFFR_X1 \core.keymem.key_mem[13][76]$_DFFE_PN0P_  (.D(_01450_),
    .RN(net93),
    .CK(clknet_leaf_283_clk),
    .Q(\core.keymem.key_mem[13][76] ),
    .QN(_21154_));
 DFFR_X1 \core.keymem.key_mem[13][77]$_DFFE_PN0P_  (.D(_01451_),
    .RN(net97),
    .CK(clknet_leaf_159_clk),
    .Q(\core.keymem.key_mem[13][77] ),
    .QN(_21153_));
 DFFR_X1 \core.keymem.key_mem[13][78]$_DFFE_PN0P_  (.D(_01452_),
    .RN(net97),
    .CK(clknet_leaf_172_clk),
    .Q(\core.keymem.key_mem[13][78] ),
    .QN(_21152_));
 DFFR_X1 \core.keymem.key_mem[13][79]$_DFFE_PN0P_  (.D(_01453_),
    .RN(net96),
    .CK(clknet_leaf_230_clk),
    .Q(\core.keymem.key_mem[13][79] ),
    .QN(_21151_));
 DFFR_X1 \core.keymem.key_mem[13][7]$_DFFE_PN0P_  (.D(_01454_),
    .RN(net98),
    .CK(clknet_leaf_170_clk),
    .Q(\core.keymem.key_mem[13][7] ),
    .QN(_21150_));
 DFFR_X1 \core.keymem.key_mem[13][80]$_DFFE_PN0P_  (.D(_01455_),
    .RN(net97),
    .CK(clknet_leaf_157_clk),
    .Q(\core.keymem.key_mem[13][80] ),
    .QN(_21149_));
 DFFR_X1 \core.keymem.key_mem[13][81]$_DFFE_PN0P_  (.D(_01456_),
    .RN(net97),
    .CK(clknet_leaf_153_clk),
    .Q(\core.keymem.key_mem[13][81] ),
    .QN(_21148_));
 DFFR_X1 \core.keymem.key_mem[13][82]$_DFFE_PN0P_  (.D(_01457_),
    .RN(net98),
    .CK(clknet_leaf_180_clk),
    .Q(\core.keymem.key_mem[13][82] ),
    .QN(_21147_));
 DFFR_X1 \core.keymem.key_mem[13][83]$_DFFE_PN0P_  (.D(_01458_),
    .RN(net94),
    .CK(clknet_leaf_181_clk),
    .Q(\core.keymem.key_mem[13][83] ),
    .QN(_21146_));
 DFFR_X1 \core.keymem.key_mem[13][84]$_DFFE_PN0P_  (.D(_01459_),
    .RN(net95),
    .CK(clknet_leaf_179_clk),
    .Q(\core.keymem.key_mem[13][84] ),
    .QN(_21145_));
 DFFR_X1 \core.keymem.key_mem[13][85]$_DFFE_PN0P_  (.D(_01460_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[13][85] ),
    .QN(_21144_));
 DFFR_X1 \core.keymem.key_mem[13][86]$_DFFE_PN0P_  (.D(_01461_),
    .RN(net97),
    .CK(clknet_leaf_160_clk),
    .Q(\core.keymem.key_mem[13][86] ),
    .QN(_21143_));
 DFFR_X1 \core.keymem.key_mem[13][87]$_DFFE_PN0P_  (.D(_01462_),
    .RN(net93),
    .CK(clknet_leaf_56_clk),
    .Q(\core.keymem.key_mem[13][87] ),
    .QN(_21142_));
 DFFR_X1 \core.keymem.key_mem[13][88]$_DFFE_PN0P_  (.D(_01463_),
    .RN(net93),
    .CK(clknet_leaf_282_clk),
    .Q(\core.keymem.key_mem[13][88] ),
    .QN(_21141_));
 DFFR_X1 \core.keymem.key_mem[13][89]$_DFFE_PN0P_  (.D(_01464_),
    .RN(net93),
    .CK(clknet_leaf_200_clk),
    .Q(\core.keymem.key_mem[13][89] ),
    .QN(_21140_));
 DFFR_X1 \core.keymem.key_mem[13][8]$_DFFE_PN0P_  (.D(_01465_),
    .RN(net89),
    .CK(clknet_leaf_378_clk),
    .Q(\core.keymem.key_mem[13][8] ),
    .QN(_21139_));
 DFFR_X1 \core.keymem.key_mem[13][90]$_DFFE_PN0P_  (.D(_01466_),
    .RN(net97),
    .CK(clknet_leaf_156_clk),
    .Q(\core.keymem.key_mem[13][90] ),
    .QN(_21138_));
 DFFR_X1 \core.keymem.key_mem[13][91]$_DFFE_PN0P_  (.D(_01467_),
    .RN(net94),
    .CK(clknet_leaf_186_clk),
    .Q(\core.keymem.key_mem[13][91] ),
    .QN(_21137_));
 DFFR_X1 \core.keymem.key_mem[13][92]$_DFFE_PN0P_  (.D(_01468_),
    .RN(net95),
    .CK(clknet_leaf_63_clk),
    .Q(\core.keymem.key_mem[13][92] ),
    .QN(_21136_));
 DFFR_X1 \core.keymem.key_mem[13][93]$_DFFE_PN0P_  (.D(_01469_),
    .RN(net98),
    .CK(clknet_leaf_189_clk),
    .Q(\core.keymem.key_mem[13][93] ),
    .QN(_21135_));
 DFFR_X1 \core.keymem.key_mem[13][94]$_DFFE_PN0P_  (.D(_01470_),
    .RN(net94),
    .CK(clknet_leaf_214_clk),
    .Q(\core.keymem.key_mem[13][94] ),
    .QN(_21134_));
 DFFR_X1 \core.keymem.key_mem[13][95]$_DFFE_PN0P_  (.D(_01471_),
    .RN(net96),
    .CK(clknet_leaf_242_clk),
    .Q(\core.keymem.key_mem[13][95] ),
    .QN(_21133_));
 DFFR_X1 \core.keymem.key_mem[13][96]$_DFFE_PN0P_  (.D(_01472_),
    .RN(net92),
    .CK(clknet_leaf_204_clk),
    .Q(\core.keymem.key_mem[13][96] ),
    .QN(_21132_));
 DFFR_X1 \core.keymem.key_mem[13][97]$_DFFE_PN0P_  (.D(_01473_),
    .RN(net93),
    .CK(clknet_leaf_194_clk),
    .Q(\core.keymem.key_mem[13][97] ),
    .QN(_21131_));
 DFFR_X1 \core.keymem.key_mem[13][98]$_DFFE_PN0P_  (.D(_01474_),
    .RN(net95),
    .CK(clknet_leaf_194_clk),
    .Q(\core.keymem.key_mem[13][98] ),
    .QN(_21130_));
 DFFR_X1 \core.keymem.key_mem[13][99]$_DFFE_PN0P_  (.D(_01475_),
    .RN(net92),
    .CK(clknet_leaf_207_clk),
    .Q(\core.keymem.key_mem[13][99] ),
    .QN(_21129_));
 DFFR_X1 \core.keymem.key_mem[13][9]$_DFFE_PN0P_  (.D(_01476_),
    .RN(net92),
    .CK(clknet_leaf_203_clk),
    .Q(\core.keymem.key_mem[13][9] ),
    .QN(_21128_));
 DFFR_X1 \core.keymem.key_mem[14][0]$_DFFE_PN0P_  (.D(_01477_),
    .RN(net96),
    .CK(clknet_leaf_248_clk),
    .Q(\core.keymem.key_mem[14][0] ),
    .QN(_21127_));
 DFFR_X1 \core.keymem.key_mem[14][100]$_DFFE_PN0P_  (.D(_01478_),
    .RN(net98),
    .CK(clknet_leaf_226_clk),
    .Q(\core.keymem.key_mem[14][100] ),
    .QN(_21126_));
 DFFR_X1 \core.keymem.key_mem[14][101]$_DFFE_PN0P_  (.D(_01479_),
    .RN(net96),
    .CK(clknet_leaf_245_clk),
    .Q(\core.keymem.key_mem[14][101] ),
    .QN(_21125_));
 DFFR_X1 \core.keymem.key_mem[14][102]$_DFFE_PN0P_  (.D(_01480_),
    .RN(net96),
    .CK(clknet_leaf_233_clk),
    .Q(\core.keymem.key_mem[14][102] ),
    .QN(_21124_));
 DFFR_X1 \core.keymem.key_mem[14][103]$_DFFE_PN0P_  (.D(_01481_),
    .RN(net96),
    .CK(clknet_leaf_245_clk),
    .Q(\core.keymem.key_mem[14][103] ),
    .QN(_21123_));
 DFFR_X1 \core.keymem.key_mem[14][104]$_DFFE_PN0P_  (.D(_01482_),
    .RN(net93),
    .CK(clknet_leaf_196_clk),
    .Q(\core.keymem.key_mem[14][104] ),
    .QN(_21122_));
 DFFR_X1 \core.keymem.key_mem[14][105]$_DFFE_PN0P_  (.D(_01483_),
    .RN(net96),
    .CK(clknet_leaf_245_clk),
    .Q(\core.keymem.key_mem[14][105] ),
    .QN(_21121_));
 DFFR_X1 \core.keymem.key_mem[14][106]$_DFFE_PN0P_  (.D(_01484_),
    .RN(net92),
    .CK(clknet_leaf_258_clk),
    .Q(\core.keymem.key_mem[14][106] ),
    .QN(_21120_));
 DFFR_X1 \core.keymem.key_mem[14][107]$_DFFE_PN0P_  (.D(_01485_),
    .RN(net92),
    .CK(clknet_leaf_270_clk),
    .Q(\core.keymem.key_mem[14][107] ),
    .QN(_21119_));
 DFFR_X1 \core.keymem.key_mem[14][108]$_DFFE_PN0P_  (.D(_01486_),
    .RN(net91),
    .CK(clknet_leaf_277_clk),
    .Q(\core.keymem.key_mem[14][108] ),
    .QN(_21118_));
 DFFR_X1 \core.keymem.key_mem[14][109]$_DFFE_PN0P_  (.D(_01487_),
    .RN(net94),
    .CK(clknet_leaf_260_clk),
    .Q(\core.keymem.key_mem[14][109] ),
    .QN(_21117_));
 DFFR_X1 \core.keymem.key_mem[14][10]$_DFFE_PN0P_  (.D(_01488_),
    .RN(net98),
    .CK(clknet_leaf_187_clk),
    .Q(\core.keymem.key_mem[14][10] ),
    .QN(_21116_));
 DFFR_X1 \core.keymem.key_mem[14][110]$_DFFE_PN0P_  (.D(_01489_),
    .RN(net96),
    .CK(clknet_leaf_250_clk),
    .Q(\core.keymem.key_mem[14][110] ),
    .QN(_21115_));
 DFFR_X1 \core.keymem.key_mem[14][111]$_DFFE_PN0P_  (.D(_01490_),
    .RN(net96),
    .CK(clknet_leaf_224_clk),
    .Q(\core.keymem.key_mem[14][111] ),
    .QN(_21114_));
 DFFR_X1 \core.keymem.key_mem[14][112]$_DFFE_PN0P_  (.D(_01491_),
    .RN(net94),
    .CK(clknet_leaf_261_clk),
    .Q(\core.keymem.key_mem[14][112] ),
    .QN(_21113_));
 DFFR_X1 \core.keymem.key_mem[14][113]$_DFFE_PN0P_  (.D(_01492_),
    .RN(net92),
    .CK(clknet_leaf_272_clk),
    .Q(\core.keymem.key_mem[14][113] ),
    .QN(_21112_));
 DFFR_X1 \core.keymem.key_mem[14][114]$_DFFE_PN0P_  (.D(_01493_),
    .RN(net91),
    .CK(clknet_leaf_278_clk),
    .Q(\core.keymem.key_mem[14][114] ),
    .QN(_21111_));
 DFFR_X1 \core.keymem.key_mem[14][115]$_DFFE_PN0P_  (.D(_01494_),
    .RN(net92),
    .CK(clknet_leaf_275_clk),
    .Q(\core.keymem.key_mem[14][115] ),
    .QN(_21110_));
 DFFR_X1 \core.keymem.key_mem[14][116]$_DFFE_PN0P_  (.D(_01495_),
    .RN(net94),
    .CK(clknet_leaf_262_clk),
    .Q(\core.keymem.key_mem[14][116] ),
    .QN(_21109_));
 DFFR_X1 \core.keymem.key_mem[14][117]$_DFFE_PN0P_  (.D(_01496_),
    .RN(net96),
    .CK(clknet_leaf_223_clk),
    .Q(\core.keymem.key_mem[14][117] ),
    .QN(_21108_));
 DFFR_X1 \core.keymem.key_mem[14][118]$_DFFE_PN0P_  (.D(_01497_),
    .RN(net97),
    .CK(clknet_leaf_244_clk),
    .Q(\core.keymem.key_mem[14][118] ),
    .QN(_21107_));
 DFFR_X1 \core.keymem.key_mem[14][119]$_DFFE_PN0P_  (.D(_01498_),
    .RN(net94),
    .CK(clknet_leaf_220_clk),
    .Q(\core.keymem.key_mem[14][119] ),
    .QN(_21106_));
 DFFR_X1 \core.keymem.key_mem[14][11]$_DFFE_PN0P_  (.D(_01499_),
    .RN(net95),
    .CK(clknet_leaf_61_clk),
    .Q(\core.keymem.key_mem[14][11] ),
    .QN(_21105_));
 DFFR_X1 \core.keymem.key_mem[14][120]$_DFFE_PN0P_  (.D(_01500_),
    .RN(net94),
    .CK(clknet_leaf_215_clk),
    .Q(\core.keymem.key_mem[14][120] ),
    .QN(_21104_));
 DFFR_X1 \core.keymem.key_mem[14][121]$_DFFE_PN0P_  (.D(_01501_),
    .RN(net94),
    .CK(clknet_leaf_265_clk),
    .Q(\core.keymem.key_mem[14][121] ),
    .QN(_21103_));
 DFFR_X1 \core.keymem.key_mem[14][122]$_DFFE_PN0P_  (.D(_01502_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[14][122] ),
    .QN(_21102_));
 DFFR_X1 \core.keymem.key_mem[14][123]$_DFFE_PN0P_  (.D(_01503_),
    .RN(net93),
    .CK(clknet_leaf_197_clk),
    .Q(\core.keymem.key_mem[14][123] ),
    .QN(_21101_));
 DFFR_X1 \core.keymem.key_mem[14][124]$_DFFE_PN0P_  (.D(_01504_),
    .RN(net93),
    .CK(clknet_leaf_198_clk),
    .Q(\core.keymem.key_mem[14][124] ),
    .QN(_21100_));
 DFFR_X1 \core.keymem.key_mem[14][125]$_DFFE_PN0P_  (.D(_01505_),
    .RN(net96),
    .CK(clknet_leaf_232_clk),
    .Q(\core.keymem.key_mem[14][125] ),
    .QN(_21099_));
 DFFR_X1 \core.keymem.key_mem[14][126]$_DFFE_PN0P_  (.D(_01506_),
    .RN(net98),
    .CK(clknet_leaf_166_clk),
    .Q(\core.keymem.key_mem[14][126] ),
    .QN(_21098_));
 DFFR_X1 \core.keymem.key_mem[14][127]$_DFFE_PN0P_  (.D(_01507_),
    .RN(net97),
    .CK(clknet_leaf_240_clk),
    .Q(\core.keymem.key_mem[14][127] ),
    .QN(_21097_));
 DFFR_X1 \core.keymem.key_mem[14][12]$_DFFE_PN0P_  (.D(_01508_),
    .RN(net93),
    .CK(clknet_leaf_206_clk),
    .Q(\core.keymem.key_mem[14][12] ),
    .QN(_21096_));
 DFFR_X1 \core.keymem.key_mem[14][13]$_DFFE_PN0P_  (.D(_01509_),
    .RN(net88),
    .CK(clknet_leaf_31_clk),
    .Q(\core.keymem.key_mem[14][13] ),
    .QN(_21095_));
 DFFR_X1 \core.keymem.key_mem[14][14]$_DFFE_PN0P_  (.D(_01510_),
    .RN(net94),
    .CK(clknet_leaf_211_clk),
    .Q(\core.keymem.key_mem[14][14] ),
    .QN(_21094_));
 DFFR_X1 \core.keymem.key_mem[14][15]$_DFFE_PN0P_  (.D(_01511_),
    .RN(net96),
    .CK(clknet_leaf_165_clk),
    .Q(\core.keymem.key_mem[14][15] ),
    .QN(_21093_));
 DFFR_X1 \core.keymem.key_mem[14][16]$_DFFE_PN0P_  (.D(_01512_),
    .RN(net89),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[14][16] ),
    .QN(_21092_));
 DFFR_X1 \core.keymem.key_mem[14][17]$_DFFE_PN0P_  (.D(_01513_),
    .RN(net98),
    .CK(clknet_leaf_168_clk),
    .Q(\core.keymem.key_mem[14][17] ),
    .QN(_21091_));
 DFFR_X1 \core.keymem.key_mem[14][18]$_DFFE_PN0P_  (.D(_01514_),
    .RN(net89),
    .CK(clknet_leaf_26_clk),
    .Q(\core.keymem.key_mem[14][18] ),
    .QN(_21090_));
 DFFR_X1 \core.keymem.key_mem[14][19]$_DFFE_PN0P_  (.D(_01515_),
    .RN(net89),
    .CK(clknet_leaf_59_clk),
    .Q(\core.keymem.key_mem[14][19] ),
    .QN(_21089_));
 DFFR_X1 \core.keymem.key_mem[14][1]$_DFFE_PN0P_  (.D(_01516_),
    .RN(net89),
    .CK(clknet_leaf_25_clk),
    .Q(\core.keymem.key_mem[14][1] ),
    .QN(_21088_));
 DFFR_X1 \core.keymem.key_mem[14][20]$_DFFE_PN0P_  (.D(_01517_),
    .RN(net100),
    .CK(clknet_leaf_21_clk),
    .Q(\core.keymem.key_mem[14][20] ),
    .QN(_21087_));
 DFFR_X1 \core.keymem.key_mem[14][21]$_DFFE_PN0P_  (.D(_01518_),
    .RN(net85),
    .CK(clknet_leaf_68_clk),
    .Q(\core.keymem.key_mem[14][21] ),
    .QN(_21086_));
 DFFR_X1 \core.keymem.key_mem[14][22]$_DFFE_PN0P_  (.D(_01519_),
    .RN(net94),
    .CK(clknet_leaf_221_clk),
    .Q(\core.keymem.key_mem[14][22] ),
    .QN(_21085_));
 DFFR_X1 \core.keymem.key_mem[14][23]$_DFFE_PN0P_  (.D(_01520_),
    .RN(net89),
    .CK(clknet_leaf_54_clk),
    .Q(\core.keymem.key_mem[14][23] ),
    .QN(_21084_));
 DFFR_X1 \core.keymem.key_mem[14][24]$_DFFE_PN0P_  (.D(_01521_),
    .RN(net89),
    .CK(clknet_leaf_64_clk),
    .Q(\core.keymem.key_mem[14][24] ),
    .QN(_21083_));
 DFFR_X1 \core.keymem.key_mem[14][25]$_DFFE_PN0P_  (.D(_01522_),
    .RN(net85),
    .CK(clknet_leaf_47_clk),
    .Q(\core.keymem.key_mem[14][25] ),
    .QN(_21082_));
 DFFR_X1 \core.keymem.key_mem[14][26]$_DFFE_PN0P_  (.D(_01523_),
    .RN(net100),
    .CK(clknet_leaf_96_clk),
    .Q(\core.keymem.key_mem[14][26] ),
    .QN(_21081_));
 DFFR_X1 \core.keymem.key_mem[14][27]$_DFFE_PN0P_  (.D(_01524_),
    .RN(net16),
    .CK(clknet_leaf_151_clk),
    .Q(\core.keymem.key_mem[14][27] ),
    .QN(_21080_));
 DFFR_X1 \core.keymem.key_mem[14][28]$_DFFE_PN0P_  (.D(_01525_),
    .RN(net16),
    .CK(clknet_leaf_131_clk),
    .Q(\core.keymem.key_mem[14][28] ),
    .QN(_21079_));
 DFFR_X1 \core.keymem.key_mem[14][29]$_DFFE_PN0P_  (.D(_01526_),
    .RN(net16),
    .CK(clknet_leaf_132_clk),
    .Q(\core.keymem.key_mem[14][29] ),
    .QN(_21078_));
 DFFR_X1 \core.keymem.key_mem[14][2]$_DFFE_PN0P_  (.D(_01527_),
    .RN(net95),
    .CK(clknet_leaf_60_clk),
    .Q(\core.keymem.key_mem[14][2] ),
    .QN(_21077_));
 DFFR_X1 \core.keymem.key_mem[14][30]$_DFFE_PN0P_  (.D(_01528_),
    .RN(net98),
    .CK(clknet_leaf_149_clk),
    .Q(\core.keymem.key_mem[14][30] ),
    .QN(_21076_));
 DFFR_X1 \core.keymem.key_mem[14][31]$_DFFE_PN0P_  (.D(_01529_),
    .RN(net98),
    .CK(clknet_leaf_139_clk),
    .Q(\core.keymem.key_mem[14][31] ),
    .QN(_21075_));
 DFFR_X1 \core.keymem.key_mem[14][32]$_DFFE_PN0P_  (.D(_01530_),
    .RN(net100),
    .CK(clknet_leaf_110_clk),
    .Q(\core.keymem.key_mem[14][32] ),
    .QN(_21074_));
 DFFR_X1 \core.keymem.key_mem[14][33]$_DFFE_PN0P_  (.D(_01531_),
    .RN(net16),
    .CK(clknet_leaf_127_clk),
    .Q(\core.keymem.key_mem[14][33] ),
    .QN(_21073_));
 DFFR_X1 \core.keymem.key_mem[14][34]$_DFFE_PN0P_  (.D(_01532_),
    .RN(net16),
    .CK(clknet_leaf_136_clk),
    .Q(\core.keymem.key_mem[14][34] ),
    .QN(_21072_));
 DFFR_X1 \core.keymem.key_mem[14][35]$_DFFE_PN0P_  (.D(_01533_),
    .RN(net99),
    .CK(clknet_leaf_122_clk),
    .Q(\core.keymem.key_mem[14][35] ),
    .QN(_21071_));
 DFFR_X1 \core.keymem.key_mem[14][36]$_DFFE_PN0P_  (.D(_01534_),
    .RN(net88),
    .CK(clknet_leaf_89_clk),
    .Q(\core.keymem.key_mem[14][36] ),
    .QN(_21070_));
 DFFR_X1 \core.keymem.key_mem[14][37]$_DFFE_PN0P_  (.D(_01535_),
    .RN(net89),
    .CK(clknet_leaf_84_clk),
    .Q(\core.keymem.key_mem[14][37] ),
    .QN(_21069_));
 DFFR_X1 \core.keymem.key_mem[14][38]$_DFFE_PN0P_  (.D(_01536_),
    .RN(net99),
    .CK(clknet_leaf_127_clk),
    .Q(\core.keymem.key_mem[14][38] ),
    .QN(_21068_));
 DFFR_X1 \core.keymem.key_mem[14][39]$_DFFE_PN0P_  (.D(_01537_),
    .RN(net85),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[14][39] ),
    .QN(_21067_));
 DFFR_X1 \core.keymem.key_mem[14][3]$_DFFE_PN0P_  (.D(_01538_),
    .RN(net85),
    .CK(clknet_leaf_67_clk),
    .Q(\core.keymem.key_mem[14][3] ),
    .QN(_21066_));
 DFFR_X1 \core.keymem.key_mem[14][40]$_DFFE_PN0P_  (.D(_01539_),
    .RN(net88),
    .CK(clknet_leaf_89_clk),
    .Q(\core.keymem.key_mem[14][40] ),
    .QN(_21065_));
 DFFR_X1 \core.keymem.key_mem[14][41]$_DFFE_PN0P_  (.D(_01540_),
    .RN(net89),
    .CK(clknet_leaf_114_clk),
    .Q(\core.keymem.key_mem[14][41] ),
    .QN(_21064_));
 DFFR_X1 \core.keymem.key_mem[14][42]$_DFFE_PN0P_  (.D(_01541_),
    .RN(net100),
    .CK(clknet_leaf_111_clk),
    .Q(\core.keymem.key_mem[14][42] ),
    .QN(_21063_));
 DFFR_X1 \core.keymem.key_mem[14][43]$_DFFE_PN0P_  (.D(_01542_),
    .RN(net85),
    .CK(clknet_leaf_68_clk),
    .Q(\core.keymem.key_mem[14][43] ),
    .QN(_21062_));
 DFFR_X1 \core.keymem.key_mem[14][44]$_DFFE_PN0P_  (.D(_01543_),
    .RN(net100),
    .CK(clknet_leaf_105_clk),
    .Q(\core.keymem.key_mem[14][44] ),
    .QN(_21061_));
 DFFR_X1 \core.keymem.key_mem[14][45]$_DFFE_PN0P_  (.D(_01544_),
    .RN(net89),
    .CK(clknet_leaf_68_clk),
    .Q(\core.keymem.key_mem[14][45] ),
    .QN(_21060_));
 DFFR_X1 \core.keymem.key_mem[14][46]$_DFFE_PN0P_  (.D(_01545_),
    .RN(net99),
    .CK(clknet_leaf_79_clk),
    .Q(\core.keymem.key_mem[14][46] ),
    .QN(_21059_));
 DFFR_X1 \core.keymem.key_mem[14][47]$_DFFE_PN0P_  (.D(_01546_),
    .RN(net98),
    .CK(clknet_leaf_145_clk),
    .Q(\core.keymem.key_mem[14][47] ),
    .QN(_21058_));
 DFFR_X1 \core.keymem.key_mem[14][48]$_DFFE_PN0P_  (.D(_01547_),
    .RN(net98),
    .CK(clknet_leaf_141_clk),
    .Q(\core.keymem.key_mem[14][48] ),
    .QN(_21057_));
 DFFR_X1 \core.keymem.key_mem[14][49]$_DFFE_PN0P_  (.D(_01548_),
    .RN(net99),
    .CK(clknet_leaf_118_clk),
    .Q(\core.keymem.key_mem[14][49] ),
    .QN(_21056_));
 DFFR_X1 \core.keymem.key_mem[14][4]$_DFFE_PN0P_  (.D(_01549_),
    .RN(net100),
    .CK(clknet_leaf_105_clk),
    .Q(\core.keymem.key_mem[14][4] ),
    .QN(_21055_));
 DFFR_X1 \core.keymem.key_mem[14][50]$_DFFE_PN0P_  (.D(_01550_),
    .RN(net98),
    .CK(clknet_leaf_137_clk),
    .Q(\core.keymem.key_mem[14][50] ),
    .QN(_21054_));
 DFFR_X1 \core.keymem.key_mem[14][51]$_DFFE_PN0P_  (.D(_01551_),
    .RN(net100),
    .CK(clknet_leaf_129_clk),
    .Q(\core.keymem.key_mem[14][51] ),
    .QN(_21053_));
 DFFR_X1 \core.keymem.key_mem[14][52]$_DFFE_PN0P_  (.D(_01552_),
    .RN(net99),
    .CK(clknet_leaf_74_clk),
    .Q(\core.keymem.key_mem[14][52] ),
    .QN(_21052_));
 DFFR_X1 \core.keymem.key_mem[14][53]$_DFFE_PN0P_  (.D(_01553_),
    .RN(net98),
    .CK(clknet_leaf_145_clk),
    .Q(\core.keymem.key_mem[14][53] ),
    .QN(_21051_));
 DFFR_X1 \core.keymem.key_mem[14][54]$_DFFE_PN0P_  (.D(_01554_),
    .RN(net98),
    .CK(clknet_leaf_143_clk),
    .Q(\core.keymem.key_mem[14][54] ),
    .QN(_21050_));
 DFFR_X1 \core.keymem.key_mem[14][55]$_DFFE_PN0P_  (.D(_01555_),
    .RN(net16),
    .CK(clknet_leaf_135_clk),
    .Q(\core.keymem.key_mem[14][55] ),
    .QN(_21049_));
 DFFR_X1 \core.keymem.key_mem[14][56]$_DFFE_PN0P_  (.D(_01556_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[14][56] ),
    .QN(_21048_));
 DFFR_X1 \core.keymem.key_mem[14][57]$_DFFE_PN0P_  (.D(_01557_),
    .RN(net100),
    .CK(clknet_leaf_108_clk),
    .Q(\core.keymem.key_mem[14][57] ),
    .QN(_21047_));
 DFFR_X1 \core.keymem.key_mem[14][58]$_DFFE_PN0P_  (.D(_01558_),
    .RN(net100),
    .CK(clknet_leaf_107_clk),
    .Q(\core.keymem.key_mem[14][58] ),
    .QN(_21046_));
 DFFR_X1 \core.keymem.key_mem[14][59]$_DFFE_PN0P_  (.D(_01559_),
    .RN(net100),
    .CK(clknet_leaf_17_clk),
    .Q(\core.keymem.key_mem[14][59] ),
    .QN(_21045_));
 DFFR_X1 \core.keymem.key_mem[14][5]$_DFFE_PN0P_  (.D(_01560_),
    .RN(net100),
    .CK(clknet_leaf_19_clk),
    .Q(\core.keymem.key_mem[14][5] ),
    .QN(_21044_));
 DFFR_X1 \core.keymem.key_mem[14][60]$_DFFE_PN0P_  (.D(_01561_),
    .RN(net82),
    .CK(clknet_leaf_24_clk),
    .Q(\core.keymem.key_mem[14][60] ),
    .QN(_21043_));
 DFFR_X1 \core.keymem.key_mem[14][61]$_DFFE_PN0P_  (.D(_01562_),
    .RN(net89),
    .CK(clknet_leaf_94_clk),
    .Q(\core.keymem.key_mem[14][61] ),
    .QN(_21042_));
 DFFR_X1 \core.keymem.key_mem[14][62]$_DFFE_PN0P_  (.D(_01563_),
    .RN(net100),
    .CK(clknet_leaf_99_clk),
    .Q(\core.keymem.key_mem[14][62] ),
    .QN(_21041_));
 DFFR_X1 \core.keymem.key_mem[14][63]$_DFFE_PN0P_  (.D(_01564_),
    .RN(net100),
    .CK(clknet_leaf_103_clk),
    .Q(\core.keymem.key_mem[14][63] ),
    .QN(_21040_));
 DFFR_X1 \core.keymem.key_mem[14][64]$_DFFE_PN0P_  (.D(_01565_),
    .RN(net100),
    .CK(clknet_leaf_15_clk),
    .Q(\core.keymem.key_mem[14][64] ),
    .QN(_21039_));
 DFFR_X1 \core.keymem.key_mem[14][65]$_DFFE_PN0P_  (.D(_01566_),
    .RN(net98),
    .CK(clknet_leaf_121_clk),
    .Q(\core.keymem.key_mem[14][65] ),
    .QN(_21038_));
 DFFR_X1 \core.keymem.key_mem[14][66]$_DFFE_PN0P_  (.D(_01567_),
    .RN(net100),
    .CK(clknet_leaf_17_clk),
    .Q(\core.keymem.key_mem[14][66] ),
    .QN(_21037_));
 DFFR_X1 \core.keymem.key_mem[14][67]$_DFFE_PN0P_  (.D(_01568_),
    .RN(net95),
    .CK(clknet_leaf_178_clk),
    .Q(\core.keymem.key_mem[14][67] ),
    .QN(_21036_));
 DFFR_X1 \core.keymem.key_mem[14][68]$_DFFE_PN0P_  (.D(_01569_),
    .RN(net99),
    .CK(clknet_leaf_118_clk),
    .Q(\core.keymem.key_mem[14][68] ),
    .QN(_21035_));
 DFFR_X1 \core.keymem.key_mem[14][69]$_DFFE_PN0P_  (.D(_01570_),
    .RN(net95),
    .CK(clknet_leaf_177_clk),
    .Q(\core.keymem.key_mem[14][69] ),
    .QN(_21034_));
 DFFR_X1 \core.keymem.key_mem[14][6]$_DFFE_PN0P_  (.D(_01571_),
    .RN(net100),
    .CK(clknet_leaf_101_clk),
    .Q(\core.keymem.key_mem[14][6] ),
    .QN(_21033_));
 DFFR_X1 \core.keymem.key_mem[14][70]$_DFFE_PN0P_  (.D(_01572_),
    .RN(net100),
    .CK(clknet_leaf_98_clk),
    .Q(\core.keymem.key_mem[14][70] ),
    .QN(_21032_));
 DFFR_X1 \core.keymem.key_mem[14][71]$_DFFE_PN0P_  (.D(_01573_),
    .RN(net99),
    .CK(clknet_leaf_73_clk),
    .Q(\core.keymem.key_mem[14][71] ),
    .QN(_21031_));
 DFFR_X1 \core.keymem.key_mem[14][72]$_DFFE_PN0P_  (.D(_01574_),
    .RN(net95),
    .CK(clknet_leaf_76_clk),
    .Q(\core.keymem.key_mem[14][72] ),
    .QN(_21030_));
 DFFR_X1 \core.keymem.key_mem[14][73]$_DFFE_PN0P_  (.D(_01575_),
    .RN(net97),
    .CK(clknet_leaf_147_clk),
    .Q(\core.keymem.key_mem[14][73] ),
    .QN(_21029_));
 DFFR_X1 \core.keymem.key_mem[14][74]$_DFFE_PN0P_  (.D(_01576_),
    .RN(net97),
    .CK(clknet_leaf_155_clk),
    .Q(\core.keymem.key_mem[14][74] ),
    .QN(_21028_));
 DFFR_X1 \core.keymem.key_mem[14][75]$_DFFE_PN0P_  (.D(_01577_),
    .RN(net97),
    .CK(clknet_leaf_152_clk),
    .Q(\core.keymem.key_mem[14][75] ),
    .QN(_21027_));
 DFFR_X1 \core.keymem.key_mem[14][76]$_DFFE_PN0P_  (.D(_01578_),
    .RN(net93),
    .CK(clknet_leaf_282_clk),
    .Q(\core.keymem.key_mem[14][76] ),
    .QN(_21026_));
 DFFR_X1 \core.keymem.key_mem[14][77]$_DFFE_PN0P_  (.D(_01579_),
    .RN(net97),
    .CK(clknet_leaf_160_clk),
    .Q(\core.keymem.key_mem[14][77] ),
    .QN(_21025_));
 DFFR_X1 \core.keymem.key_mem[14][78]$_DFFE_PN0P_  (.D(_01580_),
    .RN(net97),
    .CK(clknet_leaf_164_clk),
    .Q(\core.keymem.key_mem[14][78] ),
    .QN(_21024_));
 DFFR_X1 \core.keymem.key_mem[14][79]$_DFFE_PN0P_  (.D(_01581_),
    .RN(net96),
    .CK(clknet_leaf_230_clk),
    .Q(\core.keymem.key_mem[14][79] ),
    .QN(_21023_));
 DFFR_X1 \core.keymem.key_mem[14][7]$_DFFE_PN0P_  (.D(_01582_),
    .RN(net98),
    .CK(clknet_leaf_174_clk),
    .Q(\core.keymem.key_mem[14][7] ),
    .QN(_21022_));
 DFFR_X1 \core.keymem.key_mem[14][80]$_DFFE_PN0P_  (.D(_01583_),
    .RN(net97),
    .CK(clknet_leaf_158_clk),
    .Q(\core.keymem.key_mem[14][80] ),
    .QN(_21021_));
 DFFR_X1 \core.keymem.key_mem[14][81]$_DFFE_PN0P_  (.D(_01584_),
    .RN(net97),
    .CK(clknet_leaf_153_clk),
    .Q(\core.keymem.key_mem[14][81] ),
    .QN(_21020_));
 DFFR_X1 \core.keymem.key_mem[14][82]$_DFFE_PN0P_  (.D(_01585_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[14][82] ),
    .QN(_21019_));
 DFFR_X1 \core.keymem.key_mem[14][83]$_DFFE_PN0P_  (.D(_01586_),
    .RN(net95),
    .CK(clknet_leaf_185_clk),
    .Q(\core.keymem.key_mem[14][83] ),
    .QN(_21018_));
 DFFR_X1 \core.keymem.key_mem[14][84]$_DFFE_PN0P_  (.D(_01587_),
    .RN(net95),
    .CK(clknet_leaf_179_clk),
    .Q(\core.keymem.key_mem[14][84] ),
    .QN(_21017_));
 DFFR_X1 \core.keymem.key_mem[14][85]$_DFFE_PN0P_  (.D(_01588_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[14][85] ),
    .QN(_21016_));
 DFFR_X1 \core.keymem.key_mem[14][86]$_DFFE_PN0P_  (.D(_01589_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[14][86] ),
    .QN(_21015_));
 DFFR_X1 \core.keymem.key_mem[14][87]$_DFFE_PN0P_  (.D(_01590_),
    .RN(net89),
    .CK(clknet_leaf_56_clk),
    .Q(\core.keymem.key_mem[14][87] ),
    .QN(_21014_));
 DFFR_X1 \core.keymem.key_mem[14][88]$_DFFE_PN0P_  (.D(_01591_),
    .RN(net93),
    .CK(clknet_leaf_280_clk),
    .Q(\core.keymem.key_mem[14][88] ),
    .QN(_21013_));
 DFFR_X1 \core.keymem.key_mem[14][89]$_DFFE_PN0P_  (.D(_01592_),
    .RN(net93),
    .CK(clknet_leaf_199_clk),
    .Q(\core.keymem.key_mem[14][89] ),
    .QN(_21012_));
 DFFR_X1 \core.keymem.key_mem[14][8]$_DFFE_PN0P_  (.D(_01593_),
    .RN(net93),
    .CK(clknet_leaf_377_clk),
    .Q(\core.keymem.key_mem[14][8] ),
    .QN(_21011_));
 DFFR_X1 \core.keymem.key_mem[14][90]$_DFFE_PN0P_  (.D(_01594_),
    .RN(net97),
    .CK(clknet_leaf_163_clk),
    .Q(\core.keymem.key_mem[14][90] ),
    .QN(_21010_));
 DFFR_X1 \core.keymem.key_mem[14][91]$_DFFE_PN0P_  (.D(_01595_),
    .RN(net94),
    .CK(clknet_leaf_186_clk),
    .Q(\core.keymem.key_mem[14][91] ),
    .QN(_21009_));
 DFFR_X1 \core.keymem.key_mem[14][92]$_DFFE_PN0P_  (.D(_01596_),
    .RN(net95),
    .CK(clknet_leaf_62_clk),
    .Q(\core.keymem.key_mem[14][92] ),
    .QN(_21008_));
 DFFR_X1 \core.keymem.key_mem[14][93]$_DFFE_PN0P_  (.D(_01597_),
    .RN(net96),
    .CK(clknet_leaf_231_clk),
    .Q(\core.keymem.key_mem[14][93] ),
    .QN(_21007_));
 DFFR_X1 \core.keymem.key_mem[14][94]$_DFFE_PN0P_  (.D(_01598_),
    .RN(net96),
    .CK(clknet_leaf_226_clk),
    .Q(\core.keymem.key_mem[14][94] ),
    .QN(_21006_));
 DFFR_X1 \core.keymem.key_mem[14][95]$_DFFE_PN0P_  (.D(_01599_),
    .RN(net96),
    .CK(clknet_leaf_242_clk),
    .Q(\core.keymem.key_mem[14][95] ),
    .QN(_21005_));
 DFFR_X1 \core.keymem.key_mem[14][96]$_DFFE_PN0P_  (.D(_01600_),
    .RN(net92),
    .CK(clknet_leaf_216_clk),
    .Q(\core.keymem.key_mem[14][96] ),
    .QN(_21004_));
 DFFR_X1 \core.keymem.key_mem[14][97]$_DFFE_PN0P_  (.D(_01601_),
    .RN(net93),
    .CK(clknet_leaf_193_clk),
    .Q(\core.keymem.key_mem[14][97] ),
    .QN(_21003_));
 DFFR_X1 \core.keymem.key_mem[14][98]$_DFFE_PN0P_  (.D(_01602_),
    .RN(net93),
    .CK(clknet_leaf_193_clk),
    .Q(\core.keymem.key_mem[14][98] ),
    .QN(_21002_));
 DFFR_X1 \core.keymem.key_mem[14][99]$_DFFE_PN0P_  (.D(_01603_),
    .RN(net92),
    .CK(clknet_leaf_207_clk),
    .Q(\core.keymem.key_mem[14][99] ),
    .QN(_21001_));
 DFFR_X1 \core.keymem.key_mem[14][9]$_DFFE_PN0P_  (.D(_01604_),
    .RN(net92),
    .CK(clknet_leaf_207_clk),
    .Q(\core.keymem.key_mem[14][9] ),
    .QN(_21000_));
 DFFR_X1 \core.keymem.key_mem[1][0]$_DFFE_PN0P_  (.D(_01605_),
    .RN(net96),
    .CK(clknet_leaf_221_clk),
    .Q(\core.keymem.key_mem[1][0] ),
    .QN(_20999_));
 DFFR_X1 \core.keymem.key_mem[1][100]$_DFFE_PN0P_  (.D(_01606_),
    .RN(net94),
    .CK(clknet_leaf_210_clk),
    .Q(\core.keymem.key_mem[1][100] ),
    .QN(_20998_));
 DFFR_X1 \core.keymem.key_mem[1][101]$_DFFE_PN0P_  (.D(_01607_),
    .RN(net94),
    .CK(clknet_leaf_212_clk),
    .Q(\core.keymem.key_mem[1][101] ),
    .QN(_20997_));
 DFFR_X1 \core.keymem.key_mem[1][102]$_DFFE_PN0P_  (.D(_01608_),
    .RN(net96),
    .CK(clknet_leaf_230_clk),
    .Q(\core.keymem.key_mem[1][102] ),
    .QN(_20996_));
 DFFR_X1 \core.keymem.key_mem[1][103]$_DFFE_PN0P_  (.D(_01609_),
    .RN(net96),
    .CK(clknet_leaf_224_clk),
    .Q(\core.keymem.key_mem[1][103] ),
    .QN(_20995_));
 DFFR_X1 \core.keymem.key_mem[1][104]$_DFFE_PN0P_  (.D(_01610_),
    .RN(net92),
    .CK(clknet_leaf_192_clk),
    .Q(\core.keymem.key_mem[1][104] ),
    .QN(_20994_));
 DFFR_X1 \core.keymem.key_mem[1][105]$_DFFE_PN0P_  (.D(_01611_),
    .RN(net96),
    .CK(clknet_leaf_223_clk),
    .Q(\core.keymem.key_mem[1][105] ),
    .QN(_20993_));
 DFFR_X1 \core.keymem.key_mem[1][106]$_DFFE_PN0P_  (.D(_01612_),
    .RN(net92),
    .CK(clknet_leaf_276_clk),
    .Q(\core.keymem.key_mem[1][106] ),
    .QN(_20992_));
 DFFR_X1 \core.keymem.key_mem[1][107]$_DFFE_PN0P_  (.D(_01613_),
    .RN(net92),
    .CK(clknet_leaf_276_clk),
    .Q(\core.keymem.key_mem[1][107] ),
    .QN(_20991_));
 DFFR_X1 \core.keymem.key_mem[1][108]$_DFFE_PN0P_  (.D(_01614_),
    .RN(net91),
    .CK(clknet_leaf_280_clk),
    .Q(\core.keymem.key_mem[1][108] ),
    .QN(_20990_));
 DFFR_X1 \core.keymem.key_mem[1][109]$_DFFE_PN0P_  (.D(_01615_),
    .RN(net94),
    .CK(clknet_leaf_264_clk),
    .Q(\core.keymem.key_mem[1][109] ),
    .QN(_20989_));
 DFFR_X2 \core.keymem.key_mem[1][10]$_DFFE_PN0P_  (.D(_01616_),
    .RN(net89),
    .CK(clknet_leaf_53_clk),
    .Q(\core.keymem.key_mem[1][10] ),
    .QN(_20988_));
 DFFR_X1 \core.keymem.key_mem[1][110]$_DFFE_PN0P_  (.D(_01617_),
    .RN(net96),
    .CK(clknet_leaf_213_clk),
    .Q(\core.keymem.key_mem[1][110] ),
    .QN(_20987_));
 DFFR_X1 \core.keymem.key_mem[1][111]$_DFFE_PN0P_  (.D(_01618_),
    .RN(net96),
    .CK(clknet_leaf_225_clk),
    .Q(\core.keymem.key_mem[1][111] ),
    .QN(_20986_));
 DFFR_X1 \core.keymem.key_mem[1][112]$_DFFE_PN0P_  (.D(_01619_),
    .RN(net94),
    .CK(clknet_leaf_262_clk),
    .Q(\core.keymem.key_mem[1][112] ),
    .QN(_20985_));
 DFFR_X1 \core.keymem.key_mem[1][113]$_DFFE_PN0P_  (.D(_01620_),
    .RN(net91),
    .CK(clknet_leaf_279_clk),
    .Q(\core.keymem.key_mem[1][113] ),
    .QN(_20984_));
 DFFR_X1 \core.keymem.key_mem[1][114]$_DFFE_PN0P_  (.D(_01621_),
    .RN(net91),
    .CK(clknet_leaf_279_clk),
    .Q(\core.keymem.key_mem[1][114] ),
    .QN(_20983_));
 DFFR_X1 \core.keymem.key_mem[1][115]$_DFFE_PN0P_  (.D(_01622_),
    .RN(net92),
    .CK(clknet_leaf_275_clk),
    .Q(\core.keymem.key_mem[1][115] ),
    .QN(_20982_));
 DFFR_X1 \core.keymem.key_mem[1][116]$_DFFE_PN0P_  (.D(_01623_),
    .RN(net94),
    .CK(clknet_leaf_264_clk),
    .Q(\core.keymem.key_mem[1][116] ),
    .QN(_20981_));
 DFFR_X1 \core.keymem.key_mem[1][117]$_DFFE_PN0P_  (.D(_01624_),
    .RN(net94),
    .CK(clknet_leaf_213_clk),
    .Q(\core.keymem.key_mem[1][117] ),
    .QN(_20980_));
 DFFR_X1 \core.keymem.key_mem[1][118]$_DFFE_PN0P_  (.D(_01625_),
    .RN(net96),
    .CK(clknet_leaf_228_clk),
    .Q(\core.keymem.key_mem[1][118] ),
    .QN(_20979_));
 DFFR_X1 \core.keymem.key_mem[1][119]$_DFFE_PN0P_  (.D(_01626_),
    .RN(net94),
    .CK(clknet_leaf_219_clk),
    .Q(\core.keymem.key_mem[1][119] ),
    .QN(_20978_));
 DFFR_X1 \core.keymem.key_mem[1][11]$_DFFE_PN0P_  (.D(_01627_),
    .RN(net95),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[1][11] ),
    .QN(_20977_));
 DFFR_X1 \core.keymem.key_mem[1][120]$_DFFE_PN0P_  (.D(_01628_),
    .RN(net93),
    .CK(clknet_leaf_205_clk),
    .Q(\core.keymem.key_mem[1][120] ),
    .QN(_20976_));
 DFFR_X1 \core.keymem.key_mem[1][121]$_DFFE_PN0P_  (.D(_01629_),
    .RN(net92),
    .CK(clknet_leaf_266_clk),
    .Q(\core.keymem.key_mem[1][121] ),
    .QN(_20975_));
 DFFR_X1 \core.keymem.key_mem[1][122]$_DFFE_PN0P_  (.D(_01630_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[1][122] ),
    .QN(_20974_));
 DFFR_X1 \core.keymem.key_mem[1][123]$_DFFE_PN0P_  (.D(_01631_),
    .RN(net93),
    .CK(clknet_leaf_197_clk),
    .Q(\core.keymem.key_mem[1][123] ),
    .QN(_20973_));
 DFFR_X1 \core.keymem.key_mem[1][124]$_DFFE_PN0P_  (.D(_01632_),
    .RN(net93),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[1][124] ),
    .QN(_20972_));
 DFFR_X2 \core.keymem.key_mem[1][125]$_DFFE_PN0P_  (.D(_01633_),
    .RN(net85),
    .CK(clknet_leaf_53_clk),
    .Q(\core.keymem.key_mem[1][125] ),
    .QN(_20971_));
 DFFR_X1 \core.keymem.key_mem[1][126]$_DFFE_PN0P_  (.D(_01634_),
    .RN(net98),
    .CK(clknet_leaf_166_clk),
    .Q(\core.keymem.key_mem[1][126] ),
    .QN(_20970_));
 DFFR_X1 \core.keymem.key_mem[1][127]$_DFFE_PN0P_  (.D(_01635_),
    .RN(net97),
    .CK(clknet_leaf_241_clk),
    .Q(\core.keymem.key_mem[1][127] ),
    .QN(_20969_));
 DFFR_X1 \core.keymem.key_mem[1][12]$_DFFE_PN0P_  (.D(_01636_),
    .RN(net93),
    .CK(clknet_leaf_191_clk),
    .Q(\core.keymem.key_mem[1][12] ),
    .QN(_20968_));
 DFFR_X2 \core.keymem.key_mem[1][13]$_DFFE_PN0P_  (.D(_01637_),
    .RN(net85),
    .CK(clknet_leaf_52_clk),
    .Q(\core.keymem.key_mem[1][13] ),
    .QN(_20967_));
 DFFR_X2 \core.keymem.key_mem[1][14]$_DFFE_PN0P_  (.D(_01638_),
    .RN(net93),
    .CK(clknet_leaf_377_clk),
    .Q(\core.keymem.key_mem[1][14] ),
    .QN(_20966_));
 DFFR_X1 \core.keymem.key_mem[1][15]$_DFFE_PN0P_  (.D(_01639_),
    .RN(net98),
    .CK(clknet_leaf_229_clk),
    .Q(\core.keymem.key_mem[1][15] ),
    .QN(_20965_));
 DFFR_X1 \core.keymem.key_mem[1][16]$_DFFE_PN0P_  (.D(_01640_),
    .RN(net87),
    .CK(clknet_leaf_31_clk),
    .Q(\core.keymem.key_mem[1][16] ),
    .QN(_20964_));
 DFFR_X1 \core.keymem.key_mem[1][17]$_DFFE_PN0P_  (.D(_01641_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[1][17] ),
    .QN(_20963_));
 DFFR_X1 \core.keymem.key_mem[1][18]$_DFFE_PN0P_  (.D(_01642_),
    .RN(net88),
    .CK(clknet_leaf_28_clk),
    .Q(\core.keymem.key_mem[1][18] ),
    .QN(_20962_));
 DFFR_X1 \core.keymem.key_mem[1][19]$_DFFE_PN0P_  (.D(_01643_),
    .RN(net85),
    .CK(clknet_leaf_54_clk),
    .Q(\core.keymem.key_mem[1][19] ),
    .QN(_20961_));
 DFFR_X1 \core.keymem.key_mem[1][1]$_DFFE_PN0P_  (.D(_01644_),
    .RN(net82),
    .CK(clknet_leaf_10_clk),
    .Q(\core.keymem.key_mem[1][1] ),
    .QN(_20960_));
 DFFR_X1 \core.keymem.key_mem[1][20]$_DFFE_PN0P_  (.D(_01645_),
    .RN(net89),
    .CK(clknet_leaf_96_clk),
    .Q(\core.keymem.key_mem[1][20] ),
    .QN(_20959_));
 DFFR_X1 \core.keymem.key_mem[1][21]$_DFFE_PN0P_  (.D(_01646_),
    .RN(net85),
    .CK(clknet_leaf_51_clk),
    .Q(\core.keymem.key_mem[1][21] ),
    .QN(_20958_));
 DFFR_X1 \core.keymem.key_mem[1][22]$_DFFE_PN0P_  (.D(_01647_),
    .RN(net98),
    .CK(clknet_leaf_228_clk),
    .Q(\core.keymem.key_mem[1][22] ),
    .QN(_20957_));
 DFFR_X1 \core.keymem.key_mem[1][23]$_DFFE_PN0P_  (.D(_01648_),
    .RN(net89),
    .CK(clknet_leaf_55_clk),
    .Q(\core.keymem.key_mem[1][23] ),
    .QN(_20956_));
 DFFR_X1 \core.keymem.key_mem[1][24]$_DFFE_PN0P_  (.D(_01649_),
    .RN(net85),
    .CK(clknet_leaf_43_clk),
    .Q(\core.keymem.key_mem[1][24] ),
    .QN(_20955_));
 DFFR_X1 \core.keymem.key_mem[1][25]$_DFFE_PN0P_  (.D(_01650_),
    .RN(net85),
    .CK(clknet_leaf_51_clk),
    .Q(\core.keymem.key_mem[1][25] ),
    .QN(_20954_));
 DFFR_X1 \core.keymem.key_mem[1][26]$_DFFE_PN0P_  (.D(_01651_),
    .RN(net89),
    .CK(clknet_leaf_92_clk),
    .Q(\core.keymem.key_mem[1][26] ),
    .QN(_20953_));
 DFFR_X1 \core.keymem.key_mem[1][27]$_DFFE_PN0P_  (.D(_01652_),
    .RN(net88),
    .CK(clknet_leaf_46_clk),
    .Q(\core.keymem.key_mem[1][27] ),
    .QN(_20952_));
 DFFR_X2 \core.keymem.key_mem[1][28]$_DFFE_PN0P_  (.D(_01653_),
    .RN(net82),
    .CK(clknet_leaf_13_clk),
    .Q(\core.keymem.key_mem[1][28] ),
    .QN(_20951_));
 DFFR_X2 \core.keymem.key_mem[1][29]$_DFFE_PN0P_  (.D(_01654_),
    .RN(net85),
    .CK(clknet_leaf_50_clk),
    .Q(\core.keymem.key_mem[1][29] ),
    .QN(_20950_));
 DFFR_X1 \core.keymem.key_mem[1][2]$_DFFE_PN0P_  (.D(_01655_),
    .RN(net89),
    .CK(clknet_leaf_66_clk),
    .Q(\core.keymem.key_mem[1][2] ),
    .QN(_20949_));
 DFFR_X2 \core.keymem.key_mem[1][30]$_DFFE_PN0P_  (.D(_01656_),
    .RN(net88),
    .CK(clknet_leaf_46_clk),
    .Q(\core.keymem.key_mem[1][30] ),
    .QN(_20948_));
 DFFR_X1 \core.keymem.key_mem[1][31]$_DFFE_PN0P_  (.D(_01657_),
    .RN(net99),
    .CK(clknet_leaf_80_clk),
    .Q(\core.keymem.key_mem[1][31] ),
    .QN(_20947_));
 DFFR_X1 \core.keymem.key_mem[1][32]$_DFFE_PN0P_  (.D(_01658_),
    .RN(net99),
    .CK(clknet_leaf_116_clk),
    .Q(\core.keymem.key_mem[1][32] ),
    .QN(_20946_));
 DFFR_X2 \core.keymem.key_mem[1][33]$_DFFE_PN0P_  (.D(_01659_),
    .RN(net100),
    .CK(clknet_leaf_115_clk),
    .Q(\core.keymem.key_mem[1][33] ),
    .QN(_20945_));
 DFFR_X1 \core.keymem.key_mem[1][34]$_DFFE_PN0P_  (.D(_01660_),
    .RN(net99),
    .CK(clknet_leaf_122_clk),
    .Q(\core.keymem.key_mem[1][34] ),
    .QN(_20944_));
 DFFR_X1 \core.keymem.key_mem[1][35]$_DFFE_PN0P_  (.D(_01661_),
    .RN(net88),
    .CK(clknet_leaf_83_clk),
    .Q(\core.keymem.key_mem[1][35] ),
    .QN(_20943_));
 DFFR_X1 \core.keymem.key_mem[1][36]$_DFFE_PN0P_  (.D(_01662_),
    .RN(net87),
    .CK(clknet_leaf_28_clk),
    .Q(\core.keymem.key_mem[1][36] ),
    .QN(_20942_));
 DFFR_X1 \core.keymem.key_mem[1][37]$_DFFE_PN0P_  (.D(_01663_),
    .RN(net88),
    .CK(clknet_leaf_93_clk),
    .Q(\core.keymem.key_mem[1][37] ),
    .QN(_20941_));
 DFFR_X2 \core.keymem.key_mem[1][38]$_DFFE_PN0P_  (.D(_01664_),
    .RN(net88),
    .CK(clknet_leaf_28_clk),
    .Q(\core.keymem.key_mem[1][38] ),
    .QN(_20940_));
 DFFR_X1 \core.keymem.key_mem[1][39]$_DFFE_PN0P_  (.D(_01665_),
    .RN(net85),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[1][39] ),
    .QN(_20939_));
 DFFR_X1 \core.keymem.key_mem[1][3]$_DFFE_PN0P_  (.D(_01666_),
    .RN(net89),
    .CK(clknet_leaf_91_clk),
    .Q(\core.keymem.key_mem[1][3] ),
    .QN(_20938_));
 DFFR_X1 \core.keymem.key_mem[1][40]$_DFFE_PN0P_  (.D(_01667_),
    .RN(net85),
    .CK(clknet_leaf_89_clk),
    .Q(\core.keymem.key_mem[1][40] ),
    .QN(_20937_));
 DFFR_X1 \core.keymem.key_mem[1][41]$_DFFE_PN0P_  (.D(_01668_),
    .RN(net89),
    .CK(clknet_leaf_83_clk),
    .Q(\core.keymem.key_mem[1][41] ),
    .QN(_20936_));
 DFFR_X1 \core.keymem.key_mem[1][42]$_DFFE_PN0P_  (.D(_01669_),
    .RN(net99),
    .CK(clknet_leaf_117_clk),
    .Q(\core.keymem.key_mem[1][42] ),
    .QN(_20935_));
 DFFR_X1 \core.keymem.key_mem[1][43]$_DFFE_PN0P_  (.D(_01670_),
    .RN(net85),
    .CK(clknet_leaf_88_clk),
    .Q(\core.keymem.key_mem[1][43] ),
    .QN(_20934_));
 DFFR_X1 \core.keymem.key_mem[1][44]$_DFFE_PN0P_  (.D(_01671_),
    .RN(net99),
    .CK(clknet_leaf_115_clk),
    .Q(\core.keymem.key_mem[1][44] ),
    .QN(_20933_));
 DFFR_X1 \core.keymem.key_mem[1][45]$_DFFE_PN0P_  (.D(_01672_),
    .RN(net99),
    .CK(clknet_leaf_69_clk),
    .Q(\core.keymem.key_mem[1][45] ),
    .QN(_20932_));
 DFFR_X1 \core.keymem.key_mem[1][46]$_DFFE_PN0P_  (.D(_01673_),
    .RN(net89),
    .CK(clknet_leaf_84_clk),
    .Q(\core.keymem.key_mem[1][46] ),
    .QN(_20931_));
 DFFR_X1 \core.keymem.key_mem[1][47]$_DFFE_PN0P_  (.D(_01674_),
    .RN(net98),
    .CK(clknet_leaf_146_clk),
    .Q(\core.keymem.key_mem[1][47] ),
    .QN(_20930_));
 DFFR_X1 \core.keymem.key_mem[1][48]$_DFFE_PN0P_  (.D(_01675_),
    .RN(net95),
    .CK(clknet_leaf_121_clk),
    .Q(\core.keymem.key_mem[1][48] ),
    .QN(_20929_));
 DFFR_X1 \core.keymem.key_mem[1][49]$_DFFE_PN0P_  (.D(_01676_),
    .RN(net99),
    .CK(clknet_leaf_82_clk),
    .Q(\core.keymem.key_mem[1][49] ),
    .QN(_20928_));
 DFFR_X1 \core.keymem.key_mem[1][4]$_DFFE_PN0P_  (.D(_01677_),
    .RN(net88),
    .CK(clknet_leaf_92_clk),
    .Q(\core.keymem.key_mem[1][4] ),
    .QN(_20927_));
 DFFR_X1 \core.keymem.key_mem[1][50]$_DFFE_PN0P_  (.D(_01678_),
    .RN(net98),
    .CK(clknet_leaf_139_clk),
    .Q(\core.keymem.key_mem[1][50] ),
    .QN(_20926_));
 DFFR_X1 \core.keymem.key_mem[1][51]$_DFFE_PN0P_  (.D(_01679_),
    .RN(net99),
    .CK(clknet_leaf_121_clk),
    .Q(\core.keymem.key_mem[1][51] ),
    .QN(_20925_));
 DFFR_X1 \core.keymem.key_mem[1][52]$_DFFE_PN0P_  (.D(_01680_),
    .RN(net89),
    .CK(clknet_leaf_83_clk),
    .Q(\core.keymem.key_mem[1][52] ),
    .QN(_20924_));
 DFFR_X1 \core.keymem.key_mem[1][53]$_DFFE_PN0P_  (.D(_01681_),
    .RN(net97),
    .CK(clknet_leaf_144_clk),
    .Q(\core.keymem.key_mem[1][53] ),
    .QN(_20923_));
 DFFR_X1 \core.keymem.key_mem[1][54]$_DFFE_PN0P_  (.D(_01682_),
    .RN(net98),
    .CK(clknet_leaf_142_clk),
    .Q(\core.keymem.key_mem[1][54] ),
    .QN(_20922_));
 DFFR_X1 \core.keymem.key_mem[1][55]$_DFFE_PN0P_  (.D(_01683_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[1][55] ),
    .QN(_20921_));
 DFFR_X2 \core.keymem.key_mem[1][56]$_DFFE_PN0P_  (.D(_01684_),
    .RN(net88),
    .CK(clknet_leaf_44_clk),
    .Q(\core.keymem.key_mem[1][56] ),
    .QN(_20920_));
 DFFR_X1 \core.keymem.key_mem[1][57]$_DFFE_PN0P_  (.D(_01685_),
    .RN(net100),
    .CK(clknet_leaf_108_clk),
    .Q(\core.keymem.key_mem[1][57] ),
    .QN(_20919_));
 DFFR_X1 \core.keymem.key_mem[1][58]$_DFFE_PN0P_  (.D(_01686_),
    .RN(net100),
    .CK(clknet_leaf_103_clk),
    .Q(\core.keymem.key_mem[1][58] ),
    .QN(_20918_));
 DFFR_X1 \core.keymem.key_mem[1][59]$_DFFE_PN0P_  (.D(_01687_),
    .RN(net89),
    .CK(clknet_leaf_27_clk),
    .Q(\core.keymem.key_mem[1][59] ),
    .QN(_20917_));
 DFFR_X1 \core.keymem.key_mem[1][5]$_DFFE_PN0P_  (.D(_01688_),
    .RN(net100),
    .CK(clknet_leaf_20_clk),
    .Q(\core.keymem.key_mem[1][5] ),
    .QN(_20916_));
 DFFR_X1 \core.keymem.key_mem[1][60]$_DFFE_PN0P_  (.D(_01689_),
    .RN(net87),
    .CK(clknet_leaf_31_clk),
    .Q(\core.keymem.key_mem[1][60] ),
    .QN(_20915_));
 DFFR_X1 \core.keymem.key_mem[1][61]$_DFFE_PN0P_  (.D(_01690_),
    .RN(net89),
    .CK(clknet_leaf_84_clk),
    .Q(\core.keymem.key_mem[1][61] ),
    .QN(_20914_));
 DFFR_X1 \core.keymem.key_mem[1][62]$_DFFE_PN0P_  (.D(_01691_),
    .RN(net89),
    .CK(clknet_leaf_27_clk),
    .Q(\core.keymem.key_mem[1][62] ),
    .QN(_20913_));
 DFFR_X1 \core.keymem.key_mem[1][63]$_DFFE_PN0P_  (.D(_01692_),
    .RN(net100),
    .CK(clknet_leaf_21_clk),
    .Q(\core.keymem.key_mem[1][63] ),
    .QN(_20912_));
 DFFR_X1 \core.keymem.key_mem[1][64]$_DFFE_PN0P_  (.D(_01693_),
    .RN(net82),
    .CK(clknet_leaf_15_clk),
    .Q(\core.keymem.key_mem[1][64] ),
    .QN(_20911_));
 DFFR_X1 \core.keymem.key_mem[1][65]$_DFFE_PN0P_  (.D(_01694_),
    .RN(net99),
    .CK(clknet_leaf_121_clk),
    .Q(\core.keymem.key_mem[1][65] ),
    .QN(_20910_));
 DFFR_X2 \core.keymem.key_mem[1][66]$_DFFE_PN0P_  (.D(_01695_),
    .RN(net82),
    .CK(clknet_leaf_35_clk),
    .Q(\core.keymem.key_mem[1][66] ),
    .QN(_20909_));
 DFFR_X1 \core.keymem.key_mem[1][67]$_DFFE_PN0P_  (.D(_01696_),
    .RN(net99),
    .CK(clknet_leaf_74_clk),
    .Q(\core.keymem.key_mem[1][67] ),
    .QN(_20908_));
 DFFR_X1 \core.keymem.key_mem[1][68]$_DFFE_PN0P_  (.D(_01697_),
    .RN(net99),
    .CK(clknet_leaf_116_clk),
    .Q(\core.keymem.key_mem[1][68] ),
    .QN(_20907_));
 DFFR_X1 \core.keymem.key_mem[1][69]$_DFFE_PN0P_  (.D(_01698_),
    .RN(net98),
    .CK(clknet_leaf_177_clk),
    .Q(\core.keymem.key_mem[1][69] ),
    .QN(_20906_));
 DFFR_X1 \core.keymem.key_mem[1][6]$_DFFE_PN0P_  (.D(_01699_),
    .RN(net100),
    .CK(clknet_leaf_103_clk),
    .Q(\core.keymem.key_mem[1][6] ),
    .QN(_20905_));
 DFFR_X1 \core.keymem.key_mem[1][70]$_DFFE_PN0P_  (.D(_01700_),
    .RN(net88),
    .CK(clknet_leaf_92_clk),
    .Q(\core.keymem.key_mem[1][70] ),
    .QN(_20904_));
 DFFR_X1 \core.keymem.key_mem[1][71]$_DFFE_PN0P_  (.D(_01701_),
    .RN(net99),
    .CK(clknet_leaf_71_clk),
    .Q(\core.keymem.key_mem[1][71] ),
    .QN(_20903_));
 DFFR_X1 \core.keymem.key_mem[1][72]$_DFFE_PN0P_  (.D(_01702_),
    .RN(net95),
    .CK(clknet_leaf_76_clk),
    .Q(\core.keymem.key_mem[1][72] ),
    .QN(_20902_));
 DFFR_X1 \core.keymem.key_mem[1][73]$_DFFE_PN0P_  (.D(_01703_),
    .RN(net97),
    .CK(clknet_leaf_146_clk),
    .Q(\core.keymem.key_mem[1][73] ),
    .QN(_20901_));
 DFFR_X1 \core.keymem.key_mem[1][74]$_DFFE_PN0P_  (.D(_01704_),
    .RN(net97),
    .CK(clknet_leaf_164_clk),
    .Q(\core.keymem.key_mem[1][74] ),
    .QN(_20900_));
 DFFR_X1 \core.keymem.key_mem[1][75]$_DFFE_PN0P_  (.D(_01705_),
    .RN(net97),
    .CK(clknet_leaf_148_clk),
    .Q(\core.keymem.key_mem[1][75] ),
    .QN(_20899_));
 DFFR_X1 \core.keymem.key_mem[1][76]$_DFFE_PN0P_  (.D(_01706_),
    .RN(net93),
    .CK(clknet_leaf_283_clk),
    .Q(\core.keymem.key_mem[1][76] ),
    .QN(_20898_));
 DFFR_X1 \core.keymem.key_mem[1][77]$_DFFE_PN0P_  (.D(_01707_),
    .RN(net97),
    .CK(clknet_leaf_164_clk),
    .Q(\core.keymem.key_mem[1][77] ),
    .QN(_20897_));
 DFFR_X1 \core.keymem.key_mem[1][78]$_DFFE_PN0P_  (.D(_01708_),
    .RN(net96),
    .CK(clknet_leaf_171_clk),
    .Q(\core.keymem.key_mem[1][78] ),
    .QN(_20896_));
 DFFR_X1 \core.keymem.key_mem[1][79]$_DFFE_PN0P_  (.D(_01709_),
    .RN(net98),
    .CK(clknet_leaf_228_clk),
    .Q(\core.keymem.key_mem[1][79] ),
    .QN(_20895_));
 DFFR_X1 \core.keymem.key_mem[1][7]$_DFFE_PN0P_  (.D(_01710_),
    .RN(net98),
    .CK(clknet_leaf_172_clk),
    .Q(\core.keymem.key_mem[1][7] ),
    .QN(_20894_));
 DFFR_X1 \core.keymem.key_mem[1][80]$_DFFE_PN0P_  (.D(_01711_),
    .RN(net97),
    .CK(clknet_leaf_163_clk),
    .Q(\core.keymem.key_mem[1][80] ),
    .QN(_20893_));
 DFFR_X1 \core.keymem.key_mem[1][81]$_DFFE_PN0P_  (.D(_01712_),
    .RN(net97),
    .CK(clknet_leaf_155_clk),
    .Q(\core.keymem.key_mem[1][81] ),
    .QN(_20892_));
 DFFR_X1 \core.keymem.key_mem[1][82]$_DFFE_PN0P_  (.D(_01713_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[1][82] ),
    .QN(_20891_));
 DFFR_X1 \core.keymem.key_mem[1][83]$_DFFE_PN0P_  (.D(_01714_),
    .RN(net93),
    .CK(clknet_leaf_183_clk),
    .Q(\core.keymem.key_mem[1][83] ),
    .QN(_20890_));
 DFFR_X1 \core.keymem.key_mem[1][84]$_DFFE_PN0P_  (.D(_01715_),
    .RN(net94),
    .CK(clknet_leaf_181_clk),
    .Q(\core.keymem.key_mem[1][84] ),
    .QN(_20889_));
 DFFR_X1 \core.keymem.key_mem[1][85]$_DFFE_PN0P_  (.D(_01716_),
    .RN(net96),
    .CK(clknet_leaf_230_clk),
    .Q(\core.keymem.key_mem[1][85] ),
    .QN(_20888_));
 DFFR_X1 \core.keymem.key_mem[1][86]$_DFFE_PN0P_  (.D(_01717_),
    .RN(net98),
    .CK(clknet_leaf_166_clk),
    .Q(\core.keymem.key_mem[1][86] ),
    .QN(_20887_));
 DFFR_X1 \core.keymem.key_mem[1][87]$_DFFE_PN0P_  (.D(_01718_),
    .RN(net89),
    .CK(clknet_leaf_378_clk),
    .Q(\core.keymem.key_mem[1][87] ),
    .QN(_20886_));
 DFFR_X1 \core.keymem.key_mem[1][88]$_DFFE_PN0P_  (.D(_01719_),
    .RN(net93),
    .CK(clknet_leaf_282_clk),
    .Q(\core.keymem.key_mem[1][88] ),
    .QN(_20885_));
 DFFR_X1 \core.keymem.key_mem[1][89]$_DFFE_PN0P_  (.D(_01720_),
    .RN(net93),
    .CK(clknet_leaf_199_clk),
    .Q(\core.keymem.key_mem[1][89] ),
    .QN(_20884_));
 DFFR_X1 \core.keymem.key_mem[1][8]$_DFFE_PN0P_  (.D(_01721_),
    .RN(net89),
    .CK(clknet_leaf_57_clk),
    .Q(\core.keymem.key_mem[1][8] ),
    .QN(_20883_));
 DFFR_X1 \core.keymem.key_mem[1][90]$_DFFE_PN0P_  (.D(_01722_),
    .RN(net97),
    .CK(clknet_leaf_163_clk),
    .Q(\core.keymem.key_mem[1][90] ),
    .QN(_20882_));
 DFFR_X1 \core.keymem.key_mem[1][91]$_DFFE_PN0P_  (.D(_01723_),
    .RN(net93),
    .CK(clknet_leaf_184_clk),
    .Q(\core.keymem.key_mem[1][91] ),
    .QN(_20881_));
 DFFR_X1 \core.keymem.key_mem[1][92]$_DFFE_PN0P_  (.D(_01724_),
    .RN(net95),
    .CK(clknet_leaf_62_clk),
    .Q(\core.keymem.key_mem[1][92] ),
    .QN(_20880_));
 DFFR_X1 \core.keymem.key_mem[1][93]$_DFFE_PN0P_  (.D(_01725_),
    .RN(net95),
    .CK(clknet_leaf_190_clk),
    .Q(\core.keymem.key_mem[1][93] ),
    .QN(_20879_));
 DFFR_X1 \core.keymem.key_mem[1][94]$_DFFE_PN0P_  (.D(_01726_),
    .RN(net94),
    .CK(clknet_leaf_214_clk),
    .Q(\core.keymem.key_mem[1][94] ),
    .QN(_20878_));
 DFFR_X1 \core.keymem.key_mem[1][95]$_DFFE_PN0P_  (.D(_01727_),
    .RN(net96),
    .CK(clknet_leaf_234_clk),
    .Q(\core.keymem.key_mem[1][95] ),
    .QN(_20877_));
 DFFR_X1 \core.keymem.key_mem[1][96]$_DFFE_PN0P_  (.D(_01728_),
    .RN(net89),
    .CK(clknet_leaf_374_clk),
    .Q(\core.keymem.key_mem[1][96] ),
    .QN(_20876_));
 DFFR_X1 \core.keymem.key_mem[1][97]$_DFFE_PN0P_  (.D(_01729_),
    .RN(net95),
    .CK(clknet_leaf_194_clk),
    .Q(\core.keymem.key_mem[1][97] ),
    .QN(_20875_));
 DFFR_X1 \core.keymem.key_mem[1][98]$_DFFE_PN0P_  (.D(_01730_),
    .RN(net89),
    .CK(clknet_leaf_59_clk),
    .Q(\core.keymem.key_mem[1][98] ),
    .QN(_20874_));
 DFFR_X1 \core.keymem.key_mem[1][99]$_DFFE_PN0P_  (.D(_01731_),
    .RN(net93),
    .CK(clknet_leaf_201_clk),
    .Q(\core.keymem.key_mem[1][99] ),
    .QN(_20873_));
 DFFR_X1 \core.keymem.key_mem[1][9]$_DFFE_PN0P_  (.D(_01732_),
    .RN(net91),
    .CK(clknet_leaf_200_clk),
    .Q(\core.keymem.key_mem[1][9] ),
    .QN(_20872_));
 DFFR_X1 \core.keymem.key_mem[2][0]$_DFFE_PN0P_  (.D(_01733_),
    .RN(net96),
    .CK(clknet_leaf_248_clk),
    .Q(\core.keymem.key_mem[2][0] ),
    .QN(_20871_));
 DFFR_X1 \core.keymem.key_mem[2][100]$_DFFE_PN0P_  (.D(_01734_),
    .RN(net94),
    .CK(clknet_leaf_210_clk),
    .Q(\core.keymem.key_mem[2][100] ),
    .QN(_20870_));
 DFFR_X1 \core.keymem.key_mem[2][101]$_DFFE_PN0P_  (.D(_01735_),
    .RN(net94),
    .CK(clknet_leaf_212_clk),
    .Q(\core.keymem.key_mem[2][101] ),
    .QN(_20869_));
 DFFR_X1 \core.keymem.key_mem[2][102]$_DFFE_PN0P_  (.D(_01736_),
    .RN(net96),
    .CK(clknet_leaf_233_clk),
    .Q(\core.keymem.key_mem[2][102] ),
    .QN(_20868_));
 DFFR_X1 \core.keymem.key_mem[2][103]$_DFFE_PN0P_  (.D(_01737_),
    .RN(net96),
    .CK(clknet_leaf_246_clk),
    .Q(\core.keymem.key_mem[2][103] ),
    .QN(_20867_));
 DFFR_X1 \core.keymem.key_mem[2][104]$_DFFE_PN0P_  (.D(_01738_),
    .RN(net93),
    .CK(clknet_leaf_191_clk),
    .Q(\core.keymem.key_mem[2][104] ),
    .QN(_20866_));
 DFFR_X1 \core.keymem.key_mem[2][105]$_DFFE_PN0P_  (.D(_01739_),
    .RN(net96),
    .CK(clknet_leaf_247_clk),
    .Q(\core.keymem.key_mem[2][105] ),
    .QN(_20865_));
 DFFR_X1 \core.keymem.key_mem[2][106]$_DFFE_PN0P_  (.D(_01740_),
    .RN(net92),
    .CK(clknet_leaf_268_clk),
    .Q(\core.keymem.key_mem[2][106] ),
    .QN(_20864_));
 DFFR_X1 \core.keymem.key_mem[2][107]$_DFFE_PN0P_  (.D(_01741_),
    .RN(net92),
    .CK(clknet_leaf_269_clk),
    .Q(\core.keymem.key_mem[2][107] ),
    .QN(_20863_));
 DFFR_X1 \core.keymem.key_mem[2][108]$_DFFE_PN0P_  (.D(_01742_),
    .RN(net91),
    .CK(clknet_leaf_203_clk),
    .Q(\core.keymem.key_mem[2][108] ),
    .QN(_20862_));
 DFFR_X1 \core.keymem.key_mem[2][109]$_DFFE_PN0P_  (.D(_01743_),
    .RN(net94),
    .CK(clknet_leaf_263_clk),
    .Q(\core.keymem.key_mem[2][109] ),
    .QN(_20861_));
 DFFR_X1 \core.keymem.key_mem[2][10]$_DFFE_PN0P_  (.D(_01744_),
    .RN(net95),
    .CK(clknet_leaf_189_clk),
    .Q(\core.keymem.key_mem[2][10] ),
    .QN(_20860_));
 DFFR_X1 \core.keymem.key_mem[2][110]$_DFFE_PN0P_  (.D(_01745_),
    .RN(net96),
    .CK(clknet_leaf_249_clk),
    .Q(\core.keymem.key_mem[2][110] ),
    .QN(_20859_));
 DFFR_X1 \core.keymem.key_mem[2][111]$_DFFE_PN0P_  (.D(_01746_),
    .RN(net96),
    .CK(clknet_leaf_225_clk),
    .Q(\core.keymem.key_mem[2][111] ),
    .QN(_20858_));
 DFFR_X1 \core.keymem.key_mem[2][112]$_DFFE_PN0P_  (.D(_01747_),
    .RN(net94),
    .CK(clknet_leaf_262_clk),
    .Q(\core.keymem.key_mem[2][112] ),
    .QN(_20857_));
 DFFR_X1 \core.keymem.key_mem[2][113]$_DFFE_PN0P_  (.D(_01748_),
    .RN(net91),
    .CK(clknet_leaf_280_clk),
    .Q(\core.keymem.key_mem[2][113] ),
    .QN(_20856_));
 DFFR_X1 \core.keymem.key_mem[2][114]$_DFFE_PN0P_  (.D(_01749_),
    .RN(net91),
    .CK(clknet_leaf_278_clk),
    .Q(\core.keymem.key_mem[2][114] ),
    .QN(_20855_));
 DFFR_X1 \core.keymem.key_mem[2][115]$_DFFE_PN0P_  (.D(_01750_),
    .RN(net92),
    .CK(clknet_leaf_275_clk),
    .Q(\core.keymem.key_mem[2][115] ),
    .QN(_20854_));
 DFFR_X1 \core.keymem.key_mem[2][116]$_DFFE_PN0P_  (.D(_01751_),
    .RN(net94),
    .CK(clknet_leaf_262_clk),
    .Q(\core.keymem.key_mem[2][116] ),
    .QN(_20853_));
 DFFR_X1 \core.keymem.key_mem[2][117]$_DFFE_PN0P_  (.D(_01752_),
    .RN(net94),
    .CK(clknet_leaf_212_clk),
    .Q(\core.keymem.key_mem[2][117] ),
    .QN(_20852_));
 DFFR_X1 \core.keymem.key_mem[2][118]$_DFFE_PN0P_  (.D(_01753_),
    .RN(net98),
    .CK(clknet_leaf_227_clk),
    .Q(\core.keymem.key_mem[2][118] ),
    .QN(_20851_));
 DFFR_X1 \core.keymem.key_mem[2][119]$_DFFE_PN0P_  (.D(_01754_),
    .RN(net94),
    .CK(clknet_leaf_262_clk),
    .Q(\core.keymem.key_mem[2][119] ),
    .QN(_20850_));
 DFFR_X1 \core.keymem.key_mem[2][11]$_DFFE_PN0P_  (.D(_01755_),
    .RN(net95),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[2][11] ),
    .QN(_20849_));
 DFFR_X1 \core.keymem.key_mem[2][120]$_DFFE_PN0P_  (.D(_01756_),
    .RN(net94),
    .CK(clknet_leaf_215_clk),
    .Q(\core.keymem.key_mem[2][120] ),
    .QN(_20848_));
 DFFR_X1 \core.keymem.key_mem[2][121]$_DFFE_PN0P_  (.D(_01757_),
    .RN(net94),
    .CK(clknet_leaf_268_clk),
    .Q(\core.keymem.key_mem[2][121] ),
    .QN(_20847_));
 DFFR_X1 \core.keymem.key_mem[2][122]$_DFFE_PN0P_  (.D(_01758_),
    .RN(net97),
    .CK(clknet_leaf_237_clk),
    .Q(\core.keymem.key_mem[2][122] ),
    .QN(_20846_));
 DFFR_X1 \core.keymem.key_mem[2][123]$_DFFE_PN0P_  (.D(_01759_),
    .RN(net93),
    .CK(clknet_leaf_198_clk),
    .Q(\core.keymem.key_mem[2][123] ),
    .QN(_20845_));
 DFFR_X1 \core.keymem.key_mem[2][124]$_DFFE_PN0P_  (.D(_01760_),
    .RN(net93),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[2][124] ),
    .QN(_20844_));
 DFFR_X1 \core.keymem.key_mem[2][125]$_DFFE_PN0P_  (.D(_01761_),
    .RN(net97),
    .CK(clknet_leaf_234_clk),
    .Q(\core.keymem.key_mem[2][125] ),
    .QN(_20843_));
 DFFR_X1 \core.keymem.key_mem[2][126]$_DFFE_PN0P_  (.D(_01762_),
    .RN(net98),
    .CK(clknet_leaf_166_clk),
    .Q(\core.keymem.key_mem[2][126] ),
    .QN(_20842_));
 DFFR_X1 \core.keymem.key_mem[2][127]$_DFFE_PN0P_  (.D(_01763_),
    .RN(net97),
    .CK(clknet_leaf_240_clk),
    .Q(\core.keymem.key_mem[2][127] ),
    .QN(_20841_));
 DFFR_X1 \core.keymem.key_mem[2][12]$_DFFE_PN0P_  (.D(_01764_),
    .RN(net93),
    .CK(clknet_leaf_207_clk),
    .Q(\core.keymem.key_mem[2][12] ),
    .QN(_20840_));
 DFFR_X1 \core.keymem.key_mem[2][13]$_DFFE_PN0P_  (.D(_01765_),
    .RN(net85),
    .CK(clknet_leaf_53_clk),
    .Q(\core.keymem.key_mem[2][13] ),
    .QN(_20839_));
 DFFR_X1 \core.keymem.key_mem[2][14]$_DFFE_PN0P_  (.D(_01766_),
    .RN(net89),
    .CK(clknet_leaf_379_clk),
    .Q(\core.keymem.key_mem[2][14] ),
    .QN(_20838_));
 DFFR_X1 \core.keymem.key_mem[2][15]$_DFFE_PN0P_  (.D(_01767_),
    .RN(net96),
    .CK(clknet_leaf_230_clk),
    .Q(\core.keymem.key_mem[2][15] ),
    .QN(_20837_));
 DFFR_X1 \core.keymem.key_mem[2][16]$_DFFE_PN0P_  (.D(_01768_),
    .RN(net87),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[2][16] ),
    .QN(_20836_));
 DFFR_X1 \core.keymem.key_mem[2][17]$_DFFE_PN0P_  (.D(_01769_),
    .RN(net98),
    .CK(clknet_leaf_168_clk),
    .Q(\core.keymem.key_mem[2][17] ),
    .QN(_20835_));
 DFFR_X1 \core.keymem.key_mem[2][18]$_DFFE_PN0P_  (.D(_01770_),
    .RN(net82),
    .CK(clknet_leaf_34_clk),
    .Q(\core.keymem.key_mem[2][18] ),
    .QN(_20834_));
 DFFR_X1 \core.keymem.key_mem[2][19]$_DFFE_PN0P_  (.D(_01771_),
    .RN(net85),
    .CK(clknet_leaf_54_clk),
    .Q(\core.keymem.key_mem[2][19] ),
    .QN(_20833_));
 DFFR_X1 \core.keymem.key_mem[2][1]$_DFFE_PN0P_  (.D(_01772_),
    .RN(net82),
    .CK(clknet_leaf_13_clk),
    .Q(\core.keymem.key_mem[2][1] ),
    .QN(_20832_));
 DFFR_X1 \core.keymem.key_mem[2][20]$_DFFE_PN0P_  (.D(_01773_),
    .RN(net89),
    .CK(clknet_leaf_92_clk),
    .Q(\core.keymem.key_mem[2][20] ),
    .QN(_20831_));
 DFFR_X1 \core.keymem.key_mem[2][21]$_DFFE_PN0P_  (.D(_01774_),
    .RN(net85),
    .CK(clknet_leaf_65_clk),
    .Q(\core.keymem.key_mem[2][21] ),
    .QN(_20830_));
 DFFR_X1 \core.keymem.key_mem[2][22]$_DFFE_PN0P_  (.D(_01775_),
    .RN(net94),
    .CK(clknet_leaf_219_clk),
    .Q(\core.keymem.key_mem[2][22] ),
    .QN(_20829_));
 DFFR_X1 \core.keymem.key_mem[2][23]$_DFFE_PN0P_  (.D(_01776_),
    .RN(net89),
    .CK(clknet_leaf_56_clk),
    .Q(\core.keymem.key_mem[2][23] ),
    .QN(_20828_));
 DFFR_X1 \core.keymem.key_mem[2][24]$_DFFE_PN0P_  (.D(_01777_),
    .RN(net85),
    .CK(clknet_leaf_65_clk),
    .Q(\core.keymem.key_mem[2][24] ),
    .QN(_20827_));
 DFFR_X1 \core.keymem.key_mem[2][25]$_DFFE_PN0P_  (.D(_01778_),
    .RN(net85),
    .CK(clknet_leaf_47_clk),
    .Q(\core.keymem.key_mem[2][25] ),
    .QN(_20826_));
 DFFR_X1 \core.keymem.key_mem[2][26]$_DFFE_PN0P_  (.D(_01779_),
    .RN(net100),
    .CK(clknet_leaf_96_clk),
    .Q(\core.keymem.key_mem[2][26] ),
    .QN(_20825_));
 DFFR_X1 \core.keymem.key_mem[2][27]$_DFFE_PN0P_  (.D(_01780_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[2][27] ),
    .QN(_20824_));
 DFFR_X1 \core.keymem.key_mem[2][28]$_DFFE_PN0P_  (.D(_01781_),
    .RN(net16),
    .CK(clknet_leaf_125_clk),
    .Q(\core.keymem.key_mem[2][28] ),
    .QN(_20823_));
 DFFR_X1 \core.keymem.key_mem[2][29]$_DFFE_PN0P_  (.D(_01782_),
    .RN(net16),
    .CK(clknet_leaf_132_clk),
    .Q(\core.keymem.key_mem[2][29] ),
    .QN(_20822_));
 DFFR_X1 \core.keymem.key_mem[2][2]$_DFFE_PN0P_  (.D(_01783_),
    .RN(net89),
    .CK(clknet_leaf_66_clk),
    .Q(\core.keymem.key_mem[2][2] ),
    .QN(_20821_));
 DFFR_X1 \core.keymem.key_mem[2][30]$_DFFE_PN0P_  (.D(_01784_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[2][30] ),
    .QN(_20820_));
 DFFR_X1 \core.keymem.key_mem[2][31]$_DFFE_PN0P_  (.D(_01785_),
    .RN(net98),
    .CK(clknet_leaf_144_clk),
    .Q(\core.keymem.key_mem[2][31] ),
    .QN(_20819_));
 DFFR_X1 \core.keymem.key_mem[2][32]$_DFFE_PN0P_  (.D(_01786_),
    .RN(net100),
    .CK(clknet_leaf_111_clk),
    .Q(\core.keymem.key_mem[2][32] ),
    .QN(_20818_));
 DFFR_X1 \core.keymem.key_mem[2][33]$_DFFE_PN0P_  (.D(_01787_),
    .RN(net99),
    .CK(clknet_leaf_127_clk),
    .Q(\core.keymem.key_mem[2][33] ),
    .QN(_20817_));
 DFFR_X1 \core.keymem.key_mem[2][34]$_DFFE_PN0P_  (.D(_01788_),
    .RN(net16),
    .CK(clknet_leaf_124_clk),
    .Q(\core.keymem.key_mem[2][34] ),
    .QN(_20816_));
 DFFR_X1 \core.keymem.key_mem[2][35]$_DFFE_PN0P_  (.D(_01789_),
    .RN(net99),
    .CK(clknet_leaf_127_clk),
    .Q(\core.keymem.key_mem[2][35] ),
    .QN(_20815_));
 DFFR_X1 \core.keymem.key_mem[2][36]$_DFFE_PN0P_  (.D(_01790_),
    .RN(net88),
    .CK(clknet_leaf_90_clk),
    .Q(\core.keymem.key_mem[2][36] ),
    .QN(_20814_));
 DFFR_X1 \core.keymem.key_mem[2][37]$_DFFE_PN0P_  (.D(_01791_),
    .RN(net88),
    .CK(clknet_leaf_93_clk),
    .Q(\core.keymem.key_mem[2][37] ),
    .QN(_20813_));
 DFFR_X1 \core.keymem.key_mem[2][38]$_DFFE_PN0P_  (.D(_01792_),
    .RN(net16),
    .CK(clknet_leaf_124_clk),
    .Q(\core.keymem.key_mem[2][38] ),
    .QN(_20812_));
 DFFR_X1 \core.keymem.key_mem[2][39]$_DFFE_PN0P_  (.D(_01793_),
    .RN(net85),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[2][39] ),
    .QN(_20811_));
 DFFR_X1 \core.keymem.key_mem[2][3]$_DFFE_PN0P_  (.D(_01794_),
    .RN(net88),
    .CK(clknet_leaf_92_clk),
    .Q(\core.keymem.key_mem[2][3] ),
    .QN(_20810_));
 DFFR_X1 \core.keymem.key_mem[2][40]$_DFFE_PN0P_  (.D(_01795_),
    .RN(net85),
    .CK(clknet_leaf_89_clk),
    .Q(\core.keymem.key_mem[2][40] ),
    .QN(_20809_));
 DFFR_X1 \core.keymem.key_mem[2][41]$_DFFE_PN0P_  (.D(_01796_),
    .RN(net99),
    .CK(clknet_leaf_115_clk),
    .Q(\core.keymem.key_mem[2][41] ),
    .QN(_20808_));
 DFFR_X1 \core.keymem.key_mem[2][42]$_DFFE_PN0P_  (.D(_01797_),
    .RN(net95),
    .CK(clknet_leaf_122_clk),
    .Q(\core.keymem.key_mem[2][42] ),
    .QN(_20807_));
 DFFR_X1 \core.keymem.key_mem[2][43]$_DFFE_PN0P_  (.D(_01798_),
    .RN(net85),
    .CK(clknet_leaf_67_clk),
    .Q(\core.keymem.key_mem[2][43] ),
    .QN(_20806_));
 DFFR_X1 \core.keymem.key_mem[2][44]$_DFFE_PN0P_  (.D(_01799_),
    .RN(net100),
    .CK(clknet_leaf_113_clk),
    .Q(\core.keymem.key_mem[2][44] ),
    .QN(_20805_));
 DFFR_X1 \core.keymem.key_mem[2][45]$_DFFE_PN0P_  (.D(_01800_),
    .RN(net99),
    .CK(clknet_leaf_71_clk),
    .Q(\core.keymem.key_mem[2][45] ),
    .QN(_20804_));
 DFFR_X1 \core.keymem.key_mem[2][46]$_DFFE_PN0P_  (.D(_01801_),
    .RN(net99),
    .CK(clknet_leaf_85_clk),
    .Q(\core.keymem.key_mem[2][46] ),
    .QN(_20803_));
 DFFR_X1 \core.keymem.key_mem[2][47]$_DFFE_PN0P_  (.D(_01802_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[2][47] ),
    .QN(_20802_));
 DFFR_X1 \core.keymem.key_mem[2][48]$_DFFE_PN0P_  (.D(_01803_),
    .RN(net98),
    .CK(clknet_leaf_141_clk),
    .Q(\core.keymem.key_mem[2][48] ),
    .QN(_20801_));
 DFFR_X1 \core.keymem.key_mem[2][49]$_DFFE_PN0P_  (.D(_01804_),
    .RN(net99),
    .CK(clknet_leaf_116_clk),
    .Q(\core.keymem.key_mem[2][49] ),
    .QN(_20800_));
 DFFR_X1 \core.keymem.key_mem[2][4]$_DFFE_PN0P_  (.D(_01805_),
    .RN(net100),
    .CK(clknet_leaf_104_clk),
    .Q(\core.keymem.key_mem[2][4] ),
    .QN(_20799_));
 DFFR_X1 \core.keymem.key_mem[2][50]$_DFFE_PN0P_  (.D(_01806_),
    .RN(net98),
    .CK(clknet_leaf_141_clk),
    .Q(\core.keymem.key_mem[2][50] ),
    .QN(_20798_));
 DFFR_X1 \core.keymem.key_mem[2][51]$_DFFE_PN0P_  (.D(_01807_),
    .RN(net100),
    .CK(clknet_leaf_128_clk),
    .Q(\core.keymem.key_mem[2][51] ),
    .QN(_20797_));
 DFFR_X1 \core.keymem.key_mem[2][52]$_DFFE_PN0P_  (.D(_01808_),
    .RN(net99),
    .CK(clknet_leaf_80_clk),
    .Q(\core.keymem.key_mem[2][52] ),
    .QN(_20796_));
 DFFR_X1 \core.keymem.key_mem[2][53]$_DFFE_PN0P_  (.D(_01809_),
    .RN(net97),
    .CK(clknet_leaf_144_clk),
    .Q(\core.keymem.key_mem[2][53] ),
    .QN(_20795_));
 DFFR_X1 \core.keymem.key_mem[2][54]$_DFFE_PN0P_  (.D(_01810_),
    .RN(net98),
    .CK(clknet_leaf_142_clk),
    .Q(\core.keymem.key_mem[2][54] ),
    .QN(_20794_));
 DFFR_X1 \core.keymem.key_mem[2][55]$_DFFE_PN0P_  (.D(_01811_),
    .RN(net16),
    .CK(clknet_leaf_137_clk),
    .Q(\core.keymem.key_mem[2][55] ),
    .QN(_20793_));
 DFFR_X1 \core.keymem.key_mem[2][56]$_DFFE_PN0P_  (.D(_01812_),
    .RN(net97),
    .CK(clknet_leaf_144_clk),
    .Q(\core.keymem.key_mem[2][56] ),
    .QN(_20792_));
 DFFR_X1 \core.keymem.key_mem[2][57]$_DFFE_PN0P_  (.D(_01813_),
    .RN(net100),
    .CK(clknet_leaf_109_clk),
    .Q(\core.keymem.key_mem[2][57] ),
    .QN(_20791_));
 DFFR_X1 \core.keymem.key_mem[2][58]$_DFFE_PN0P_  (.D(_01814_),
    .RN(net100),
    .CK(clknet_leaf_103_clk),
    .Q(\core.keymem.key_mem[2][58] ),
    .QN(_20790_));
 DFFR_X1 \core.keymem.key_mem[2][59]$_DFFE_PN0P_  (.D(_01815_),
    .RN(net89),
    .CK(clknet_leaf_25_clk),
    .Q(\core.keymem.key_mem[2][59] ),
    .QN(_20789_));
 DFFR_X1 \core.keymem.key_mem[2][5]$_DFFE_PN0P_  (.D(_01816_),
    .RN(net100),
    .CK(clknet_leaf_19_clk),
    .Q(\core.keymem.key_mem[2][5] ),
    .QN(_20788_));
 DFFR_X1 \core.keymem.key_mem[2][60]$_DFFE_PN0P_  (.D(_01817_),
    .RN(net89),
    .CK(clknet_leaf_25_clk),
    .Q(\core.keymem.key_mem[2][60] ),
    .QN(_20787_));
 DFFR_X1 \core.keymem.key_mem[2][61]$_DFFE_PN0P_  (.D(_01818_),
    .RN(net89),
    .CK(clknet_leaf_84_clk),
    .Q(\core.keymem.key_mem[2][61] ),
    .QN(_20786_));
 DFFR_X1 \core.keymem.key_mem[2][62]$_DFFE_PN0P_  (.D(_01819_),
    .RN(net100),
    .CK(clknet_leaf_98_clk),
    .Q(\core.keymem.key_mem[2][62] ),
    .QN(_20785_));
 DFFR_X1 \core.keymem.key_mem[2][63]$_DFFE_PN0P_  (.D(_01820_),
    .RN(net100),
    .CK(clknet_leaf_97_clk),
    .Q(\core.keymem.key_mem[2][63] ),
    .QN(_20784_));
 DFFR_X1 \core.keymem.key_mem[2][64]$_DFFE_PN0P_  (.D(_01821_),
    .RN(net100),
    .CK(clknet_leaf_14_clk),
    .Q(\core.keymem.key_mem[2][64] ),
    .QN(_20783_));
 DFFR_X1 \core.keymem.key_mem[2][65]$_DFFE_PN0P_  (.D(_01822_),
    .RN(net99),
    .CK(clknet_leaf_121_clk),
    .Q(\core.keymem.key_mem[2][65] ),
    .QN(_20782_));
 DFFR_X1 \core.keymem.key_mem[2][66]$_DFFE_PN0P_  (.D(_01823_),
    .RN(net100),
    .CK(clknet_leaf_16_clk),
    .Q(\core.keymem.key_mem[2][66] ),
    .QN(_20781_));
 DFFR_X1 \core.keymem.key_mem[2][67]$_DFFE_PN0P_  (.D(_01824_),
    .RN(net95),
    .CK(clknet_leaf_77_clk),
    .Q(\core.keymem.key_mem[2][67] ),
    .QN(_20780_));
 DFFR_X1 \core.keymem.key_mem[2][68]$_DFFE_PN0P_  (.D(_01825_),
    .RN(net95),
    .CK(clknet_leaf_77_clk),
    .Q(\core.keymem.key_mem[2][68] ),
    .QN(_20779_));
 DFFR_X1 \core.keymem.key_mem[2][69]$_DFFE_PN0P_  (.D(_01826_),
    .RN(net98),
    .CK(clknet_leaf_177_clk),
    .Q(\core.keymem.key_mem[2][69] ),
    .QN(_20778_));
 DFFR_X1 \core.keymem.key_mem[2][6]$_DFFE_PN0P_  (.D(_01827_),
    .RN(net100),
    .CK(clknet_leaf_102_clk),
    .Q(\core.keymem.key_mem[2][6] ),
    .QN(_20777_));
 DFFR_X1 \core.keymem.key_mem[2][70]$_DFFE_PN0P_  (.D(_01828_),
    .RN(net100),
    .CK(clknet_leaf_100_clk),
    .Q(\core.keymem.key_mem[2][70] ),
    .QN(_20776_));
 DFFR_X1 \core.keymem.key_mem[2][71]$_DFFE_PN0P_  (.D(_01829_),
    .RN(net99),
    .CK(clknet_leaf_73_clk),
    .Q(\core.keymem.key_mem[2][71] ),
    .QN(_20775_));
 DFFR_X1 \core.keymem.key_mem[2][72]$_DFFE_PN0P_  (.D(_01830_),
    .RN(net95),
    .CK(clknet_leaf_179_clk),
    .Q(\core.keymem.key_mem[2][72] ),
    .QN(_20774_));
 DFFR_X1 \core.keymem.key_mem[2][73]$_DFFE_PN0P_  (.D(_01831_),
    .RN(net97),
    .CK(clknet_leaf_146_clk),
    .Q(\core.keymem.key_mem[2][73] ),
    .QN(_20773_));
 DFFR_X1 \core.keymem.key_mem[2][74]$_DFFE_PN0P_  (.D(_01832_),
    .RN(net97),
    .CK(clknet_leaf_163_clk),
    .Q(\core.keymem.key_mem[2][74] ),
    .QN(_20772_));
 DFFR_X1 \core.keymem.key_mem[2][75]$_DFFE_PN0P_  (.D(_01833_),
    .RN(net97),
    .CK(clknet_leaf_148_clk),
    .Q(\core.keymem.key_mem[2][75] ),
    .QN(_20771_));
 DFFR_X1 \core.keymem.key_mem[2][76]$_DFFE_PN0P_  (.D(_01834_),
    .RN(net91),
    .CK(clknet_leaf_284_clk),
    .Q(\core.keymem.key_mem[2][76] ),
    .QN(_20770_));
 DFFR_X1 \core.keymem.key_mem[2][77]$_DFFE_PN0P_  (.D(_01835_),
    .RN(net97),
    .CK(clknet_leaf_162_clk),
    .Q(\core.keymem.key_mem[2][77] ),
    .QN(_20769_));
 DFFR_X1 \core.keymem.key_mem[2][78]$_DFFE_PN0P_  (.D(_01836_),
    .RN(net97),
    .CK(clknet_leaf_164_clk),
    .Q(\core.keymem.key_mem[2][78] ),
    .QN(_20768_));
 DFFR_X1 \core.keymem.key_mem[2][79]$_DFFE_PN0P_  (.D(_01837_),
    .RN(net98),
    .CK(clknet_leaf_170_clk),
    .Q(\core.keymem.key_mem[2][79] ),
    .QN(_20767_));
 DFFR_X1 \core.keymem.key_mem[2][7]$_DFFE_PN0P_  (.D(_01838_),
    .RN(net98),
    .CK(clknet_leaf_175_clk),
    .Q(\core.keymem.key_mem[2][7] ),
    .QN(_20766_));
 DFFR_X1 \core.keymem.key_mem[2][80]$_DFFE_PN0P_  (.D(_01839_),
    .RN(net97),
    .CK(clknet_leaf_158_clk),
    .Q(\core.keymem.key_mem[2][80] ),
    .QN(_20765_));
 DFFR_X1 \core.keymem.key_mem[2][81]$_DFFE_PN0P_  (.D(_01840_),
    .RN(net97),
    .CK(clknet_leaf_155_clk),
    .Q(\core.keymem.key_mem[2][81] ),
    .QN(_20764_));
 DFFR_X1 \core.keymem.key_mem[2][82]$_DFFE_PN0P_  (.D(_01841_),
    .RN(net98),
    .CK(clknet_leaf_186_clk),
    .Q(\core.keymem.key_mem[2][82] ),
    .QN(_20763_));
 DFFR_X1 \core.keymem.key_mem[2][83]$_DFFE_PN0P_  (.D(_01842_),
    .RN(net94),
    .CK(clknet_leaf_186_clk),
    .Q(\core.keymem.key_mem[2][83] ),
    .QN(_20762_));
 DFFR_X1 \core.keymem.key_mem[2][84]$_DFFE_PN0P_  (.D(_01843_),
    .RN(net94),
    .CK(clknet_leaf_180_clk),
    .Q(\core.keymem.key_mem[2][84] ),
    .QN(_20761_));
 DFFR_X1 \core.keymem.key_mem[2][85]$_DFFE_PN0P_  (.D(_01844_),
    .RN(net94),
    .CK(clknet_leaf_210_clk),
    .Q(\core.keymem.key_mem[2][85] ),
    .QN(_20760_));
 DFFR_X1 \core.keymem.key_mem[2][86]$_DFFE_PN0P_  (.D(_01845_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[2][86] ),
    .QN(_20759_));
 DFFR_X1 \core.keymem.key_mem[2][87]$_DFFE_PN0P_  (.D(_01846_),
    .RN(net93),
    .CK(clknet_leaf_57_clk),
    .Q(\core.keymem.key_mem[2][87] ),
    .QN(_20758_));
 DFFR_X1 \core.keymem.key_mem[2][88]$_DFFE_PN0P_  (.D(_01847_),
    .RN(net93),
    .CK(clknet_leaf_281_clk),
    .Q(\core.keymem.key_mem[2][88] ),
    .QN(_20757_));
 DFFR_X1 \core.keymem.key_mem[2][89]$_DFFE_PN0P_  (.D(_01848_),
    .RN(net93),
    .CK(clknet_leaf_199_clk),
    .Q(\core.keymem.key_mem[2][89] ),
    .QN(_20756_));
 DFFR_X1 \core.keymem.key_mem[2][8]$_DFFE_PN0P_  (.D(_01849_),
    .RN(net89),
    .CK(clknet_leaf_378_clk),
    .Q(\core.keymem.key_mem[2][8] ),
    .QN(_20755_));
 DFFR_X1 \core.keymem.key_mem[2][90]$_DFFE_PN0P_  (.D(_01850_),
    .RN(net97),
    .CK(clknet_leaf_156_clk),
    .Q(\core.keymem.key_mem[2][90] ),
    .QN(_20754_));
 DFFR_X1 \core.keymem.key_mem[2][91]$_DFFE_PN0P_  (.D(_01851_),
    .RN(net93),
    .CK(clknet_leaf_184_clk),
    .Q(\core.keymem.key_mem[2][91] ),
    .QN(_20753_));
 DFFR_X1 \core.keymem.key_mem[2][92]$_DFFE_PN0P_  (.D(_01852_),
    .RN(net95),
    .CK(clknet_leaf_62_clk),
    .Q(\core.keymem.key_mem[2][92] ),
    .QN(_20752_));
 DFFR_X1 \core.keymem.key_mem[2][93]$_DFFE_PN0P_  (.D(_01853_),
    .RN(net95),
    .CK(clknet_leaf_190_clk),
    .Q(\core.keymem.key_mem[2][93] ),
    .QN(_20751_));
 DFFR_X1 \core.keymem.key_mem[2][94]$_DFFE_PN0P_  (.D(_01854_),
    .RN(net94),
    .CK(clknet_leaf_214_clk),
    .Q(\core.keymem.key_mem[2][94] ),
    .QN(_20750_));
 DFFR_X1 \core.keymem.key_mem[2][95]$_DFFE_PN0P_  (.D(_01855_),
    .RN(net96),
    .CK(clknet_leaf_242_clk),
    .Q(\core.keymem.key_mem[2][95] ),
    .QN(_20749_));
 DFFR_X1 \core.keymem.key_mem[2][96]$_DFFE_PN0P_  (.D(_01856_),
    .RN(net92),
    .CK(clknet_leaf_203_clk),
    .Q(\core.keymem.key_mem[2][96] ),
    .QN(_20748_));
 DFFR_X1 \core.keymem.key_mem[2][97]$_DFFE_PN0P_  (.D(_01857_),
    .RN(net93),
    .CK(clknet_leaf_190_clk),
    .Q(\core.keymem.key_mem[2][97] ),
    .QN(_20747_));
 DFFR_X1 \core.keymem.key_mem[2][98]$_DFFE_PN0P_  (.D(_01858_),
    .RN(net93),
    .CK(clknet_leaf_193_clk),
    .Q(\core.keymem.key_mem[2][98] ),
    .QN(_20746_));
 DFFR_X1 \core.keymem.key_mem[2][99]$_DFFE_PN0P_  (.D(_01859_),
    .RN(net91),
    .CK(clknet_leaf_201_clk),
    .Q(\core.keymem.key_mem[2][99] ),
    .QN(_20745_));
 DFFR_X1 \core.keymem.key_mem[2][9]$_DFFE_PN0P_  (.D(_01860_),
    .RN(net91),
    .CK(clknet_leaf_200_clk),
    .Q(\core.keymem.key_mem[2][9] ),
    .QN(_20744_));
 DFFR_X1 \core.keymem.key_mem[3][0]$_DFFE_PN0P_  (.D(_01861_),
    .RN(net94),
    .CK(clknet_leaf_221_clk),
    .Q(\core.keymem.key_mem[3][0] ),
    .QN(_20743_));
 DFFR_X1 \core.keymem.key_mem[3][100]$_DFFE_PN0P_  (.D(_01862_),
    .RN(net94),
    .CK(clknet_leaf_210_clk),
    .Q(\core.keymem.key_mem[3][100] ),
    .QN(_20742_));
 DFFR_X1 \core.keymem.key_mem[3][101]$_DFFE_PN0P_  (.D(_01863_),
    .RN(net94),
    .CK(clknet_leaf_212_clk),
    .Q(\core.keymem.key_mem[3][101] ),
    .QN(_20741_));
 DFFR_X1 \core.keymem.key_mem[3][102]$_DFFE_PN0P_  (.D(_01864_),
    .RN(net96),
    .CK(clknet_leaf_233_clk),
    .Q(\core.keymem.key_mem[3][102] ),
    .QN(_20740_));
 DFFR_X1 \core.keymem.key_mem[3][103]$_DFFE_PN0P_  (.D(_01865_),
    .RN(net96),
    .CK(clknet_leaf_245_clk),
    .Q(\core.keymem.key_mem[3][103] ),
    .QN(_20739_));
 DFFR_X1 \core.keymem.key_mem[3][104]$_DFFE_PN0P_  (.D(_01866_),
    .RN(net92),
    .CK(clknet_leaf_191_clk),
    .Q(\core.keymem.key_mem[3][104] ),
    .QN(_20738_));
 DFFR_X1 \core.keymem.key_mem[3][105]$_DFFE_PN0P_  (.D(_01867_),
    .RN(net96),
    .CK(clknet_leaf_246_clk),
    .Q(\core.keymem.key_mem[3][105] ),
    .QN(_20737_));
 DFFR_X1 \core.keymem.key_mem[3][106]$_DFFE_PN0P_  (.D(_01868_),
    .RN(net92),
    .CK(clknet_leaf_267_clk),
    .Q(\core.keymem.key_mem[3][106] ),
    .QN(_20736_));
 DFFR_X1 \core.keymem.key_mem[3][107]$_DFFE_PN0P_  (.D(_01869_),
    .RN(net92),
    .CK(clknet_leaf_266_clk),
    .Q(\core.keymem.key_mem[3][107] ),
    .QN(_20735_));
 DFFR_X1 \core.keymem.key_mem[3][108]$_DFFE_PN0P_  (.D(_01870_),
    .RN(net91),
    .CK(clknet_leaf_280_clk),
    .Q(\core.keymem.key_mem[3][108] ),
    .QN(_20734_));
 DFFR_X1 \core.keymem.key_mem[3][109]$_DFFE_PN0P_  (.D(_01871_),
    .RN(net94),
    .CK(clknet_leaf_263_clk),
    .Q(\core.keymem.key_mem[3][109] ),
    .QN(_20733_));
 DFFR_X1 \core.keymem.key_mem[3][10]$_DFFE_PN0P_  (.D(_01872_),
    .RN(net95),
    .CK(clknet_leaf_189_clk),
    .Q(\core.keymem.key_mem[3][10] ),
    .QN(_20732_));
 DFFR_X1 \core.keymem.key_mem[3][110]$_DFFE_PN0P_  (.D(_01873_),
    .RN(net96),
    .CK(clknet_leaf_250_clk),
    .Q(\core.keymem.key_mem[3][110] ),
    .QN(_20731_));
 DFFR_X1 \core.keymem.key_mem[3][111]$_DFFE_PN0P_  (.D(_01874_),
    .RN(net96),
    .CK(clknet_leaf_225_clk),
    .Q(\core.keymem.key_mem[3][111] ),
    .QN(_20730_));
 DFFR_X1 \core.keymem.key_mem[3][112]$_DFFE_PN0P_  (.D(_01875_),
    .RN(net94),
    .CK(clknet_leaf_260_clk),
    .Q(\core.keymem.key_mem[3][112] ),
    .QN(_20729_));
 DFFR_X1 \core.keymem.key_mem[3][113]$_DFFE_PN0P_  (.D(_01876_),
    .RN(net91),
    .CK(clknet_leaf_279_clk),
    .Q(\core.keymem.key_mem[3][113] ),
    .QN(_20728_));
 DFFR_X1 \core.keymem.key_mem[3][114]$_DFFE_PN0P_  (.D(_01877_),
    .RN(net91),
    .CK(clknet_leaf_274_clk),
    .Q(\core.keymem.key_mem[3][114] ),
    .QN(_20727_));
 DFFR_X1 \core.keymem.key_mem[3][115]$_DFFE_PN0P_  (.D(_01878_),
    .RN(net92),
    .CK(clknet_leaf_275_clk),
    .Q(\core.keymem.key_mem[3][115] ),
    .QN(_20726_));
 DFFR_X1 \core.keymem.key_mem[3][116]$_DFFE_PN0P_  (.D(_01879_),
    .RN(net92),
    .CK(clknet_leaf_264_clk),
    .Q(\core.keymem.key_mem[3][116] ),
    .QN(_20725_));
 DFFR_X1 \core.keymem.key_mem[3][117]$_DFFE_PN0P_  (.D(_01880_),
    .RN(net94),
    .CK(clknet_leaf_213_clk),
    .Q(\core.keymem.key_mem[3][117] ),
    .QN(_20724_));
 DFFR_X1 \core.keymem.key_mem[3][118]$_DFFE_PN0P_  (.D(_01881_),
    .RN(net98),
    .CK(clknet_leaf_228_clk),
    .Q(\core.keymem.key_mem[3][118] ),
    .QN(_20723_));
 DFFR_X1 \core.keymem.key_mem[3][119]$_DFFE_PN0P_  (.D(_01882_),
    .RN(net94),
    .CK(clknet_leaf_220_clk),
    .Q(\core.keymem.key_mem[3][119] ),
    .QN(_20722_));
 DFFR_X1 \core.keymem.key_mem[3][11]$_DFFE_PN0P_  (.D(_01883_),
    .RN(net95),
    .CK(clknet_leaf_59_clk),
    .Q(\core.keymem.key_mem[3][11] ),
    .QN(_20721_));
 DFFR_X1 \core.keymem.key_mem[3][120]$_DFFE_PN0P_  (.D(_01884_),
    .RN(net93),
    .CK(clknet_leaf_205_clk),
    .Q(\core.keymem.key_mem[3][120] ),
    .QN(_20720_));
 DFFR_X1 \core.keymem.key_mem[3][121]$_DFFE_PN0P_  (.D(_01885_),
    .RN(net92),
    .CK(clknet_leaf_266_clk),
    .Q(\core.keymem.key_mem[3][121] ),
    .QN(_20719_));
 DFFR_X1 \core.keymem.key_mem[3][122]$_DFFE_PN0P_  (.D(_01886_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[3][122] ),
    .QN(_20718_));
 DFFR_X1 \core.keymem.key_mem[3][123]$_DFFE_PN0P_  (.D(_01887_),
    .RN(net93),
    .CK(clknet_leaf_201_clk),
    .Q(\core.keymem.key_mem[3][123] ),
    .QN(_20717_));
 DFFR_X1 \core.keymem.key_mem[3][124]$_DFFE_PN0P_  (.D(_01888_),
    .RN(net93),
    .CK(clknet_leaf_198_clk),
    .Q(\core.keymem.key_mem[3][124] ),
    .QN(_20716_));
 DFFR_X1 \core.keymem.key_mem[3][125]$_DFFE_PN0P_  (.D(_01889_),
    .RN(net97),
    .CK(clknet_leaf_162_clk),
    .Q(\core.keymem.key_mem[3][125] ),
    .QN(_20715_));
 DFFR_X1 \core.keymem.key_mem[3][126]$_DFFE_PN0P_  (.D(_01890_),
    .RN(net98),
    .CK(clknet_leaf_167_clk),
    .Q(\core.keymem.key_mem[3][126] ),
    .QN(_20714_));
 DFFR_X1 \core.keymem.key_mem[3][127]$_DFFE_PN0P_  (.D(_01891_),
    .RN(net97),
    .CK(clknet_leaf_240_clk),
    .Q(\core.keymem.key_mem[3][127] ),
    .QN(_20713_));
 DFFR_X1 \core.keymem.key_mem[3][12]$_DFFE_PN0P_  (.D(_01892_),
    .RN(net93),
    .CK(clknet_leaf_207_clk),
    .Q(\core.keymem.key_mem[3][12] ),
    .QN(_20712_));
 DFFR_X1 \core.keymem.key_mem[3][13]$_DFFE_PN0P_  (.D(_01893_),
    .RN(net85),
    .CK(clknet_leaf_50_clk),
    .Q(\core.keymem.key_mem[3][13] ),
    .QN(_20711_));
 DFFR_X1 \core.keymem.key_mem[3][14]$_DFFE_PN0P_  (.D(_01894_),
    .RN(net89),
    .CK(clknet_leaf_376_clk),
    .Q(\core.keymem.key_mem[3][14] ),
    .QN(_20710_));
 DFFR_X1 \core.keymem.key_mem[3][15]$_DFFE_PN0P_  (.D(_01895_),
    .RN(net96),
    .CK(clknet_leaf_230_clk),
    .Q(\core.keymem.key_mem[3][15] ),
    .QN(_20709_));
 DFFR_X1 \core.keymem.key_mem[3][16]$_DFFE_PN0P_  (.D(_01896_),
    .RN(net89),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[3][16] ),
    .QN(_20708_));
 DFFR_X1 \core.keymem.key_mem[3][17]$_DFFE_PN0P_  (.D(_01897_),
    .RN(net98),
    .CK(clknet_leaf_167_clk),
    .Q(\core.keymem.key_mem[3][17] ),
    .QN(_20707_));
 DFFR_X1 \core.keymem.key_mem[3][18]$_DFFE_PN0P_  (.D(_01898_),
    .RN(net82),
    .CK(clknet_leaf_35_clk),
    .Q(\core.keymem.key_mem[3][18] ),
    .QN(_20706_));
 DFFR_X1 \core.keymem.key_mem[3][19]$_DFFE_PN0P_  (.D(_01899_),
    .RN(net89),
    .CK(clknet_leaf_59_clk),
    .Q(\core.keymem.key_mem[3][19] ),
    .QN(_20705_));
 DFFR_X1 \core.keymem.key_mem[3][1]$_DFFE_PN0P_  (.D(_01900_),
    .RN(net82),
    .CK(clknet_leaf_10_clk),
    .Q(\core.keymem.key_mem[3][1] ),
    .QN(_20704_));
 DFFR_X1 \core.keymem.key_mem[3][20]$_DFFE_PN0P_  (.D(_01901_),
    .RN(net89),
    .CK(clknet_leaf_92_clk),
    .Q(\core.keymem.key_mem[3][20] ),
    .QN(_20703_));
 DFFR_X1 \core.keymem.key_mem[3][21]$_DFFE_PN0P_  (.D(_01902_),
    .RN(net85),
    .CK(clknet_leaf_67_clk),
    .Q(\core.keymem.key_mem[3][21] ),
    .QN(_20702_));
 DFFR_X1 \core.keymem.key_mem[3][22]$_DFFE_PN0P_  (.D(_01903_),
    .RN(net94),
    .CK(clknet_leaf_219_clk),
    .Q(\core.keymem.key_mem[3][22] ),
    .QN(_20701_));
 DFFR_X1 \core.keymem.key_mem[3][23]$_DFFE_PN0P_  (.D(_01904_),
    .RN(net93),
    .CK(clknet_leaf_59_clk),
    .Q(\core.keymem.key_mem[3][23] ),
    .QN(_20700_));
 DFFR_X1 \core.keymem.key_mem[3][24]$_DFFE_PN0P_  (.D(_01905_),
    .RN(net89),
    .CK(clknet_leaf_65_clk),
    .Q(\core.keymem.key_mem[3][24] ),
    .QN(_20699_));
 DFFR_X1 \core.keymem.key_mem[3][25]$_DFFE_PN0P_  (.D(_01906_),
    .RN(net85),
    .CK(clknet_leaf_49_clk),
    .Q(\core.keymem.key_mem[3][25] ),
    .QN(_20698_));
 DFFR_X1 \core.keymem.key_mem[3][26]$_DFFE_PN0P_  (.D(_01907_),
    .RN(net89),
    .CK(clknet_leaf_96_clk),
    .Q(\core.keymem.key_mem[3][26] ),
    .QN(_20697_));
 DFFR_X1 \core.keymem.key_mem[3][27]$_DFFE_PN0P_  (.D(_01908_),
    .RN(net16),
    .CK(clknet_leaf_151_clk),
    .Q(\core.keymem.key_mem[3][27] ),
    .QN(_20696_));
 DFFR_X1 \core.keymem.key_mem[3][28]$_DFFE_PN0P_  (.D(_01909_),
    .RN(net16),
    .CK(clknet_leaf_131_clk),
    .Q(\core.keymem.key_mem[3][28] ),
    .QN(_20695_));
 DFFR_X1 \core.keymem.key_mem[3][29]$_DFFE_PN0P_  (.D(_01910_),
    .RN(net97),
    .CK(clknet_leaf_148_clk),
    .Q(\core.keymem.key_mem[3][29] ),
    .QN(_20694_));
 DFFR_X1 \core.keymem.key_mem[3][2]$_DFFE_PN0P_  (.D(_01911_),
    .RN(net89),
    .CK(clknet_leaf_66_clk),
    .Q(\core.keymem.key_mem[3][2] ),
    .QN(_20693_));
 DFFR_X1 \core.keymem.key_mem[3][30]$_DFFE_PN0P_  (.D(_01912_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[3][30] ),
    .QN(_20692_));
 DFFR_X1 \core.keymem.key_mem[3][31]$_DFFE_PN0P_  (.D(_01913_),
    .RN(net98),
    .CK(clknet_leaf_144_clk),
    .Q(\core.keymem.key_mem[3][31] ),
    .QN(_20691_));
 DFFR_X1 \core.keymem.key_mem[3][32]$_DFFE_PN0P_  (.D(_01914_),
    .RN(net99),
    .CK(clknet_leaf_112_clk),
    .Q(\core.keymem.key_mem[3][32] ),
    .QN(_20690_));
 DFFR_X1 \core.keymem.key_mem[3][33]$_DFFE_PN0P_  (.D(_01915_),
    .RN(net16),
    .CK(clknet_leaf_126_clk),
    .Q(\core.keymem.key_mem[3][33] ),
    .QN(_20689_));
 DFFR_X1 \core.keymem.key_mem[3][34]$_DFFE_PN0P_  (.D(_01916_),
    .RN(net16),
    .CK(clknet_leaf_137_clk),
    .Q(\core.keymem.key_mem[3][34] ),
    .QN(_20688_));
 DFFR_X1 \core.keymem.key_mem[3][35]$_DFFE_PN0P_  (.D(_01917_),
    .RN(net99),
    .CK(clknet_leaf_122_clk),
    .Q(\core.keymem.key_mem[3][35] ),
    .QN(_20687_));
 DFFR_X1 \core.keymem.key_mem[3][36]$_DFFE_PN0P_  (.D(_01918_),
    .RN(net88),
    .CK(clknet_leaf_90_clk),
    .Q(\core.keymem.key_mem[3][36] ),
    .QN(_20686_));
 DFFR_X1 \core.keymem.key_mem[3][37]$_DFFE_PN0P_  (.D(_01919_),
    .RN(net88),
    .CK(clknet_leaf_92_clk),
    .Q(\core.keymem.key_mem[3][37] ),
    .QN(_20685_));
 DFFR_X1 \core.keymem.key_mem[3][38]$_DFFE_PN0P_  (.D(_01920_),
    .RN(net16),
    .CK(clknet_leaf_124_clk),
    .Q(\core.keymem.key_mem[3][38] ),
    .QN(_20684_));
 DFFR_X1 \core.keymem.key_mem[3][39]$_DFFE_PN0P_  (.D(_01921_),
    .RN(net89),
    .CK(clknet_leaf_85_clk),
    .Q(\core.keymem.key_mem[3][39] ),
    .QN(_20683_));
 DFFR_X1 \core.keymem.key_mem[3][3]$_DFFE_PN0P_  (.D(_01922_),
    .RN(net88),
    .CK(clknet_leaf_91_clk),
    .Q(\core.keymem.key_mem[3][3] ),
    .QN(_20682_));
 DFFR_X1 \core.keymem.key_mem[3][40]$_DFFE_PN0P_  (.D(_01923_),
    .RN(net88),
    .CK(clknet_leaf_89_clk),
    .Q(\core.keymem.key_mem[3][40] ),
    .QN(_20681_));
 DFFR_X1 \core.keymem.key_mem[3][41]$_DFFE_PN0P_  (.D(_01924_),
    .RN(net89),
    .CK(clknet_leaf_82_clk),
    .Q(\core.keymem.key_mem[3][41] ),
    .QN(_20680_));
 DFFR_X1 \core.keymem.key_mem[3][42]$_DFFE_PN0P_  (.D(_01925_),
    .RN(net99),
    .CK(clknet_leaf_117_clk),
    .Q(\core.keymem.key_mem[3][42] ),
    .QN(_20679_));
 DFFR_X1 \core.keymem.key_mem[3][43]$_DFFE_PN0P_  (.D(_01926_),
    .RN(net85),
    .CK(clknet_leaf_67_clk),
    .Q(\core.keymem.key_mem[3][43] ),
    .QN(_20678_));
 DFFR_X1 \core.keymem.key_mem[3][44]$_DFFE_PN0P_  (.D(_01927_),
    .RN(net100),
    .CK(clknet_leaf_114_clk),
    .Q(\core.keymem.key_mem[3][44] ),
    .QN(_20677_));
 DFFR_X1 \core.keymem.key_mem[3][45]$_DFFE_PN0P_  (.D(_01928_),
    .RN(net99),
    .CK(clknet_leaf_71_clk),
    .Q(\core.keymem.key_mem[3][45] ),
    .QN(_20676_));
 DFFR_X1 \core.keymem.key_mem[3][46]$_DFFE_PN0P_  (.D(_01929_),
    .RN(net99),
    .CK(clknet_leaf_86_clk),
    .Q(\core.keymem.key_mem[3][46] ),
    .QN(_20675_));
 DFFR_X1 \core.keymem.key_mem[3][47]$_DFFE_PN0P_  (.D(_01930_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[3][47] ),
    .QN(_20674_));
 DFFR_X1 \core.keymem.key_mem[3][48]$_DFFE_PN0P_  (.D(_01931_),
    .RN(net95),
    .CK(clknet_leaf_120_clk),
    .Q(\core.keymem.key_mem[3][48] ),
    .QN(_20673_));
 DFFR_X1 \core.keymem.key_mem[3][49]$_DFFE_PN0P_  (.D(_01932_),
    .RN(net99),
    .CK(clknet_leaf_118_clk),
    .Q(\core.keymem.key_mem[3][49] ),
    .QN(_20672_));
 DFFR_X1 \core.keymem.key_mem[3][4]$_DFFE_PN0P_  (.D(_01933_),
    .RN(net100),
    .CK(clknet_leaf_104_clk),
    .Q(\core.keymem.key_mem[3][4] ),
    .QN(_20671_));
 DFFR_X1 \core.keymem.key_mem[3][50]$_DFFE_PN0P_  (.D(_01934_),
    .RN(net98),
    .CK(clknet_leaf_139_clk),
    .Q(\core.keymem.key_mem[3][50] ),
    .QN(_20670_));
 DFFR_X1 \core.keymem.key_mem[3][51]$_DFFE_PN0P_  (.D(_01935_),
    .RN(net16),
    .CK(clknet_leaf_126_clk),
    .Q(\core.keymem.key_mem[3][51] ),
    .QN(_20669_));
 DFFR_X1 \core.keymem.key_mem[3][52]$_DFFE_PN0P_  (.D(_01936_),
    .RN(net89),
    .CK(clknet_leaf_83_clk),
    .Q(\core.keymem.key_mem[3][52] ),
    .QN(_20668_));
 DFFR_X1 \core.keymem.key_mem[3][53]$_DFFE_PN0P_  (.D(_01937_),
    .RN(net97),
    .CK(clknet_leaf_145_clk),
    .Q(\core.keymem.key_mem[3][53] ),
    .QN(_20667_));
 DFFR_X1 \core.keymem.key_mem[3][54]$_DFFE_PN0P_  (.D(_01938_),
    .RN(net98),
    .CK(clknet_leaf_143_clk),
    .Q(\core.keymem.key_mem[3][54] ),
    .QN(_20666_));
 DFFR_X1 \core.keymem.key_mem[3][55]$_DFFE_PN0P_  (.D(_01939_),
    .RN(net16),
    .CK(clknet_leaf_136_clk),
    .Q(\core.keymem.key_mem[3][55] ),
    .QN(_20665_));
 DFFR_X1 \core.keymem.key_mem[3][56]$_DFFE_PN0P_  (.D(_01940_),
    .RN(net97),
    .CK(clknet_leaf_144_clk),
    .Q(\core.keymem.key_mem[3][56] ),
    .QN(_20664_));
 DFFR_X1 \core.keymem.key_mem[3][57]$_DFFE_PN0P_  (.D(_01941_),
    .RN(net100),
    .CK(clknet_leaf_109_clk),
    .Q(\core.keymem.key_mem[3][57] ),
    .QN(_20663_));
 DFFR_X1 \core.keymem.key_mem[3][58]$_DFFE_PN0P_  (.D(_01942_),
    .RN(net100),
    .CK(clknet_leaf_102_clk),
    .Q(\core.keymem.key_mem[3][58] ),
    .QN(_20662_));
 DFFR_X1 \core.keymem.key_mem[3][59]$_DFFE_PN0P_  (.D(_01943_),
    .RN(net89),
    .CK(clknet_leaf_25_clk),
    .Q(\core.keymem.key_mem[3][59] ),
    .QN(_20661_));
 DFFR_X1 \core.keymem.key_mem[3][5]$_DFFE_PN0P_  (.D(_01944_),
    .RN(net100),
    .CK(clknet_leaf_19_clk),
    .Q(\core.keymem.key_mem[3][5] ),
    .QN(_20660_));
 DFFR_X1 \core.keymem.key_mem[3][60]$_DFFE_PN0P_  (.D(_01945_),
    .RN(net89),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[3][60] ),
    .QN(_20659_));
 DFFR_X1 \core.keymem.key_mem[3][61]$_DFFE_PN0P_  (.D(_01946_),
    .RN(net89),
    .CK(clknet_leaf_84_clk),
    .Q(\core.keymem.key_mem[3][61] ),
    .QN(_20658_));
 DFFR_X1 \core.keymem.key_mem[3][62]$_DFFE_PN0P_  (.D(_01947_),
    .RN(net100),
    .CK(clknet_leaf_98_clk),
    .Q(\core.keymem.key_mem[3][62] ),
    .QN(_20657_));
 DFFR_X1 \core.keymem.key_mem[3][63]$_DFFE_PN0P_  (.D(_01948_),
    .RN(net100),
    .CK(clknet_leaf_20_clk),
    .Q(\core.keymem.key_mem[3][63] ),
    .QN(_20656_));
 DFFR_X1 \core.keymem.key_mem[3][64]$_DFFE_PN0P_  (.D(_01949_),
    .RN(net100),
    .CK(clknet_leaf_14_clk),
    .Q(\core.keymem.key_mem[3][64] ),
    .QN(_20655_));
 DFFR_X1 \core.keymem.key_mem[3][65]$_DFFE_PN0P_  (.D(_01950_),
    .RN(net98),
    .CK(clknet_leaf_121_clk),
    .Q(\core.keymem.key_mem[3][65] ),
    .QN(_20654_));
 DFFR_X1 \core.keymem.key_mem[3][66]$_DFFE_PN0P_  (.D(_01951_),
    .RN(net100),
    .CK(clknet_leaf_15_clk),
    .Q(\core.keymem.key_mem[3][66] ),
    .QN(_20653_));
 DFFR_X1 \core.keymem.key_mem[3][67]$_DFFE_PN0P_  (.D(_01952_),
    .RN(net95),
    .CK(clknet_leaf_76_clk),
    .Q(\core.keymem.key_mem[3][67] ),
    .QN(_20652_));
 DFFR_X1 \core.keymem.key_mem[3][68]$_DFFE_PN0P_  (.D(_01953_),
    .RN(net99),
    .CK(clknet_leaf_116_clk),
    .Q(\core.keymem.key_mem[3][68] ),
    .QN(_20651_));
 DFFR_X1 \core.keymem.key_mem[3][69]$_DFFE_PN0P_  (.D(_01954_),
    .RN(net95),
    .CK(clknet_leaf_177_clk),
    .Q(\core.keymem.key_mem[3][69] ),
    .QN(_20650_));
 DFFR_X1 \core.keymem.key_mem[3][6]$_DFFE_PN0P_  (.D(_01955_),
    .RN(net100),
    .CK(clknet_leaf_102_clk),
    .Q(\core.keymem.key_mem[3][6] ),
    .QN(_20649_));
 DFFR_X1 \core.keymem.key_mem[3][70]$_DFFE_PN0P_  (.D(_01956_),
    .RN(net100),
    .CK(clknet_leaf_100_clk),
    .Q(\core.keymem.key_mem[3][70] ),
    .QN(_20648_));
 DFFR_X1 \core.keymem.key_mem[3][71]$_DFFE_PN0P_  (.D(_01957_),
    .RN(net99),
    .CK(clknet_leaf_73_clk),
    .Q(\core.keymem.key_mem[3][71] ),
    .QN(_20647_));
 DFFR_X1 \core.keymem.key_mem[3][72]$_DFFE_PN0P_  (.D(_01958_),
    .RN(net95),
    .CK(clknet_leaf_178_clk),
    .Q(\core.keymem.key_mem[3][72] ),
    .QN(_20646_));
 DFFR_X1 \core.keymem.key_mem[3][73]$_DFFE_PN0P_  (.D(_01959_),
    .RN(net97),
    .CK(clknet_leaf_152_clk),
    .Q(\core.keymem.key_mem[3][73] ),
    .QN(_20645_));
 DFFR_X1 \core.keymem.key_mem[3][74]$_DFFE_PN0P_  (.D(_01960_),
    .RN(net97),
    .CK(clknet_leaf_156_clk),
    .Q(\core.keymem.key_mem[3][74] ),
    .QN(_20644_));
 DFFR_X1 \core.keymem.key_mem[3][75]$_DFFE_PN0P_  (.D(_01961_),
    .RN(net97),
    .CK(clknet_leaf_152_clk),
    .Q(\core.keymem.key_mem[3][75] ),
    .QN(_20643_));
 DFFR_X1 \core.keymem.key_mem[3][76]$_DFFE_PN0P_  (.D(_01962_),
    .RN(net91),
    .CK(clknet_leaf_284_clk),
    .Q(\core.keymem.key_mem[3][76] ),
    .QN(_20642_));
 DFFR_X1 \core.keymem.key_mem[3][77]$_DFFE_PN0P_  (.D(_01963_),
    .RN(net97),
    .CK(clknet_leaf_161_clk),
    .Q(\core.keymem.key_mem[3][77] ),
    .QN(_20641_));
 DFFR_X1 \core.keymem.key_mem[3][78]$_DFFE_PN0P_  (.D(_01964_),
    .RN(net98),
    .CK(clknet_leaf_170_clk),
    .Q(\core.keymem.key_mem[3][78] ),
    .QN(_20640_));
 DFFR_X1 \core.keymem.key_mem[3][79]$_DFFE_PN0P_  (.D(_01965_),
    .RN(net98),
    .CK(clknet_leaf_170_clk),
    .Q(\core.keymem.key_mem[3][79] ),
    .QN(_20639_));
 DFFR_X1 \core.keymem.key_mem[3][7]$_DFFE_PN0P_  (.D(_01966_),
    .RN(net98),
    .CK(clknet_leaf_170_clk),
    .Q(\core.keymem.key_mem[3][7] ),
    .QN(_20638_));
 DFFR_X1 \core.keymem.key_mem[3][80]$_DFFE_PN0P_  (.D(_01967_),
    .RN(net97),
    .CK(clknet_leaf_157_clk),
    .Q(\core.keymem.key_mem[3][80] ),
    .QN(_20637_));
 DFFR_X1 \core.keymem.key_mem[3][81]$_DFFE_PN0P_  (.D(_01968_),
    .RN(net97),
    .CK(clknet_leaf_157_clk),
    .Q(\core.keymem.key_mem[3][81] ),
    .QN(_20636_));
 DFFR_X1 \core.keymem.key_mem[3][82]$_DFFE_PN0P_  (.D(_01969_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[3][82] ),
    .QN(_20635_));
 DFFR_X1 \core.keymem.key_mem[3][83]$_DFFE_PN0P_  (.D(_01970_),
    .RN(net93),
    .CK(clknet_leaf_184_clk),
    .Q(\core.keymem.key_mem[3][83] ),
    .QN(_20634_));
 DFFR_X1 \core.keymem.key_mem[3][84]$_DFFE_PN0P_  (.D(_01971_),
    .RN(net95),
    .CK(clknet_leaf_182_clk),
    .Q(\core.keymem.key_mem[3][84] ),
    .QN(_20633_));
 DFFR_X1 \core.keymem.key_mem[3][85]$_DFFE_PN0P_  (.D(_01972_),
    .RN(net94),
    .CK(clknet_leaf_209_clk),
    .Q(\core.keymem.key_mem[3][85] ),
    .QN(_20632_));
 DFFR_X1 \core.keymem.key_mem[3][86]$_DFFE_PN0P_  (.D(_01973_),
    .RN(net98),
    .CK(clknet_leaf_229_clk),
    .Q(\core.keymem.key_mem[3][86] ),
    .QN(_20631_));
 DFFR_X1 \core.keymem.key_mem[3][87]$_DFFE_PN0P_  (.D(_01974_),
    .RN(net93),
    .CK(clknet_leaf_57_clk),
    .Q(\core.keymem.key_mem[3][87] ),
    .QN(_20630_));
 DFFR_X1 \core.keymem.key_mem[3][88]$_DFFE_PN0P_  (.D(_01975_),
    .RN(net93),
    .CK(clknet_leaf_281_clk),
    .Q(\core.keymem.key_mem[3][88] ),
    .QN(_20629_));
 DFFR_X1 \core.keymem.key_mem[3][89]$_DFFE_PN0P_  (.D(_01976_),
    .RN(net93),
    .CK(clknet_leaf_199_clk),
    .Q(\core.keymem.key_mem[3][89] ),
    .QN(_20628_));
 DFFR_X1 \core.keymem.key_mem[3][8]$_DFFE_PN0P_  (.D(_01977_),
    .RN(net93),
    .CK(clknet_leaf_57_clk),
    .Q(\core.keymem.key_mem[3][8] ),
    .QN(_20627_));
 DFFR_X1 \core.keymem.key_mem[3][90]$_DFFE_PN0P_  (.D(_01978_),
    .RN(net97),
    .CK(clknet_leaf_156_clk),
    .Q(\core.keymem.key_mem[3][90] ),
    .QN(_20626_));
 DFFR_X1 \core.keymem.key_mem[3][91]$_DFFE_PN0P_  (.D(_01979_),
    .RN(net93),
    .CK(clknet_leaf_185_clk),
    .Q(\core.keymem.key_mem[3][91] ),
    .QN(_20625_));
 DFFR_X1 \core.keymem.key_mem[3][92]$_DFFE_PN0P_  (.D(_01980_),
    .RN(net95),
    .CK(clknet_leaf_61_clk),
    .Q(\core.keymem.key_mem[3][92] ),
    .QN(_20624_));
 DFFR_X1 \core.keymem.key_mem[3][93]$_DFFE_PN0P_  (.D(_01981_),
    .RN(net95),
    .CK(clknet_leaf_190_clk),
    .Q(\core.keymem.key_mem[3][93] ),
    .QN(_20623_));
 DFFR_X1 \core.keymem.key_mem[3][94]$_DFFE_PN0P_  (.D(_01982_),
    .RN(net94),
    .CK(clknet_leaf_214_clk),
    .Q(\core.keymem.key_mem[3][94] ),
    .QN(_20622_));
 DFFR_X1 \core.keymem.key_mem[3][95]$_DFFE_PN0P_  (.D(_01983_),
    .RN(net96),
    .CK(clknet_leaf_234_clk),
    .Q(\core.keymem.key_mem[3][95] ),
    .QN(_20621_));
 DFFR_X1 \core.keymem.key_mem[3][96]$_DFFE_PN0P_  (.D(_01984_),
    .RN(net92),
    .CK(clknet_leaf_203_clk),
    .Q(\core.keymem.key_mem[3][96] ),
    .QN(_20620_));
 DFFR_X1 \core.keymem.key_mem[3][97]$_DFFE_PN0P_  (.D(_01985_),
    .RN(net93),
    .CK(clknet_leaf_192_clk),
    .Q(\core.keymem.key_mem[3][97] ),
    .QN(_20619_));
 DFFR_X1 \core.keymem.key_mem[3][98]$_DFFE_PN0P_  (.D(_01986_),
    .RN(net93),
    .CK(clknet_leaf_195_clk),
    .Q(\core.keymem.key_mem[3][98] ),
    .QN(_20618_));
 DFFR_X1 \core.keymem.key_mem[3][99]$_DFFE_PN0P_  (.D(_01987_),
    .RN(net91),
    .CK(clknet_leaf_201_clk),
    .Q(\core.keymem.key_mem[3][99] ),
    .QN(_20617_));
 DFFR_X1 \core.keymem.key_mem[3][9]$_DFFE_PN0P_  (.D(_01988_),
    .RN(net91),
    .CK(clknet_leaf_200_clk),
    .Q(\core.keymem.key_mem[3][9] ),
    .QN(_20616_));
 DFFR_X1 \core.keymem.key_mem[4][0]$_DFFE_PN0P_  (.D(_01989_),
    .RN(net96),
    .CK(clknet_leaf_248_clk),
    .Q(\core.keymem.key_mem[4][0] ),
    .QN(_20615_));
 DFFR_X1 \core.keymem.key_mem[4][100]$_DFFE_PN0P_  (.D(_01990_),
    .RN(net94),
    .CK(clknet_leaf_212_clk),
    .Q(\core.keymem.key_mem[4][100] ),
    .QN(_20614_));
 DFFR_X1 \core.keymem.key_mem[4][101]$_DFFE_PN0P_  (.D(_01991_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[4][101] ),
    .QN(_20613_));
 DFFR_X1 \core.keymem.key_mem[4][102]$_DFFE_PN0P_  (.D(_01992_),
    .RN(net96),
    .CK(clknet_leaf_233_clk),
    .Q(\core.keymem.key_mem[4][102] ),
    .QN(_20612_));
 DFFR_X1 \core.keymem.key_mem[4][103]$_DFFE_PN0P_  (.D(_01993_),
    .RN(net96),
    .CK(clknet_leaf_245_clk),
    .Q(\core.keymem.key_mem[4][103] ),
    .QN(_20611_));
 DFFR_X1 \core.keymem.key_mem[4][104]$_DFFE_PN0P_  (.D(_01994_),
    .RN(net93),
    .CK(clknet_leaf_192_clk),
    .Q(\core.keymem.key_mem[4][104] ),
    .QN(_20610_));
 DFFR_X1 \core.keymem.key_mem[4][105]$_DFFE_PN0P_  (.D(_01995_),
    .RN(net96),
    .CK(clknet_leaf_247_clk),
    .Q(\core.keymem.key_mem[4][105] ),
    .QN(_20609_));
 DFFR_X1 \core.keymem.key_mem[4][106]$_DFFE_PN0P_  (.D(_01996_),
    .RN(net92),
    .CK(clknet_leaf_268_clk),
    .Q(\core.keymem.key_mem[4][106] ),
    .QN(_20608_));
 DFFR_X1 \core.keymem.key_mem[4][107]$_DFFE_PN0P_  (.D(_01997_),
    .RN(net92),
    .CK(clknet_leaf_269_clk),
    .Q(\core.keymem.key_mem[4][107] ),
    .QN(_20607_));
 DFFR_X1 \core.keymem.key_mem[4][108]$_DFFE_PN0P_  (.D(_01998_),
    .RN(net91),
    .CK(clknet_leaf_278_clk),
    .Q(\core.keymem.key_mem[4][108] ),
    .QN(_20606_));
 DFFR_X1 \core.keymem.key_mem[4][109]$_DFFE_PN0P_  (.D(_01999_),
    .RN(net94),
    .CK(clknet_leaf_258_clk),
    .Q(\core.keymem.key_mem[4][109] ),
    .QN(_20605_));
 DFFR_X1 \core.keymem.key_mem[4][10]$_DFFE_PN0P_  (.D(_02000_),
    .RN(net98),
    .CK(clknet_leaf_188_clk),
    .Q(\core.keymem.key_mem[4][10] ),
    .QN(_20604_));
 DFFR_X1 \core.keymem.key_mem[4][110]$_DFFE_PN0P_  (.D(_02001_),
    .RN(net96),
    .CK(clknet_leaf_250_clk),
    .Q(\core.keymem.key_mem[4][110] ),
    .QN(_20603_));
 DFFR_X1 \core.keymem.key_mem[4][111]$_DFFE_PN0P_  (.D(_02002_),
    .RN(net96),
    .CK(clknet_leaf_225_clk),
    .Q(\core.keymem.key_mem[4][111] ),
    .QN(_20602_));
 DFFR_X1 \core.keymem.key_mem[4][112]$_DFFE_PN0P_  (.D(_02003_),
    .RN(net94),
    .CK(clknet_leaf_260_clk),
    .Q(\core.keymem.key_mem[4][112] ),
    .QN(_20601_));
 DFFR_X1 \core.keymem.key_mem[4][113]$_DFFE_PN0P_  (.D(_02004_),
    .RN(net92),
    .CK(clknet_leaf_273_clk),
    .Q(\core.keymem.key_mem[4][113] ),
    .QN(_20600_));
 DFFR_X1 \core.keymem.key_mem[4][114]$_DFFE_PN0P_  (.D(_02005_),
    .RN(net91),
    .CK(clknet_leaf_274_clk),
    .Q(\core.keymem.key_mem[4][114] ),
    .QN(_20599_));
 DFFR_X1 \core.keymem.key_mem[4][115]$_DFFE_PN0P_  (.D(_02006_),
    .RN(net92),
    .CK(clknet_leaf_274_clk),
    .Q(\core.keymem.key_mem[4][115] ),
    .QN(_20598_));
 DFFR_X1 \core.keymem.key_mem[4][116]$_DFFE_PN0P_  (.D(_02007_),
    .RN(net94),
    .CK(clknet_leaf_264_clk),
    .Q(\core.keymem.key_mem[4][116] ),
    .QN(_20597_));
 DFFR_X1 \core.keymem.key_mem[4][117]$_DFFE_PN0P_  (.D(_02008_),
    .RN(net96),
    .CK(clknet_leaf_222_clk),
    .Q(\core.keymem.key_mem[4][117] ),
    .QN(_20596_));
 DFFR_X1 \core.keymem.key_mem[4][118]$_DFFE_PN0P_  (.D(_02009_),
    .RN(net97),
    .CK(clknet_leaf_241_clk),
    .Q(\core.keymem.key_mem[4][118] ),
    .QN(_20595_));
 DFFR_X1 \core.keymem.key_mem[4][119]$_DFFE_PN0P_  (.D(_02010_),
    .RN(net94),
    .CK(clknet_leaf_220_clk),
    .Q(\core.keymem.key_mem[4][119] ),
    .QN(_20594_));
 DFFR_X1 \core.keymem.key_mem[4][11]$_DFFE_PN0P_  (.D(_02011_),
    .RN(net95),
    .CK(clknet_leaf_61_clk),
    .Q(\core.keymem.key_mem[4][11] ),
    .QN(_20593_));
 DFFR_X1 \core.keymem.key_mem[4][120]$_DFFE_PN0P_  (.D(_02012_),
    .RN(net94),
    .CK(clknet_leaf_216_clk),
    .Q(\core.keymem.key_mem[4][120] ),
    .QN(_20592_));
 DFFR_X1 \core.keymem.key_mem[4][121]$_DFFE_PN0P_  (.D(_02013_),
    .RN(net94),
    .CK(clknet_leaf_264_clk),
    .Q(\core.keymem.key_mem[4][121] ),
    .QN(_20591_));
 DFFR_X1 \core.keymem.key_mem[4][122]$_DFFE_PN0P_  (.D(_02014_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[4][122] ),
    .QN(_20590_));
 DFFR_X1 \core.keymem.key_mem[4][123]$_DFFE_PN0P_  (.D(_02015_),
    .RN(net93),
    .CK(clknet_leaf_197_clk),
    .Q(\core.keymem.key_mem[4][123] ),
    .QN(_20589_));
 DFFR_X1 \core.keymem.key_mem[4][124]$_DFFE_PN0P_  (.D(_02016_),
    .RN(net93),
    .CK(clknet_leaf_198_clk),
    .Q(\core.keymem.key_mem[4][124] ),
    .QN(_20588_));
 DFFR_X1 \core.keymem.key_mem[4][125]$_DFFE_PN0P_  (.D(_02017_),
    .RN(net96),
    .CK(clknet_leaf_236_clk),
    .Q(\core.keymem.key_mem[4][125] ),
    .QN(_20587_));
 DFFR_X1 \core.keymem.key_mem[4][126]$_DFFE_PN0P_  (.D(_02018_),
    .RN(net98),
    .CK(clknet_leaf_188_clk),
    .Q(\core.keymem.key_mem[4][126] ),
    .QN(_20586_));
 DFFR_X1 \core.keymem.key_mem[4][127]$_DFFE_PN0P_  (.D(_02019_),
    .RN(net97),
    .CK(clknet_leaf_240_clk),
    .Q(\core.keymem.key_mem[4][127] ),
    .QN(_20585_));
 DFFR_X1 \core.keymem.key_mem[4][12]$_DFFE_PN0P_  (.D(_02020_),
    .RN(net93),
    .CK(clknet_leaf_206_clk),
    .Q(\core.keymem.key_mem[4][12] ),
    .QN(_20584_));
 DFFR_X1 \core.keymem.key_mem[4][13]$_DFFE_PN0P_  (.D(_02021_),
    .RN(net88),
    .CK(clknet_leaf_30_clk),
    .Q(\core.keymem.key_mem[4][13] ),
    .QN(_20583_));
 DFFR_X1 \core.keymem.key_mem[4][14]$_DFFE_PN0P_  (.D(_02022_),
    .RN(net94),
    .CK(clknet_leaf_212_clk),
    .Q(\core.keymem.key_mem[4][14] ),
    .QN(_20582_));
 DFFR_X1 \core.keymem.key_mem[4][15]$_DFFE_PN0P_  (.D(_02023_),
    .RN(net96),
    .CK(clknet_leaf_165_clk),
    .Q(\core.keymem.key_mem[4][15] ),
    .QN(_20581_));
 DFFR_X1 \core.keymem.key_mem[4][16]$_DFFE_PN0P_  (.D(_02024_),
    .RN(net87),
    .CK(clknet_leaf_28_clk),
    .Q(\core.keymem.key_mem[4][16] ),
    .QN(_20580_));
 DFFR_X1 \core.keymem.key_mem[4][17]$_DFFE_PN0P_  (.D(_02025_),
    .RN(net98),
    .CK(clknet_leaf_187_clk),
    .Q(\core.keymem.key_mem[4][17] ),
    .QN(_20579_));
 DFFR_X1 \core.keymem.key_mem[4][18]$_DFFE_PN0P_  (.D(_02026_),
    .RN(net89),
    .CK(clknet_leaf_25_clk),
    .Q(\core.keymem.key_mem[4][18] ),
    .QN(_20578_));
 DFFR_X1 \core.keymem.key_mem[4][19]$_DFFE_PN0P_  (.D(_02027_),
    .RN(net89),
    .CK(clknet_leaf_65_clk),
    .Q(\core.keymem.key_mem[4][19] ),
    .QN(_20577_));
 DFFR_X1 \core.keymem.key_mem[4][1]$_DFFE_PN0P_  (.D(_02028_),
    .RN(net100),
    .CK(clknet_leaf_23_clk),
    .Q(\core.keymem.key_mem[4][1] ),
    .QN(_20576_));
 DFFR_X1 \core.keymem.key_mem[4][20]$_DFFE_PN0P_  (.D(_02029_),
    .RN(net100),
    .CK(clknet_leaf_22_clk),
    .Q(\core.keymem.key_mem[4][20] ),
    .QN(_20575_));
 DFFR_X1 \core.keymem.key_mem[4][21]$_DFFE_PN0P_  (.D(_02030_),
    .RN(net89),
    .CK(clknet_leaf_66_clk),
    .Q(\core.keymem.key_mem[4][21] ),
    .QN(_20574_));
 DFFR_X1 \core.keymem.key_mem[4][22]$_DFFE_PN0P_  (.D(_02031_),
    .RN(net96),
    .CK(clknet_leaf_249_clk),
    .Q(\core.keymem.key_mem[4][22] ),
    .QN(_20573_));
 DFFR_X1 \core.keymem.key_mem[4][23]$_DFFE_PN0P_  (.D(_02032_),
    .RN(net89),
    .CK(clknet_leaf_53_clk),
    .Q(\core.keymem.key_mem[4][23] ),
    .QN(_20572_));
 DFFR_X1 \core.keymem.key_mem[4][24]$_DFFE_PN0P_  (.D(_02033_),
    .RN(net85),
    .CK(clknet_leaf_65_clk),
    .Q(\core.keymem.key_mem[4][24] ),
    .QN(_20571_));
 DFFR_X1 \core.keymem.key_mem[4][25]$_DFFE_PN0P_  (.D(_02034_),
    .RN(net85),
    .CK(clknet_leaf_48_clk),
    .Q(\core.keymem.key_mem[4][25] ),
    .QN(_20570_));
 DFFR_X1 \core.keymem.key_mem[4][26]$_DFFE_PN0P_  (.D(_02035_),
    .RN(net100),
    .CK(clknet_leaf_96_clk),
    .Q(\core.keymem.key_mem[4][26] ),
    .QN(_20569_));
 DFFR_X1 \core.keymem.key_mem[4][27]$_DFFE_PN0P_  (.D(_02036_),
    .RN(net16),
    .CK(clknet_leaf_151_clk),
    .Q(\core.keymem.key_mem[4][27] ),
    .QN(_20568_));
 DFFR_X1 \core.keymem.key_mem[4][28]$_DFFE_PN0P_  (.D(_02037_),
    .RN(net16),
    .CK(clknet_leaf_125_clk),
    .Q(\core.keymem.key_mem[4][28] ),
    .QN(_20567_));
 DFFR_X1 \core.keymem.key_mem[4][29]$_DFFE_PN0P_  (.D(_02038_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[4][29] ),
    .QN(_20566_));
 DFFR_X1 \core.keymem.key_mem[4][2]$_DFFE_PN0P_  (.D(_02039_),
    .RN(net89),
    .CK(clknet_leaf_65_clk),
    .Q(\core.keymem.key_mem[4][2] ),
    .QN(_20565_));
 DFFR_X1 \core.keymem.key_mem[4][30]$_DFFE_PN0P_  (.D(_02040_),
    .RN(net98),
    .CK(clknet_leaf_149_clk),
    .Q(\core.keymem.key_mem[4][30] ),
    .QN(_20564_));
 DFFR_X1 \core.keymem.key_mem[4][31]$_DFFE_PN0P_  (.D(_02041_),
    .RN(net98),
    .CK(clknet_leaf_143_clk),
    .Q(\core.keymem.key_mem[4][31] ),
    .QN(_20563_));
 DFFR_X1 \core.keymem.key_mem[4][32]$_DFFE_PN0P_  (.D(_02042_),
    .RN(net100),
    .CK(clknet_leaf_110_clk),
    .Q(\core.keymem.key_mem[4][32] ),
    .QN(_20562_));
 DFFR_X1 \core.keymem.key_mem[4][33]$_DFFE_PN0P_  (.D(_02043_),
    .RN(net16),
    .CK(clknet_leaf_126_clk),
    .Q(\core.keymem.key_mem[4][33] ),
    .QN(_20561_));
 DFFR_X1 \core.keymem.key_mem[4][34]$_DFFE_PN0P_  (.D(_02044_),
    .RN(net16),
    .CK(clknet_leaf_125_clk),
    .Q(\core.keymem.key_mem[4][34] ),
    .QN(_20560_));
 DFFR_X1 \core.keymem.key_mem[4][35]$_DFFE_PN0P_  (.D(_02045_),
    .RN(net99),
    .CK(clknet_leaf_127_clk),
    .Q(\core.keymem.key_mem[4][35] ),
    .QN(_20559_));
 DFFR_X1 \core.keymem.key_mem[4][36]$_DFFE_PN0P_  (.D(_02046_),
    .RN(net88),
    .CK(clknet_leaf_90_clk),
    .Q(\core.keymem.key_mem[4][36] ),
    .QN(_20558_));
 DFFR_X1 \core.keymem.key_mem[4][37]$_DFFE_PN0P_  (.D(_02047_),
    .RN(net89),
    .CK(clknet_leaf_85_clk),
    .Q(\core.keymem.key_mem[4][37] ),
    .QN(_20557_));
 DFFR_X1 \core.keymem.key_mem[4][38]$_DFFE_PN0P_  (.D(_02048_),
    .RN(net99),
    .CK(clknet_leaf_123_clk),
    .Q(\core.keymem.key_mem[4][38] ),
    .QN(_20556_));
 DFFR_X1 \core.keymem.key_mem[4][39]$_DFFE_PN0P_  (.D(_02049_),
    .RN(net85),
    .CK(clknet_leaf_87_clk),
    .Q(\core.keymem.key_mem[4][39] ),
    .QN(_20555_));
 DFFR_X1 \core.keymem.key_mem[4][3]$_DFFE_PN0P_  (.D(_02050_),
    .RN(net88),
    .CK(clknet_leaf_91_clk),
    .Q(\core.keymem.key_mem[4][3] ),
    .QN(_20554_));
 DFFR_X1 \core.keymem.key_mem[4][40]$_DFFE_PN0P_  (.D(_02051_),
    .RN(net88),
    .CK(clknet_leaf_90_clk),
    .Q(\core.keymem.key_mem[4][40] ),
    .QN(_20553_));
 DFFR_X1 \core.keymem.key_mem[4][41]$_DFFE_PN0P_  (.D(_02052_),
    .RN(net100),
    .CK(clknet_leaf_104_clk),
    .Q(\core.keymem.key_mem[4][41] ),
    .QN(_20552_));
 DFFR_X1 \core.keymem.key_mem[4][42]$_DFFE_PN0P_  (.D(_02053_),
    .RN(net100),
    .CK(clknet_leaf_129_clk),
    .Q(\core.keymem.key_mem[4][42] ),
    .QN(_20551_));
 DFFR_X1 \core.keymem.key_mem[4][43]$_DFFE_PN0P_  (.D(_02054_),
    .RN(net85),
    .CK(clknet_leaf_88_clk),
    .Q(\core.keymem.key_mem[4][43] ),
    .QN(_20550_));
 DFFR_X1 \core.keymem.key_mem[4][44]$_DFFE_PN0P_  (.D(_02055_),
    .RN(net100),
    .CK(clknet_leaf_113_clk),
    .Q(\core.keymem.key_mem[4][44] ),
    .QN(_20549_));
 DFFR_X1 \core.keymem.key_mem[4][45]$_DFFE_PN0P_  (.D(_02056_),
    .RN(net99),
    .CK(clknet_leaf_69_clk),
    .Q(\core.keymem.key_mem[4][45] ),
    .QN(_20548_));
 DFFR_X1 \core.keymem.key_mem[4][46]$_DFFE_PN0P_  (.D(_02057_),
    .RN(net99),
    .CK(clknet_leaf_80_clk),
    .Q(\core.keymem.key_mem[4][46] ),
    .QN(_20547_));
 DFFR_X1 \core.keymem.key_mem[4][47]$_DFFE_PN0P_  (.D(_02058_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[4][47] ),
    .QN(_20546_));
 DFFR_X1 \core.keymem.key_mem[4][48]$_DFFE_PN0P_  (.D(_02059_),
    .RN(net98),
    .CK(clknet_leaf_141_clk),
    .Q(\core.keymem.key_mem[4][48] ),
    .QN(_20545_));
 DFFR_X1 \core.keymem.key_mem[4][49]$_DFFE_PN0P_  (.D(_02060_),
    .RN(net99),
    .CK(clknet_leaf_78_clk),
    .Q(\core.keymem.key_mem[4][49] ),
    .QN(_20544_));
 DFFR_X1 \core.keymem.key_mem[4][4]$_DFFE_PN0P_  (.D(_02061_),
    .RN(net100),
    .CK(clknet_leaf_105_clk),
    .Q(\core.keymem.key_mem[4][4] ),
    .QN(_20543_));
 DFFR_X1 \core.keymem.key_mem[4][50]$_DFFE_PN0P_  (.D(_02062_),
    .RN(net98),
    .CK(clknet_leaf_140_clk),
    .Q(\core.keymem.key_mem[4][50] ),
    .QN(_20542_));
 DFFR_X1 \core.keymem.key_mem[4][51]$_DFFE_PN0P_  (.D(_02063_),
    .RN(net16),
    .CK(clknet_leaf_130_clk),
    .Q(\core.keymem.key_mem[4][51] ),
    .QN(_20541_));
 DFFR_X1 \core.keymem.key_mem[4][52]$_DFFE_PN0P_  (.D(_02064_),
    .RN(net99),
    .CK(clknet_leaf_81_clk),
    .Q(\core.keymem.key_mem[4][52] ),
    .QN(_20540_));
 DFFR_X1 \core.keymem.key_mem[4][53]$_DFFE_PN0P_  (.D(_02065_),
    .RN(net98),
    .CK(clknet_leaf_146_clk),
    .Q(\core.keymem.key_mem[4][53] ),
    .QN(_20539_));
 DFFR_X1 \core.keymem.key_mem[4][54]$_DFFE_PN0P_  (.D(_02066_),
    .RN(net98),
    .CK(clknet_leaf_145_clk),
    .Q(\core.keymem.key_mem[4][54] ),
    .QN(_20538_));
 DFFR_X1 \core.keymem.key_mem[4][55]$_DFFE_PN0P_  (.D(_02067_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[4][55] ),
    .QN(_20537_));
 DFFR_X1 \core.keymem.key_mem[4][56]$_DFFE_PN0P_  (.D(_02068_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[4][56] ),
    .QN(_20536_));
 DFFR_X1 \core.keymem.key_mem[4][57]$_DFFE_PN0P_  (.D(_02069_),
    .RN(net100),
    .CK(clknet_leaf_110_clk),
    .Q(\core.keymem.key_mem[4][57] ),
    .QN(_20535_));
 DFFR_X1 \core.keymem.key_mem[4][58]$_DFFE_PN0P_  (.D(_02070_),
    .RN(net100),
    .CK(clknet_leaf_106_clk),
    .Q(\core.keymem.key_mem[4][58] ),
    .QN(_20534_));
 DFFR_X1 \core.keymem.key_mem[4][59]$_DFFE_PN0P_  (.D(_02071_),
    .RN(net100),
    .CK(clknet_leaf_15_clk),
    .Q(\core.keymem.key_mem[4][59] ),
    .QN(_20533_));
 DFFR_X1 \core.keymem.key_mem[4][5]$_DFFE_PN0P_  (.D(_02072_),
    .RN(net100),
    .CK(clknet_leaf_19_clk),
    .Q(\core.keymem.key_mem[4][5] ),
    .QN(_20532_));
 DFFR_X1 \core.keymem.key_mem[4][60]$_DFFE_PN0P_  (.D(_02073_),
    .RN(net82),
    .CK(clknet_leaf_24_clk),
    .Q(\core.keymem.key_mem[4][60] ),
    .QN(_20531_));
 DFFR_X1 \core.keymem.key_mem[4][61]$_DFFE_PN0P_  (.D(_02074_),
    .RN(net89),
    .CK(clknet_leaf_104_clk),
    .Q(\core.keymem.key_mem[4][61] ),
    .QN(_20530_));
 DFFR_X1 \core.keymem.key_mem[4][62]$_DFFE_PN0P_  (.D(_02075_),
    .RN(net100),
    .CK(clknet_leaf_99_clk),
    .Q(\core.keymem.key_mem[4][62] ),
    .QN(_20529_));
 DFFR_X1 \core.keymem.key_mem[4][63]$_DFFE_PN0P_  (.D(_02076_),
    .RN(net100),
    .CK(clknet_leaf_95_clk),
    .Q(\core.keymem.key_mem[4][63] ),
    .QN(_20528_));
 DFFR_X1 \core.keymem.key_mem[4][64]$_DFFE_PN0P_  (.D(_02077_),
    .RN(net82),
    .CK(clknet_leaf_14_clk),
    .Q(\core.keymem.key_mem[4][64] ),
    .QN(_20527_));
 DFFR_X1 \core.keymem.key_mem[4][65]$_DFFE_PN0P_  (.D(_02078_),
    .RN(net98),
    .CK(clknet_leaf_140_clk),
    .Q(\core.keymem.key_mem[4][65] ),
    .QN(_20526_));
 DFFR_X1 \core.keymem.key_mem[4][66]$_DFFE_PN0P_  (.D(_02079_),
    .RN(net100),
    .CK(clknet_leaf_15_clk),
    .Q(\core.keymem.key_mem[4][66] ),
    .QN(_20525_));
 DFFR_X1 \core.keymem.key_mem[4][67]$_DFFE_PN0P_  (.D(_02080_),
    .RN(net95),
    .CK(clknet_leaf_77_clk),
    .Q(\core.keymem.key_mem[4][67] ),
    .QN(_20524_));
 DFFR_X1 \core.keymem.key_mem[4][68]$_DFFE_PN0P_  (.D(_02081_),
    .RN(net95),
    .CK(clknet_leaf_119_clk),
    .Q(\core.keymem.key_mem[4][68] ),
    .QN(_20523_));
 DFFR_X1 \core.keymem.key_mem[4][69]$_DFFE_PN0P_  (.D(_02082_),
    .RN(net98),
    .CK(clknet_leaf_176_clk),
    .Q(\core.keymem.key_mem[4][69] ),
    .QN(_20522_));
 DFFR_X1 \core.keymem.key_mem[4][6]$_DFFE_PN0P_  (.D(_02083_),
    .RN(net100),
    .CK(clknet_leaf_102_clk),
    .Q(\core.keymem.key_mem[4][6] ),
    .QN(_20521_));
 DFFR_X1 \core.keymem.key_mem[4][70]$_DFFE_PN0P_  (.D(_02084_),
    .RN(net100),
    .CK(clknet_leaf_100_clk),
    .Q(\core.keymem.key_mem[4][70] ),
    .QN(_20520_));
 DFFR_X1 \core.keymem.key_mem[4][71]$_DFFE_PN0P_  (.D(_02085_),
    .RN(net99),
    .CK(clknet_leaf_73_clk),
    .Q(\core.keymem.key_mem[4][71] ),
    .QN(_20519_));
 DFFR_X1 \core.keymem.key_mem[4][72]$_DFFE_PN0P_  (.D(_02086_),
    .RN(net95),
    .CK(clknet_leaf_179_clk),
    .Q(\core.keymem.key_mem[4][72] ),
    .QN(_20518_));
 DFFR_X1 \core.keymem.key_mem[4][73]$_DFFE_PN0P_  (.D(_02087_),
    .RN(net97),
    .CK(clknet_leaf_148_clk),
    .Q(\core.keymem.key_mem[4][73] ),
    .QN(_20517_));
 DFFR_X1 \core.keymem.key_mem[4][74]$_DFFE_PN0P_  (.D(_02088_),
    .RN(net97),
    .CK(clknet_leaf_157_clk),
    .Q(\core.keymem.key_mem[4][74] ),
    .QN(_20516_));
 DFFR_X1 \core.keymem.key_mem[4][75]$_DFFE_PN0P_  (.D(_02089_),
    .RN(net97),
    .CK(clknet_leaf_152_clk),
    .Q(\core.keymem.key_mem[4][75] ),
    .QN(_20515_));
 DFFR_X1 \core.keymem.key_mem[4][76]$_DFFE_PN0P_  (.D(_02090_),
    .RN(net93),
    .CK(clknet_leaf_376_clk),
    .Q(\core.keymem.key_mem[4][76] ),
    .QN(_20514_));
 DFFR_X1 \core.keymem.key_mem[4][77]$_DFFE_PN0P_  (.D(_02091_),
    .RN(net97),
    .CK(clknet_leaf_159_clk),
    .Q(\core.keymem.key_mem[4][77] ),
    .QN(_20513_));
 DFFR_X1 \core.keymem.key_mem[4][78]$_DFFE_PN0P_  (.D(_02092_),
    .RN(net96),
    .CK(clknet_leaf_172_clk),
    .Q(\core.keymem.key_mem[4][78] ),
    .QN(_20512_));
 DFFR_X1 \core.keymem.key_mem[4][79]$_DFFE_PN0P_  (.D(_02093_),
    .RN(net96),
    .CK(clknet_leaf_228_clk),
    .Q(\core.keymem.key_mem[4][79] ),
    .QN(_20511_));
 DFFR_X1 \core.keymem.key_mem[4][7]$_DFFE_PN0P_  (.D(_02094_),
    .RN(net98),
    .CK(clknet_leaf_172_clk),
    .Q(\core.keymem.key_mem[4][7] ),
    .QN(_20510_));
 DFFR_X1 \core.keymem.key_mem[4][80]$_DFFE_PN0P_  (.D(_02095_),
    .RN(net97),
    .CK(clknet_leaf_159_clk),
    .Q(\core.keymem.key_mem[4][80] ),
    .QN(_20509_));
 DFFR_X1 \core.keymem.key_mem[4][81]$_DFFE_PN0P_  (.D(_02096_),
    .RN(net97),
    .CK(clknet_leaf_157_clk),
    .Q(\core.keymem.key_mem[4][81] ),
    .QN(_20508_));
 DFFR_X1 \core.keymem.key_mem[4][82]$_DFFE_PN0P_  (.D(_02097_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[4][82] ),
    .QN(_20507_));
 DFFR_X1 \core.keymem.key_mem[4][83]$_DFFE_PN0P_  (.D(_02098_),
    .RN(net93),
    .CK(clknet_leaf_183_clk),
    .Q(\core.keymem.key_mem[4][83] ),
    .QN(_20506_));
 DFFR_X1 \core.keymem.key_mem[4][84]$_DFFE_PN0P_  (.D(_02099_),
    .RN(net95),
    .CK(clknet_leaf_182_clk),
    .Q(\core.keymem.key_mem[4][84] ),
    .QN(_20505_));
 DFFR_X1 \core.keymem.key_mem[4][85]$_DFFE_PN0P_  (.D(_02100_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[4][85] ),
    .QN(_20504_));
 DFFR_X1 \core.keymem.key_mem[4][86]$_DFFE_PN0P_  (.D(_02101_),
    .RN(net95),
    .CK(clknet_leaf_189_clk),
    .Q(\core.keymem.key_mem[4][86] ),
    .QN(_20503_));
 DFFR_X1 \core.keymem.key_mem[4][87]$_DFFE_PN0P_  (.D(_02102_),
    .RN(net89),
    .CK(clknet_leaf_56_clk),
    .Q(\core.keymem.key_mem[4][87] ),
    .QN(_20502_));
 DFFR_X1 \core.keymem.key_mem[4][88]$_DFFE_PN0P_  (.D(_02103_),
    .RN(net93),
    .CK(clknet_leaf_280_clk),
    .Q(\core.keymem.key_mem[4][88] ),
    .QN(_20501_));
 DFFR_X1 \core.keymem.key_mem[4][89]$_DFFE_PN0P_  (.D(_02104_),
    .RN(net93),
    .CK(clknet_leaf_199_clk),
    .Q(\core.keymem.key_mem[4][89] ),
    .QN(_20500_));
 DFFR_X1 \core.keymem.key_mem[4][8]$_DFFE_PN0P_  (.D(_02105_),
    .RN(net93),
    .CK(clknet_leaf_376_clk),
    .Q(\core.keymem.key_mem[4][8] ),
    .QN(_20499_));
 DFFR_X1 \core.keymem.key_mem[4][90]$_DFFE_PN0P_  (.D(_02106_),
    .RN(net97),
    .CK(clknet_leaf_161_clk),
    .Q(\core.keymem.key_mem[4][90] ),
    .QN(_20498_));
 DFFR_X1 \core.keymem.key_mem[4][91]$_DFFE_PN0P_  (.D(_02107_),
    .RN(net95),
    .CK(clknet_leaf_183_clk),
    .Q(\core.keymem.key_mem[4][91] ),
    .QN(_20497_));
 DFFR_X1 \core.keymem.key_mem[4][92]$_DFFE_PN0P_  (.D(_02108_),
    .RN(net95),
    .CK(clknet_leaf_63_clk),
    .Q(\core.keymem.key_mem[4][92] ),
    .QN(_20496_));
 DFFR_X1 \core.keymem.key_mem[4][93]$_DFFE_PN0P_  (.D(_02109_),
    .RN(net98),
    .CK(clknet_leaf_166_clk),
    .Q(\core.keymem.key_mem[4][93] ),
    .QN(_20495_));
 DFFR_X1 \core.keymem.key_mem[4][94]$_DFFE_PN0P_  (.D(_02110_),
    .RN(net96),
    .CK(clknet_leaf_226_clk),
    .Q(\core.keymem.key_mem[4][94] ),
    .QN(_20494_));
 DFFR_X1 \core.keymem.key_mem[4][95]$_DFFE_PN0P_  (.D(_02111_),
    .RN(net96),
    .CK(clknet_leaf_242_clk),
    .Q(\core.keymem.key_mem[4][95] ),
    .QN(_20493_));
 DFFR_X1 \core.keymem.key_mem[4][96]$_DFFE_PN0P_  (.D(_02112_),
    .RN(net92),
    .CK(clknet_leaf_266_clk),
    .Q(\core.keymem.key_mem[4][96] ),
    .QN(_20492_));
 DFFR_X1 \core.keymem.key_mem[4][97]$_DFFE_PN0P_  (.D(_02113_),
    .RN(net93),
    .CK(clknet_leaf_184_clk),
    .Q(\core.keymem.key_mem[4][97] ),
    .QN(_20491_));
 DFFR_X1 \core.keymem.key_mem[4][98]$_DFFE_PN0P_  (.D(_02114_),
    .RN(net95),
    .CK(clknet_leaf_195_clk),
    .Q(\core.keymem.key_mem[4][98] ),
    .QN(_20490_));
 DFFR_X1 \core.keymem.key_mem[4][99]$_DFFE_PN0P_  (.D(_02115_),
    .RN(net92),
    .CK(clknet_leaf_191_clk),
    .Q(\core.keymem.key_mem[4][99] ),
    .QN(_20489_));
 DFFR_X1 \core.keymem.key_mem[4][9]$_DFFE_PN0P_  (.D(_02116_),
    .RN(net92),
    .CK(clknet_leaf_205_clk),
    .Q(\core.keymem.key_mem[4][9] ),
    .QN(_20488_));
 DFFR_X1 \core.keymem.key_mem[5][0]$_DFFE_PN0P_  (.D(_02117_),
    .RN(net96),
    .CK(clknet_leaf_248_clk),
    .Q(\core.keymem.key_mem[5][0] ),
    .QN(_20487_));
 DFFR_X1 \core.keymem.key_mem[5][100]$_DFFE_PN0P_  (.D(_02118_),
    .RN(net94),
    .CK(clknet_leaf_211_clk),
    .Q(\core.keymem.key_mem[5][100] ),
    .QN(_20486_));
 DFFR_X1 \core.keymem.key_mem[5][101]$_DFFE_PN0P_  (.D(_02119_),
    .RN(net94),
    .CK(clknet_leaf_219_clk),
    .Q(\core.keymem.key_mem[5][101] ),
    .QN(_20485_));
 DFFR_X1 \core.keymem.key_mem[5][102]$_DFFE_PN0P_  (.D(_02120_),
    .RN(net96),
    .CK(clknet_leaf_232_clk),
    .Q(\core.keymem.key_mem[5][102] ),
    .QN(_20484_));
 DFFR_X1 \core.keymem.key_mem[5][103]$_DFFE_PN0P_  (.D(_02121_),
    .RN(net96),
    .CK(clknet_leaf_233_clk),
    .Q(\core.keymem.key_mem[5][103] ),
    .QN(_20483_));
 DFFR_X1 \core.keymem.key_mem[5][104]$_DFFE_PN0P_  (.D(_02122_),
    .RN(net93),
    .CK(clknet_leaf_190_clk),
    .Q(\core.keymem.key_mem[5][104] ),
    .QN(_20482_));
 DFFR_X1 \core.keymem.key_mem[5][105]$_DFFE_PN0P_  (.D(_02123_),
    .RN(net96),
    .CK(clknet_leaf_248_clk),
    .Q(\core.keymem.key_mem[5][105] ),
    .QN(_20481_));
 DFFR_X1 \core.keymem.key_mem[5][106]$_DFFE_PN0P_  (.D(_02124_),
    .RN(net92),
    .CK(clknet_leaf_267_clk),
    .Q(\core.keymem.key_mem[5][106] ),
    .QN(_20480_));
 DFFR_X1 \core.keymem.key_mem[5][107]$_DFFE_PN0P_  (.D(_02125_),
    .RN(net92),
    .CK(clknet_leaf_276_clk),
    .Q(\core.keymem.key_mem[5][107] ),
    .QN(_20479_));
 DFFR_X1 \core.keymem.key_mem[5][108]$_DFFE_PN0P_  (.D(_02126_),
    .RN(net92),
    .CK(clknet_leaf_277_clk),
    .Q(\core.keymem.key_mem[5][108] ),
    .QN(_20478_));
 DFFR_X1 \core.keymem.key_mem[5][109]$_DFFE_PN0P_  (.D(_02127_),
    .RN(net94),
    .CK(clknet_leaf_259_clk),
    .Q(\core.keymem.key_mem[5][109] ),
    .QN(_20477_));
 DFFR_X1 \core.keymem.key_mem[5][10]$_DFFE_PN0P_  (.D(_02128_),
    .RN(net95),
    .CK(clknet_leaf_190_clk),
    .Q(\core.keymem.key_mem[5][10] ),
    .QN(_20476_));
 DFFR_X1 \core.keymem.key_mem[5][110]$_DFFE_PN0P_  (.D(_02129_),
    .RN(net96),
    .CK(clknet_leaf_250_clk),
    .Q(\core.keymem.key_mem[5][110] ),
    .QN(_20475_));
 DFFR_X1 \core.keymem.key_mem[5][111]$_DFFE_PN0P_  (.D(_02130_),
    .RN(net96),
    .CK(clknet_leaf_226_clk),
    .Q(\core.keymem.key_mem[5][111] ),
    .QN(_20474_));
 DFFR_X1 \core.keymem.key_mem[5][112]$_DFFE_PN0P_  (.D(_02131_),
    .RN(net94),
    .CK(clknet_leaf_261_clk),
    .Q(\core.keymem.key_mem[5][112] ),
    .QN(_20473_));
 DFFR_X1 \core.keymem.key_mem[5][113]$_DFFE_PN0P_  (.D(_02132_),
    .RN(net92),
    .CK(clknet_leaf_273_clk),
    .Q(\core.keymem.key_mem[5][113] ),
    .QN(_20472_));
 DFFR_X1 \core.keymem.key_mem[5][114]$_DFFE_PN0P_  (.D(_02133_),
    .RN(net91),
    .CK(clknet_leaf_279_clk),
    .Q(\core.keymem.key_mem[5][114] ),
    .QN(_20471_));
 DFFR_X1 \core.keymem.key_mem[5][115]$_DFFE_PN0P_  (.D(_02134_),
    .RN(net92),
    .CK(clknet_leaf_272_clk),
    .Q(\core.keymem.key_mem[5][115] ),
    .QN(_20470_));
 DFFR_X1 \core.keymem.key_mem[5][116]$_DFFE_PN0P_  (.D(_02135_),
    .RN(net94),
    .CK(clknet_leaf_266_clk),
    .Q(\core.keymem.key_mem[5][116] ),
    .QN(_20469_));
 DFFR_X1 \core.keymem.key_mem[5][117]$_DFFE_PN0P_  (.D(_02136_),
    .RN(net96),
    .CK(clknet_leaf_223_clk),
    .Q(\core.keymem.key_mem[5][117] ),
    .QN(_20468_));
 DFFR_X1 \core.keymem.key_mem[5][118]$_DFFE_PN0P_  (.D(_02137_),
    .RN(net97),
    .CK(clknet_leaf_241_clk),
    .Q(\core.keymem.key_mem[5][118] ),
    .QN(_20467_));
 DFFR_X1 \core.keymem.key_mem[5][119]$_DFFE_PN0P_  (.D(_02138_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[5][119] ),
    .QN(_20466_));
 DFFR_X1 \core.keymem.key_mem[5][11]$_DFFE_PN0P_  (.D(_02139_),
    .RN(net95),
    .CK(clknet_leaf_61_clk),
    .Q(\core.keymem.key_mem[5][11] ),
    .QN(_20465_));
 DFFR_X1 \core.keymem.key_mem[5][120]$_DFFE_PN0P_  (.D(_02140_),
    .RN(net93),
    .CK(clknet_leaf_205_clk),
    .Q(\core.keymem.key_mem[5][120] ),
    .QN(_20464_));
 DFFR_X1 \core.keymem.key_mem[5][121]$_DFFE_PN0P_  (.D(_02141_),
    .RN(net94),
    .CK(clknet_leaf_216_clk),
    .Q(\core.keymem.key_mem[5][121] ),
    .QN(_20463_));
 DFFR_X1 \core.keymem.key_mem[5][122]$_DFFE_PN0P_  (.D(_02142_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[5][122] ),
    .QN(_20462_));
 DFFR_X1 \core.keymem.key_mem[5][123]$_DFFE_PN0P_  (.D(_02143_),
    .RN(net93),
    .CK(clknet_leaf_197_clk),
    .Q(\core.keymem.key_mem[5][123] ),
    .QN(_20461_));
 DFFR_X1 \core.keymem.key_mem[5][124]$_DFFE_PN0P_  (.D(_02144_),
    .RN(net93),
    .CK(clknet_leaf_198_clk),
    .Q(\core.keymem.key_mem[5][124] ),
    .QN(_20460_));
 DFFR_X1 \core.keymem.key_mem[5][125]$_DFFE_PN0P_  (.D(_02145_),
    .RN(net96),
    .CK(clknet_leaf_231_clk),
    .Q(\core.keymem.key_mem[5][125] ),
    .QN(_20459_));
 DFFR_X1 \core.keymem.key_mem[5][126]$_DFFE_PN0P_  (.D(_02146_),
    .RN(net94),
    .CK(clknet_leaf_188_clk),
    .Q(\core.keymem.key_mem[5][126] ),
    .QN(_20458_));
 DFFR_X1 \core.keymem.key_mem[5][127]$_DFFE_PN0P_  (.D(_02147_),
    .RN(net97),
    .CK(clknet_leaf_240_clk),
    .Q(\core.keymem.key_mem[5][127] ),
    .QN(_20457_));
 DFFR_X1 \core.keymem.key_mem[5][12]$_DFFE_PN0P_  (.D(_02148_),
    .RN(net93),
    .CK(clknet_leaf_206_clk),
    .Q(\core.keymem.key_mem[5][12] ),
    .QN(_20456_));
 DFFR_X1 \core.keymem.key_mem[5][13]$_DFFE_PN0P_  (.D(_02149_),
    .RN(net88),
    .CK(clknet_leaf_31_clk),
    .Q(\core.keymem.key_mem[5][13] ),
    .QN(_20455_));
 DFFR_X1 \core.keymem.key_mem[5][14]$_DFFE_PN0P_  (.D(_02150_),
    .RN(net94),
    .CK(clknet_leaf_209_clk),
    .Q(\core.keymem.key_mem[5][14] ),
    .QN(_20454_));
 DFFR_X1 \core.keymem.key_mem[5][15]$_DFFE_PN0P_  (.D(_02151_),
    .RN(net96),
    .CK(clknet_leaf_168_clk),
    .Q(\core.keymem.key_mem[5][15] ),
    .QN(_20453_));
 DFFR_X1 \core.keymem.key_mem[5][16]$_DFFE_PN0P_  (.D(_02152_),
    .RN(net89),
    .CK(clknet_leaf_32_clk),
    .Q(\core.keymem.key_mem[5][16] ),
    .QN(_20452_));
 DFFR_X1 \core.keymem.key_mem[5][17]$_DFFE_PN0P_  (.D(_02153_),
    .RN(net94),
    .CK(clknet_leaf_187_clk),
    .Q(\core.keymem.key_mem[5][17] ),
    .QN(_20451_));
 DFFR_X1 \core.keymem.key_mem[5][18]$_DFFE_PN0P_  (.D(_02154_),
    .RN(net82),
    .CK(clknet_leaf_34_clk),
    .Q(\core.keymem.key_mem[5][18] ),
    .QN(_20450_));
 DFFR_X1 \core.keymem.key_mem[5][19]$_DFFE_PN0P_  (.D(_02155_),
    .RN(net85),
    .CK(clknet_leaf_54_clk),
    .Q(\core.keymem.key_mem[5][19] ),
    .QN(_20449_));
 DFFR_X1 \core.keymem.key_mem[5][1]$_DFFE_PN0P_  (.D(_02156_),
    .RN(net89),
    .CK(clknet_leaf_22_clk),
    .Q(\core.keymem.key_mem[5][1] ),
    .QN(_20448_));
 DFFR_X1 \core.keymem.key_mem[5][20]$_DFFE_PN0P_  (.D(_02157_),
    .RN(net89),
    .CK(clknet_leaf_95_clk),
    .Q(\core.keymem.key_mem[5][20] ),
    .QN(_20447_));
 DFFR_X1 \core.keymem.key_mem[5][21]$_DFFE_PN0P_  (.D(_02158_),
    .RN(net89),
    .CK(clknet_leaf_66_clk),
    .Q(\core.keymem.key_mem[5][21] ),
    .QN(_20446_));
 DFFR_X1 \core.keymem.key_mem[5][22]$_DFFE_PN0P_  (.D(_02159_),
    .RN(net94),
    .CK(clknet_leaf_219_clk),
    .Q(\core.keymem.key_mem[5][22] ),
    .QN(_20445_));
 DFFR_X1 \core.keymem.key_mem[5][23]$_DFFE_PN0P_  (.D(_02160_),
    .RN(net89),
    .CK(clknet_leaf_55_clk),
    .Q(\core.keymem.key_mem[5][23] ),
    .QN(_20444_));
 DFFR_X1 \core.keymem.key_mem[5][24]$_DFFE_PN0P_  (.D(_02161_),
    .RN(net89),
    .CK(clknet_leaf_54_clk),
    .Q(\core.keymem.key_mem[5][24] ),
    .QN(_20443_));
 DFFR_X1 \core.keymem.key_mem[5][25]$_DFFE_PN0P_  (.D(_02162_),
    .RN(net85),
    .CK(clknet_leaf_48_clk),
    .Q(\core.keymem.key_mem[5][25] ),
    .QN(_20442_));
 DFFR_X1 \core.keymem.key_mem[5][26]$_DFFE_PN0P_  (.D(_02163_),
    .RN(net89),
    .CK(clknet_leaf_96_clk),
    .Q(\core.keymem.key_mem[5][26] ),
    .QN(_20441_));
 DFFR_X1 \core.keymem.key_mem[5][27]$_DFFE_PN0P_  (.D(_02164_),
    .RN(net16),
    .CK(clknet_leaf_151_clk),
    .Q(\core.keymem.key_mem[5][27] ),
    .QN(_20440_));
 DFFR_X1 \core.keymem.key_mem[5][28]$_DFFE_PN0P_  (.D(_02165_),
    .RN(net16),
    .CK(clknet_leaf_126_clk),
    .Q(\core.keymem.key_mem[5][28] ),
    .QN(_20439_));
 DFFR_X1 \core.keymem.key_mem[5][29]$_DFFE_PN0P_  (.D(_02166_),
    .RN(net16),
    .CK(clknet_leaf_132_clk),
    .Q(\core.keymem.key_mem[5][29] ),
    .QN(_20438_));
 DFFR_X1 \core.keymem.key_mem[5][2]$_DFFE_PN0P_  (.D(_02167_),
    .RN(net89),
    .CK(clknet_leaf_60_clk),
    .Q(\core.keymem.key_mem[5][2] ),
    .QN(_20437_));
 DFFR_X1 \core.keymem.key_mem[5][30]$_DFFE_PN0P_  (.D(_02168_),
    .RN(net98),
    .CK(clknet_leaf_149_clk),
    .Q(\core.keymem.key_mem[5][30] ),
    .QN(_20436_));
 DFFR_X1 \core.keymem.key_mem[5][31]$_DFFE_PN0P_  (.D(_02169_),
    .RN(net16),
    .CK(clknet_leaf_138_clk),
    .Q(\core.keymem.key_mem[5][31] ),
    .QN(_20435_));
 DFFR_X1 \core.keymem.key_mem[5][32]$_DFFE_PN0P_  (.D(_02170_),
    .RN(net100),
    .CK(clknet_leaf_110_clk),
    .Q(\core.keymem.key_mem[5][32] ),
    .QN(_20434_));
 DFFR_X1 \core.keymem.key_mem[5][33]$_DFFE_PN0P_  (.D(_02171_),
    .RN(net99),
    .CK(clknet_leaf_111_clk),
    .Q(\core.keymem.key_mem[5][33] ),
    .QN(_20433_));
 DFFR_X1 \core.keymem.key_mem[5][34]$_DFFE_PN0P_  (.D(_02172_),
    .RN(net16),
    .CK(clknet_leaf_124_clk),
    .Q(\core.keymem.key_mem[5][34] ),
    .QN(_20432_));
 DFFR_X1 \core.keymem.key_mem[5][35]$_DFFE_PN0P_  (.D(_02173_),
    .RN(net99),
    .CK(clknet_leaf_128_clk),
    .Q(\core.keymem.key_mem[5][35] ),
    .QN(_20431_));
 DFFR_X1 \core.keymem.key_mem[5][36]$_DFFE_PN0P_  (.D(_02174_),
    .RN(net88),
    .CK(clknet_leaf_91_clk),
    .Q(\core.keymem.key_mem[5][36] ),
    .QN(_20430_));
 DFFR_X1 \core.keymem.key_mem[5][37]$_DFFE_PN0P_  (.D(_02175_),
    .RN(net89),
    .CK(clknet_leaf_84_clk),
    .Q(\core.keymem.key_mem[5][37] ),
    .QN(_20429_));
 DFFR_X1 \core.keymem.key_mem[5][38]$_DFFE_PN0P_  (.D(_02176_),
    .RN(net16),
    .CK(clknet_leaf_123_clk),
    .Q(\core.keymem.key_mem[5][38] ),
    .QN(_20428_));
 DFFR_X1 \core.keymem.key_mem[5][39]$_DFFE_PN0P_  (.D(_02177_),
    .RN(net99),
    .CK(clknet_leaf_70_clk),
    .Q(\core.keymem.key_mem[5][39] ),
    .QN(_20427_));
 DFFR_X1 \core.keymem.key_mem[5][3]$_DFFE_PN0P_  (.D(_02178_),
    .RN(net85),
    .CK(clknet_leaf_47_clk),
    .Q(\core.keymem.key_mem[5][3] ),
    .QN(_20426_));
 DFFR_X1 \core.keymem.key_mem[5][40]$_DFFE_PN0P_  (.D(_02179_),
    .RN(net85),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[5][40] ),
    .QN(_20425_));
 DFFR_X1 \core.keymem.key_mem[5][41]$_DFFE_PN0P_  (.D(_02180_),
    .RN(net89),
    .CK(clknet_leaf_83_clk),
    .Q(\core.keymem.key_mem[5][41] ),
    .QN(_20424_));
 DFFR_X1 \core.keymem.key_mem[5][42]$_DFFE_PN0P_  (.D(_02181_),
    .RN(net100),
    .CK(clknet_leaf_109_clk),
    .Q(\core.keymem.key_mem[5][42] ),
    .QN(_20423_));
 DFFR_X1 \core.keymem.key_mem[5][43]$_DFFE_PN0P_  (.D(_02182_),
    .RN(net85),
    .CK(clknet_leaf_88_clk),
    .Q(\core.keymem.key_mem[5][43] ),
    .QN(_20422_));
 DFFR_X1 \core.keymem.key_mem[5][44]$_DFFE_PN0P_  (.D(_02183_),
    .RN(net100),
    .CK(clknet_leaf_107_clk),
    .Q(\core.keymem.key_mem[5][44] ),
    .QN(_20421_));
 DFFR_X1 \core.keymem.key_mem[5][45]$_DFFE_PN0P_  (.D(_02184_),
    .RN(net99),
    .CK(clknet_leaf_70_clk),
    .Q(\core.keymem.key_mem[5][45] ),
    .QN(_20420_));
 DFFR_X1 \core.keymem.key_mem[5][46]$_DFFE_PN0P_  (.D(_02185_),
    .RN(net99),
    .CK(clknet_leaf_82_clk),
    .Q(\core.keymem.key_mem[5][46] ),
    .QN(_20419_));
 DFFR_X1 \core.keymem.key_mem[5][47]$_DFFE_PN0P_  (.D(_02186_),
    .RN(net98),
    .CK(clknet_leaf_175_clk),
    .Q(\core.keymem.key_mem[5][47] ),
    .QN(_20418_));
 DFFR_X1 \core.keymem.key_mem[5][48]$_DFFE_PN0P_  (.D(_02187_),
    .RN(net99),
    .CK(clknet_leaf_119_clk),
    .Q(\core.keymem.key_mem[5][48] ),
    .QN(_20417_));
 DFFR_X1 \core.keymem.key_mem[5][49]$_DFFE_PN0P_  (.D(_02188_),
    .RN(net99),
    .CK(clknet_leaf_118_clk),
    .Q(\core.keymem.key_mem[5][49] ),
    .QN(_20416_));
 DFFR_X1 \core.keymem.key_mem[5][4]$_DFFE_PN0P_  (.D(_02189_),
    .RN(net100),
    .CK(clknet_leaf_105_clk),
    .Q(\core.keymem.key_mem[5][4] ),
    .QN(_20415_));
 DFFR_X1 \core.keymem.key_mem[5][50]$_DFFE_PN0P_  (.D(_02190_),
    .RN(net98),
    .CK(clknet_leaf_137_clk),
    .Q(\core.keymem.key_mem[5][50] ),
    .QN(_20414_));
 DFFR_X1 \core.keymem.key_mem[5][51]$_DFFE_PN0P_  (.D(_02191_),
    .RN(net100),
    .CK(clknet_leaf_130_clk),
    .Q(\core.keymem.key_mem[5][51] ),
    .QN(_20413_));
 DFFR_X1 \core.keymem.key_mem[5][52]$_DFFE_PN0P_  (.D(_02192_),
    .RN(net99),
    .CK(clknet_leaf_81_clk),
    .Q(\core.keymem.key_mem[5][52] ),
    .QN(_20412_));
 DFFR_X1 \core.keymem.key_mem[5][53]$_DFFE_PN0P_  (.D(_02193_),
    .RN(net98),
    .CK(clknet_leaf_176_clk),
    .Q(\core.keymem.key_mem[5][53] ),
    .QN(_20411_));
 DFFR_X1 \core.keymem.key_mem[5][54]$_DFFE_PN0P_  (.D(_02194_),
    .RN(net98),
    .CK(clknet_leaf_141_clk),
    .Q(\core.keymem.key_mem[5][54] ),
    .QN(_20410_));
 DFFR_X1 \core.keymem.key_mem[5][55]$_DFFE_PN0P_  (.D(_02195_),
    .RN(net16),
    .CK(clknet_leaf_135_clk),
    .Q(\core.keymem.key_mem[5][55] ),
    .QN(_20409_));
 DFFR_X1 \core.keymem.key_mem[5][56]$_DFFE_PN0P_  (.D(_02196_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[5][56] ),
    .QN(_20408_));
 DFFR_X1 \core.keymem.key_mem[5][57]$_DFFE_PN0P_  (.D(_02197_),
    .RN(net100),
    .CK(clknet_leaf_108_clk),
    .Q(\core.keymem.key_mem[5][57] ),
    .QN(_20407_));
 DFFR_X1 \core.keymem.key_mem[5][58]$_DFFE_PN0P_  (.D(_02198_),
    .RN(net100),
    .CK(clknet_leaf_102_clk),
    .Q(\core.keymem.key_mem[5][58] ),
    .QN(_20406_));
 DFFR_X1 \core.keymem.key_mem[5][59]$_DFFE_PN0P_  (.D(_02199_),
    .RN(net82),
    .CK(clknet_leaf_23_clk),
    .Q(\core.keymem.key_mem[5][59] ),
    .QN(_20405_));
 DFFR_X1 \core.keymem.key_mem[5][5]$_DFFE_PN0P_  (.D(_02200_),
    .RN(net100),
    .CK(clknet_leaf_19_clk),
    .Q(\core.keymem.key_mem[5][5] ),
    .QN(_20404_));
 DFFR_X1 \core.keymem.key_mem[5][60]$_DFFE_PN0P_  (.D(_02201_),
    .RN(net82),
    .CK(clknet_leaf_13_clk),
    .Q(\core.keymem.key_mem[5][60] ),
    .QN(_20403_));
 DFFR_X1 \core.keymem.key_mem[5][61]$_DFFE_PN0P_  (.D(_02202_),
    .RN(net89),
    .CK(clknet_leaf_104_clk),
    .Q(\core.keymem.key_mem[5][61] ),
    .QN(_20402_));
 DFFR_X1 \core.keymem.key_mem[5][62]$_DFFE_PN0P_  (.D(_02203_),
    .RN(net100),
    .CK(clknet_leaf_99_clk),
    .Q(\core.keymem.key_mem[5][62] ),
    .QN(_20401_));
 DFFR_X1 \core.keymem.key_mem[5][63]$_DFFE_PN0P_  (.D(_02204_),
    .RN(net100),
    .CK(clknet_leaf_98_clk),
    .Q(\core.keymem.key_mem[5][63] ),
    .QN(_20400_));
 DFFR_X1 \core.keymem.key_mem[5][64]$_DFFE_PN0P_  (.D(_02205_),
    .RN(net82),
    .CK(clknet_leaf_13_clk),
    .Q(\core.keymem.key_mem[5][64] ),
    .QN(_20399_));
 DFFR_X1 \core.keymem.key_mem[5][65]$_DFFE_PN0P_  (.D(_02206_),
    .RN(net99),
    .CK(clknet_leaf_120_clk),
    .Q(\core.keymem.key_mem[5][65] ),
    .QN(_20398_));
 DFFR_X1 \core.keymem.key_mem[5][66]$_DFFE_PN0P_  (.D(_02207_),
    .RN(net100),
    .CK(clknet_leaf_17_clk),
    .Q(\core.keymem.key_mem[5][66] ),
    .QN(_20397_));
 DFFR_X1 \core.keymem.key_mem[5][67]$_DFFE_PN0P_  (.D(_02208_),
    .RN(net95),
    .CK(clknet_leaf_76_clk),
    .Q(\core.keymem.key_mem[5][67] ),
    .QN(_20396_));
 DFFR_X1 \core.keymem.key_mem[5][68]$_DFFE_PN0P_  (.D(_02209_),
    .RN(net99),
    .CK(clknet_leaf_117_clk),
    .Q(\core.keymem.key_mem[5][68] ),
    .QN(_20395_));
 DFFR_X1 \core.keymem.key_mem[5][69]$_DFFE_PN0P_  (.D(_02210_),
    .RN(net98),
    .CK(clknet_leaf_142_clk),
    .Q(\core.keymem.key_mem[5][69] ),
    .QN(_20394_));
 DFFR_X1 \core.keymem.key_mem[5][6]$_DFFE_PN0P_  (.D(_02211_),
    .RN(net100),
    .CK(clknet_leaf_103_clk),
    .Q(\core.keymem.key_mem[5][6] ),
    .QN(_20393_));
 DFFR_X1 \core.keymem.key_mem[5][70]$_DFFE_PN0P_  (.D(_02212_),
    .RN(net100),
    .CK(clknet_leaf_101_clk),
    .Q(\core.keymem.key_mem[5][70] ),
    .QN(_20392_));
 DFFR_X1 \core.keymem.key_mem[5][71]$_DFFE_PN0P_  (.D(_02213_),
    .RN(net99),
    .CK(clknet_leaf_74_clk),
    .Q(\core.keymem.key_mem[5][71] ),
    .QN(_20391_));
 DFFR_X1 \core.keymem.key_mem[5][72]$_DFFE_PN0P_  (.D(_02214_),
    .RN(net95),
    .CK(clknet_leaf_76_clk),
    .Q(\core.keymem.key_mem[5][72] ),
    .QN(_20390_));
 DFFR_X1 \core.keymem.key_mem[5][73]$_DFFE_PN0P_  (.D(_02215_),
    .RN(net97),
    .CK(clknet_leaf_147_clk),
    .Q(\core.keymem.key_mem[5][73] ),
    .QN(_20389_));
 DFFR_X1 \core.keymem.key_mem[5][74]$_DFFE_PN0P_  (.D(_02216_),
    .RN(net97),
    .CK(clknet_leaf_156_clk),
    .Q(\core.keymem.key_mem[5][74] ),
    .QN(_20388_));
 DFFR_X1 \core.keymem.key_mem[5][75]$_DFFE_PN0P_  (.D(_02217_),
    .RN(net97),
    .CK(clknet_leaf_154_clk),
    .Q(\core.keymem.key_mem[5][75] ),
    .QN(_20387_));
 DFFR_X1 \core.keymem.key_mem[5][76]$_DFFE_PN0P_  (.D(_02218_),
    .RN(net93),
    .CK(clknet_leaf_283_clk),
    .Q(\core.keymem.key_mem[5][76] ),
    .QN(_20386_));
 DFFR_X1 \core.keymem.key_mem[5][77]$_DFFE_PN0P_  (.D(_02219_),
    .RN(net97),
    .CK(clknet_leaf_160_clk),
    .Q(\core.keymem.key_mem[5][77] ),
    .QN(_20385_));
 DFFR_X1 \core.keymem.key_mem[5][78]$_DFFE_PN0P_  (.D(_02220_),
    .RN(net97),
    .CK(clknet_leaf_164_clk),
    .Q(\core.keymem.key_mem[5][78] ),
    .QN(_20384_));
 DFFR_X1 \core.keymem.key_mem[5][79]$_DFFE_PN0P_  (.D(_02221_),
    .RN(net98),
    .CK(clknet_leaf_229_clk),
    .Q(\core.keymem.key_mem[5][79] ),
    .QN(_20383_));
 DFFR_X1 \core.keymem.key_mem[5][7]$_DFFE_PN0P_  (.D(_02222_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[5][7] ),
    .QN(_20382_));
 DFFR_X1 \core.keymem.key_mem[5][80]$_DFFE_PN0P_  (.D(_02223_),
    .RN(net97),
    .CK(clknet_leaf_158_clk),
    .Q(\core.keymem.key_mem[5][80] ),
    .QN(_20381_));
 DFFR_X1 \core.keymem.key_mem[5][81]$_DFFE_PN0P_  (.D(_02224_),
    .RN(net97),
    .CK(clknet_leaf_153_clk),
    .Q(\core.keymem.key_mem[5][81] ),
    .QN(_20380_));
 DFFR_X1 \core.keymem.key_mem[5][82]$_DFFE_PN0P_  (.D(_02225_),
    .RN(net98),
    .CK(clknet_leaf_186_clk),
    .Q(\core.keymem.key_mem[5][82] ),
    .QN(_20379_));
 DFFR_X1 \core.keymem.key_mem[5][83]$_DFFE_PN0P_  (.D(_02226_),
    .RN(net95),
    .CK(clknet_leaf_185_clk),
    .Q(\core.keymem.key_mem[5][83] ),
    .QN(_20378_));
 DFFR_X1 \core.keymem.key_mem[5][84]$_DFFE_PN0P_  (.D(_02227_),
    .RN(net95),
    .CK(clknet_leaf_181_clk),
    .Q(\core.keymem.key_mem[5][84] ),
    .QN(_20377_));
 DFFR_X1 \core.keymem.key_mem[5][85]$_DFFE_PN0P_  (.D(_02228_),
    .RN(net97),
    .CK(clknet_leaf_236_clk),
    .Q(\core.keymem.key_mem[5][85] ),
    .QN(_20376_));
 DFFR_X1 \core.keymem.key_mem[5][86]$_DFFE_PN0P_  (.D(_02229_),
    .RN(net95),
    .CK(clknet_leaf_191_clk),
    .Q(\core.keymem.key_mem[5][86] ),
    .QN(_20375_));
 DFFR_X1 \core.keymem.key_mem[5][87]$_DFFE_PN0P_  (.D(_02230_),
    .RN(net89),
    .CK(clknet_leaf_56_clk),
    .Q(\core.keymem.key_mem[5][87] ),
    .QN(_20374_));
 DFFR_X1 \core.keymem.key_mem[5][88]$_DFFE_PN0P_  (.D(_02231_),
    .RN(net91),
    .CK(clknet_leaf_280_clk),
    .Q(\core.keymem.key_mem[5][88] ),
    .QN(_20373_));
 DFFR_X1 \core.keymem.key_mem[5][89]$_DFFE_PN0P_  (.D(_02232_),
    .RN(net93),
    .CK(clknet_leaf_200_clk),
    .Q(\core.keymem.key_mem[5][89] ),
    .QN(_20372_));
 DFFR_X1 \core.keymem.key_mem[5][8]$_DFFE_PN0P_  (.D(_02233_),
    .RN(net93),
    .CK(clknet_leaf_377_clk),
    .Q(\core.keymem.key_mem[5][8] ),
    .QN(_20371_));
 DFFR_X1 \core.keymem.key_mem[5][90]$_DFFE_PN0P_  (.D(_02234_),
    .RN(net97),
    .CK(clknet_leaf_163_clk),
    .Q(\core.keymem.key_mem[5][90] ),
    .QN(_20370_));
 DFFR_X1 \core.keymem.key_mem[5][91]$_DFFE_PN0P_  (.D(_02235_),
    .RN(net95),
    .CK(clknet_leaf_181_clk),
    .Q(\core.keymem.key_mem[5][91] ),
    .QN(_20369_));
 DFFR_X1 \core.keymem.key_mem[5][92]$_DFFE_PN0P_  (.D(_02236_),
    .RN(net95),
    .CK(clknet_leaf_71_clk),
    .Q(\core.keymem.key_mem[5][92] ),
    .QN(_20368_));
 DFFR_X1 \core.keymem.key_mem[5][93]$_DFFE_PN0P_  (.D(_02237_),
    .RN(net97),
    .CK(clknet_leaf_162_clk),
    .Q(\core.keymem.key_mem[5][93] ),
    .QN(_20367_));
 DFFR_X1 \core.keymem.key_mem[5][94]$_DFFE_PN0P_  (.D(_02238_),
    .RN(net94),
    .CK(clknet_leaf_213_clk),
    .Q(\core.keymem.key_mem[5][94] ),
    .QN(_20366_));
 DFFR_X1 \core.keymem.key_mem[5][95]$_DFFE_PN0P_  (.D(_02239_),
    .RN(net96),
    .CK(clknet_leaf_242_clk),
    .Q(\core.keymem.key_mem[5][95] ),
    .QN(_20365_));
 DFFR_X1 \core.keymem.key_mem[5][96]$_DFFE_PN0P_  (.D(_02240_),
    .RN(net92),
    .CK(clknet_leaf_204_clk),
    .Q(\core.keymem.key_mem[5][96] ),
    .QN(_20364_));
 DFFR_X1 \core.keymem.key_mem[5][97]$_DFFE_PN0P_  (.D(_02241_),
    .RN(net93),
    .CK(clknet_leaf_194_clk),
    .Q(\core.keymem.key_mem[5][97] ),
    .QN(_20363_));
 DFFR_X1 \core.keymem.key_mem[5][98]$_DFFE_PN0P_  (.D(_02242_),
    .RN(net93),
    .CK(clknet_leaf_195_clk),
    .Q(\core.keymem.key_mem[5][98] ),
    .QN(_20362_));
 DFFR_X1 \core.keymem.key_mem[5][99]$_DFFE_PN0P_  (.D(_02243_),
    .RN(net92),
    .CK(clknet_leaf_201_clk),
    .Q(\core.keymem.key_mem[5][99] ),
    .QN(_20361_));
 DFFR_X1 \core.keymem.key_mem[5][9]$_DFFE_PN0P_  (.D(_02244_),
    .RN(net92),
    .CK(clknet_leaf_203_clk),
    .Q(\core.keymem.key_mem[5][9] ),
    .QN(_20360_));
 DFFR_X1 \core.keymem.key_mem[6][0]$_DFFE_PN0P_  (.D(_02245_),
    .RN(net96),
    .CK(clknet_leaf_247_clk),
    .Q(\core.keymem.key_mem[6][0] ),
    .QN(_20359_));
 DFFR_X1 \core.keymem.key_mem[6][100]$_DFFE_PN0P_  (.D(_02246_),
    .RN(net98),
    .CK(clknet_leaf_210_clk),
    .Q(\core.keymem.key_mem[6][100] ),
    .QN(_20358_));
 DFFR_X1 \core.keymem.key_mem[6][101]$_DFFE_PN0P_  (.D(_02247_),
    .RN(net96),
    .CK(clknet_leaf_245_clk),
    .Q(\core.keymem.key_mem[6][101] ),
    .QN(_20357_));
 DFFR_X1 \core.keymem.key_mem[6][102]$_DFFE_PN0P_  (.D(_02248_),
    .RN(net96),
    .CK(clknet_leaf_233_clk),
    .Q(\core.keymem.key_mem[6][102] ),
    .QN(_20356_));
 DFFR_X1 \core.keymem.key_mem[6][103]$_DFFE_PN0P_  (.D(_02249_),
    .RN(net96),
    .CK(clknet_leaf_223_clk),
    .Q(\core.keymem.key_mem[6][103] ),
    .QN(_20355_));
 DFFR_X1 \core.keymem.key_mem[6][104]$_DFFE_PN0P_  (.D(_02250_),
    .RN(net93),
    .CK(clknet_leaf_192_clk),
    .Q(\core.keymem.key_mem[6][104] ),
    .QN(_20354_));
 DFFR_X1 \core.keymem.key_mem[6][105]$_DFFE_PN0P_  (.D(_02251_),
    .RN(net96),
    .CK(clknet_leaf_247_clk),
    .Q(\core.keymem.key_mem[6][105] ),
    .QN(_20353_));
 DFFR_X1 \core.keymem.key_mem[6][106]$_DFFE_PN0P_  (.D(_02252_),
    .RN(net92),
    .CK(clknet_leaf_269_clk),
    .Q(\core.keymem.key_mem[6][106] ),
    .QN(_20352_));
 DFFR_X1 \core.keymem.key_mem[6][107]$_DFFE_PN0P_  (.D(_02253_),
    .RN(net92),
    .CK(clknet_leaf_267_clk),
    .Q(\core.keymem.key_mem[6][107] ),
    .QN(_20351_));
 DFFR_X1 \core.keymem.key_mem[6][108]$_DFFE_PN0P_  (.D(_02254_),
    .RN(net92),
    .CK(clknet_leaf_277_clk),
    .Q(\core.keymem.key_mem[6][108] ),
    .QN(_20350_));
 DFFR_X1 \core.keymem.key_mem[6][109]$_DFFE_PN0P_  (.D(_02255_),
    .RN(net94),
    .CK(clknet_leaf_259_clk),
    .Q(\core.keymem.key_mem[6][109] ),
    .QN(_20349_));
 DFFR_X1 \core.keymem.key_mem[6][10]$_DFFE_PN0P_  (.D(_02256_),
    .RN(net95),
    .CK(clknet_leaf_190_clk),
    .Q(\core.keymem.key_mem[6][10] ),
    .QN(_20348_));
 DFFR_X1 \core.keymem.key_mem[6][110]$_DFFE_PN0P_  (.D(_02257_),
    .RN(net96),
    .CK(clknet_leaf_250_clk),
    .Q(\core.keymem.key_mem[6][110] ),
    .QN(_20347_));
 DFFR_X1 \core.keymem.key_mem[6][111]$_DFFE_PN0P_  (.D(_02258_),
    .RN(net96),
    .CK(clknet_leaf_227_clk),
    .Q(\core.keymem.key_mem[6][111] ),
    .QN(_20346_));
 DFFR_X1 \core.keymem.key_mem[6][112]$_DFFE_PN0P_  (.D(_02259_),
    .RN(net94),
    .CK(clknet_leaf_261_clk),
    .Q(\core.keymem.key_mem[6][112] ),
    .QN(_20345_));
 DFFR_X1 \core.keymem.key_mem[6][113]$_DFFE_PN0P_  (.D(_02260_),
    .RN(net92),
    .CK(clknet_leaf_272_clk),
    .Q(\core.keymem.key_mem[6][113] ),
    .QN(_20344_));
 DFFR_X1 \core.keymem.key_mem[6][114]$_DFFE_PN0P_  (.D(_02261_),
    .RN(net91),
    .CK(clknet_leaf_278_clk),
    .Q(\core.keymem.key_mem[6][114] ),
    .QN(_20343_));
 DFFR_X1 \core.keymem.key_mem[6][115]$_DFFE_PN0P_  (.D(_02262_),
    .RN(net92),
    .CK(clknet_leaf_272_clk),
    .Q(\core.keymem.key_mem[6][115] ),
    .QN(_20342_));
 DFFR_X1 \core.keymem.key_mem[6][116]$_DFFE_PN0P_  (.D(_02263_),
    .RN(net94),
    .CK(clknet_leaf_265_clk),
    .Q(\core.keymem.key_mem[6][116] ),
    .QN(_20341_));
 DFFR_X1 \core.keymem.key_mem[6][117]$_DFFE_PN0P_  (.D(_02264_),
    .RN(net96),
    .CK(clknet_leaf_222_clk),
    .Q(\core.keymem.key_mem[6][117] ),
    .QN(_20340_));
 DFFR_X1 \core.keymem.key_mem[6][118]$_DFFE_PN0P_  (.D(_02265_),
    .RN(net96),
    .CK(clknet_leaf_243_clk),
    .Q(\core.keymem.key_mem[6][118] ),
    .QN(_20339_));
 DFFR_X1 \core.keymem.key_mem[6][119]$_DFFE_PN0P_  (.D(_02266_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[6][119] ),
    .QN(_20338_));
 DFFR_X1 \core.keymem.key_mem[6][11]$_DFFE_PN0P_  (.D(_02267_),
    .RN(net95),
    .CK(clknet_leaf_60_clk),
    .Q(\core.keymem.key_mem[6][11] ),
    .QN(_20337_));
 DFFR_X1 \core.keymem.key_mem[6][120]$_DFFE_PN0P_  (.D(_02268_),
    .RN(net94),
    .CK(clknet_leaf_215_clk),
    .Q(\core.keymem.key_mem[6][120] ),
    .QN(_20336_));
 DFFR_X1 \core.keymem.key_mem[6][121]$_DFFE_PN0P_  (.D(_02269_),
    .RN(net94),
    .CK(clknet_leaf_265_clk),
    .Q(\core.keymem.key_mem[6][121] ),
    .QN(_20335_));
 DFFR_X1 \core.keymem.key_mem[6][122]$_DFFE_PN0P_  (.D(_02270_),
    .RN(net97),
    .CK(clknet_leaf_237_clk),
    .Q(\core.keymem.key_mem[6][122] ),
    .QN(_20334_));
 DFFR_X1 \core.keymem.key_mem[6][123]$_DFFE_PN0P_  (.D(_02271_),
    .RN(net93),
    .CK(clknet_leaf_196_clk),
    .Q(\core.keymem.key_mem[6][123] ),
    .QN(_20333_));
 DFFR_X1 \core.keymem.key_mem[6][124]$_DFFE_PN0P_  (.D(_02272_),
    .RN(net93),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[6][124] ),
    .QN(_20332_));
 DFFR_X1 \core.keymem.key_mem[6][125]$_DFFE_PN0P_  (.D(_02273_),
    .RN(net97),
    .CK(clknet_leaf_235_clk),
    .Q(\core.keymem.key_mem[6][125] ),
    .QN(_20331_));
 DFFR_X1 \core.keymem.key_mem[6][126]$_DFFE_PN0P_  (.D(_02274_),
    .RN(net98),
    .CK(clknet_leaf_167_clk),
    .Q(\core.keymem.key_mem[6][126] ),
    .QN(_20330_));
 DFFR_X1 \core.keymem.key_mem[6][127]$_DFFE_PN0P_  (.D(_02275_),
    .RN(net97),
    .CK(clknet_leaf_243_clk),
    .Q(\core.keymem.key_mem[6][127] ),
    .QN(_20329_));
 DFFR_X1 \core.keymem.key_mem[6][12]$_DFFE_PN0P_  (.D(_02276_),
    .RN(net93),
    .CK(clknet_leaf_206_clk),
    .Q(\core.keymem.key_mem[6][12] ),
    .QN(_20328_));
 DFFR_X1 \core.keymem.key_mem[6][13]$_DFFE_PN0P_  (.D(_02277_),
    .RN(net88),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[6][13] ),
    .QN(_20327_));
 DFFR_X1 \core.keymem.key_mem[6][14]$_DFFE_PN0P_  (.D(_02278_),
    .RN(net98),
    .CK(clknet_leaf_229_clk),
    .Q(\core.keymem.key_mem[6][14] ),
    .QN(_20326_));
 DFFR_X1 \core.keymem.key_mem[6][15]$_DFFE_PN0P_  (.D(_02279_),
    .RN(net96),
    .CK(clknet_leaf_171_clk),
    .Q(\core.keymem.key_mem[6][15] ),
    .QN(_20325_));
 DFFR_X1 \core.keymem.key_mem[6][16]$_DFFE_PN0P_  (.D(_02280_),
    .RN(net89),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[6][16] ),
    .QN(_20324_));
 DFFR_X1 \core.keymem.key_mem[6][17]$_DFFE_PN0P_  (.D(_02281_),
    .RN(net98),
    .CK(clknet_leaf_168_clk),
    .Q(\core.keymem.key_mem[6][17] ),
    .QN(_20323_));
 DFFR_X1 \core.keymem.key_mem[6][18]$_DFFE_PN0P_  (.D(_02282_),
    .RN(net89),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[6][18] ),
    .QN(_20322_));
 DFFR_X1 \core.keymem.key_mem[6][19]$_DFFE_PN0P_  (.D(_02283_),
    .RN(net89),
    .CK(clknet_leaf_64_clk),
    .Q(\core.keymem.key_mem[6][19] ),
    .QN(_20321_));
 DFFR_X1 \core.keymem.key_mem[6][1]$_DFFE_PN0P_  (.D(_02284_),
    .RN(net89),
    .CK(clknet_leaf_27_clk),
    .Q(\core.keymem.key_mem[6][1] ),
    .QN(_20320_));
 DFFR_X1 \core.keymem.key_mem[6][20]$_DFFE_PN0P_  (.D(_02285_),
    .RN(net89),
    .CK(clknet_leaf_93_clk),
    .Q(\core.keymem.key_mem[6][20] ),
    .QN(_20319_));
 DFFR_X1 \core.keymem.key_mem[6][21]$_DFFE_PN0P_  (.D(_02286_),
    .RN(net89),
    .CK(clknet_leaf_69_clk),
    .Q(\core.keymem.key_mem[6][21] ),
    .QN(_20318_));
 DFFR_X1 \core.keymem.key_mem[6][22]$_DFFE_PN0P_  (.D(_02287_),
    .RN(net96),
    .CK(clknet_leaf_221_clk),
    .Q(\core.keymem.key_mem[6][22] ),
    .QN(_20317_));
 DFFR_X1 \core.keymem.key_mem[6][23]$_DFFE_PN0P_  (.D(_02288_),
    .RN(net89),
    .CK(clknet_leaf_54_clk),
    .Q(\core.keymem.key_mem[6][23] ),
    .QN(_20316_));
 DFFR_X1 \core.keymem.key_mem[6][24]$_DFFE_PN0P_  (.D(_02289_),
    .RN(net85),
    .CK(clknet_leaf_49_clk),
    .Q(\core.keymem.key_mem[6][24] ),
    .QN(_20315_));
 DFFR_X1 \core.keymem.key_mem[6][25]$_DFFE_PN0P_  (.D(_02290_),
    .RN(net85),
    .CK(clknet_leaf_47_clk),
    .Q(\core.keymem.key_mem[6][25] ),
    .QN(_20314_));
 DFFR_X1 \core.keymem.key_mem[6][26]$_DFFE_PN0P_  (.D(_02291_),
    .RN(net89),
    .CK(clknet_leaf_27_clk),
    .Q(\core.keymem.key_mem[6][26] ),
    .QN(_20313_));
 DFFR_X1 \core.keymem.key_mem[6][27]$_DFFE_PN0P_  (.D(_02292_),
    .RN(net16),
    .CK(clknet_leaf_132_clk),
    .Q(\core.keymem.key_mem[6][27] ),
    .QN(_20312_));
 DFFR_X1 \core.keymem.key_mem[6][28]$_DFFE_PN0P_  (.D(_02293_),
    .RN(net16),
    .CK(clknet_leaf_126_clk),
    .Q(\core.keymem.key_mem[6][28] ),
    .QN(_20311_));
 DFFR_X1 \core.keymem.key_mem[6][29]$_DFFE_PN0P_  (.D(_02294_),
    .RN(net16),
    .CK(clknet_leaf_132_clk),
    .Q(\core.keymem.key_mem[6][29] ),
    .QN(_20310_));
 DFFR_X1 \core.keymem.key_mem[6][2]$_DFFE_PN0P_  (.D(_02295_),
    .RN(net89),
    .CK(clknet_leaf_64_clk),
    .Q(\core.keymem.key_mem[6][2] ),
    .QN(_20309_));
 DFFR_X1 \core.keymem.key_mem[6][30]$_DFFE_PN0P_  (.D(_02296_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[6][30] ),
    .QN(_20308_));
 DFFR_X1 \core.keymem.key_mem[6][31]$_DFFE_PN0P_  (.D(_02297_),
    .RN(net16),
    .CK(clknet_leaf_137_clk),
    .Q(\core.keymem.key_mem[6][31] ),
    .QN(_20307_));
 DFFR_X1 \core.keymem.key_mem[6][32]$_DFFE_PN0P_  (.D(_02298_),
    .RN(net99),
    .CK(clknet_leaf_112_clk),
    .Q(\core.keymem.key_mem[6][32] ),
    .QN(_20306_));
 DFFR_X1 \core.keymem.key_mem[6][33]$_DFFE_PN0P_  (.D(_02299_),
    .RN(net99),
    .CK(clknet_leaf_112_clk),
    .Q(\core.keymem.key_mem[6][33] ),
    .QN(_20305_));
 DFFR_X1 \core.keymem.key_mem[6][34]$_DFFE_PN0P_  (.D(_02300_),
    .RN(net16),
    .CK(clknet_leaf_136_clk),
    .Q(\core.keymem.key_mem[6][34] ),
    .QN(_20304_));
 DFFR_X1 \core.keymem.key_mem[6][35]$_DFFE_PN0P_  (.D(_02301_),
    .RN(net99),
    .CK(clknet_leaf_122_clk),
    .Q(\core.keymem.key_mem[6][35] ),
    .QN(_20303_));
 DFFR_X1 \core.keymem.key_mem[6][36]$_DFFE_PN0P_  (.D(_02302_),
    .RN(net87),
    .CK(clknet_leaf_28_clk),
    .Q(\core.keymem.key_mem[6][36] ),
    .QN(_20302_));
 DFFR_X1 \core.keymem.key_mem[6][37]$_DFFE_PN0P_  (.D(_02303_),
    .RN(net89),
    .CK(clknet_leaf_84_clk),
    .Q(\core.keymem.key_mem[6][37] ),
    .QN(_20301_));
 DFFR_X1 \core.keymem.key_mem[6][38]$_DFFE_PN0P_  (.D(_02304_),
    .RN(net16),
    .CK(clknet_leaf_124_clk),
    .Q(\core.keymem.key_mem[6][38] ),
    .QN(_20300_));
 DFFR_X1 \core.keymem.key_mem[6][39]$_DFFE_PN0P_  (.D(_02305_),
    .RN(net89),
    .CK(clknet_leaf_86_clk),
    .Q(\core.keymem.key_mem[6][39] ),
    .QN(_20299_));
 DFFR_X1 \core.keymem.key_mem[6][3]$_DFFE_PN0P_  (.D(_02306_),
    .RN(net85),
    .CK(clknet_leaf_47_clk),
    .Q(\core.keymem.key_mem[6][3] ),
    .QN(_20298_));
 DFFR_X1 \core.keymem.key_mem[6][40]$_DFFE_PN0P_  (.D(_02307_),
    .RN(net88),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[6][40] ),
    .QN(_20297_));
 DFFR_X1 \core.keymem.key_mem[6][41]$_DFFE_PN0P_  (.D(_02308_),
    .RN(net99),
    .CK(clknet_leaf_82_clk),
    .Q(\core.keymem.key_mem[6][41] ),
    .QN(_20296_));
 DFFR_X1 \core.keymem.key_mem[6][42]$_DFFE_PN0P_  (.D(_02309_),
    .RN(net100),
    .CK(clknet_leaf_109_clk),
    .Q(\core.keymem.key_mem[6][42] ),
    .QN(_20295_));
 DFFR_X1 \core.keymem.key_mem[6][43]$_DFFE_PN0P_  (.D(_02310_),
    .RN(net85),
    .CK(clknet_leaf_88_clk),
    .Q(\core.keymem.key_mem[6][43] ),
    .QN(_20294_));
 DFFR_X1 \core.keymem.key_mem[6][44]$_DFFE_PN0P_  (.D(_02311_),
    .RN(net100),
    .CK(clknet_leaf_108_clk),
    .Q(\core.keymem.key_mem[6][44] ),
    .QN(_20293_));
 DFFR_X1 \core.keymem.key_mem[6][45]$_DFFE_PN0P_  (.D(_02312_),
    .RN(net89),
    .CK(clknet_leaf_68_clk),
    .Q(\core.keymem.key_mem[6][45] ),
    .QN(_20292_));
 DFFR_X1 \core.keymem.key_mem[6][46]$_DFFE_PN0P_  (.D(_02313_),
    .RN(net99),
    .CK(clknet_leaf_82_clk),
    .Q(\core.keymem.key_mem[6][46] ),
    .QN(_20291_));
 DFFR_X1 \core.keymem.key_mem[6][47]$_DFFE_PN0P_  (.D(_02314_),
    .RN(net98),
    .CK(clknet_leaf_175_clk),
    .Q(\core.keymem.key_mem[6][47] ),
    .QN(_20290_));
 DFFR_X1 \core.keymem.key_mem[6][48]$_DFFE_PN0P_  (.D(_02315_),
    .RN(net99),
    .CK(clknet_leaf_119_clk),
    .Q(\core.keymem.key_mem[6][48] ),
    .QN(_20289_));
 DFFR_X1 \core.keymem.key_mem[6][49]$_DFFE_PN0P_  (.D(_02316_),
    .RN(net99),
    .CK(clknet_leaf_81_clk),
    .Q(\core.keymem.key_mem[6][49] ),
    .QN(_20288_));
 DFFR_X1 \core.keymem.key_mem[6][4]$_DFFE_PN0P_  (.D(_02317_),
    .RN(net100),
    .CK(clknet_leaf_106_clk),
    .Q(\core.keymem.key_mem[6][4] ),
    .QN(_20287_));
 DFFR_X1 \core.keymem.key_mem[6][50]$_DFFE_PN0P_  (.D(_02318_),
    .RN(net98),
    .CK(clknet_leaf_137_clk),
    .Q(\core.keymem.key_mem[6][50] ),
    .QN(_20286_));
 DFFR_X1 \core.keymem.key_mem[6][51]$_DFFE_PN0P_  (.D(_02319_),
    .RN(net100),
    .CK(clknet_leaf_130_clk),
    .Q(\core.keymem.key_mem[6][51] ),
    .QN(_20285_));
 DFFR_X1 \core.keymem.key_mem[6][52]$_DFFE_PN0P_  (.D(_02320_),
    .RN(net99),
    .CK(clknet_leaf_78_clk),
    .Q(\core.keymem.key_mem[6][52] ),
    .QN(_20284_));
 DFFR_X1 \core.keymem.key_mem[6][53]$_DFFE_PN0P_  (.D(_02321_),
    .RN(net98),
    .CK(clknet_leaf_176_clk),
    .Q(\core.keymem.key_mem[6][53] ),
    .QN(_20283_));
 DFFR_X1 \core.keymem.key_mem[6][54]$_DFFE_PN0P_  (.D(_02322_),
    .RN(net98),
    .CK(clknet_leaf_142_clk),
    .Q(\core.keymem.key_mem[6][54] ),
    .QN(_20282_));
 DFFR_X1 \core.keymem.key_mem[6][55]$_DFFE_PN0P_  (.D(_02323_),
    .RN(net16),
    .CK(clknet_leaf_135_clk),
    .Q(\core.keymem.key_mem[6][55] ),
    .QN(_20281_));
 DFFR_X1 \core.keymem.key_mem[6][56]$_DFFE_PN0P_  (.D(_02324_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[6][56] ),
    .QN(_20280_));
 DFFR_X1 \core.keymem.key_mem[6][57]$_DFFE_PN0P_  (.D(_02325_),
    .RN(net100),
    .CK(clknet_leaf_108_clk),
    .Q(\core.keymem.key_mem[6][57] ),
    .QN(_20279_));
 DFFR_X1 \core.keymem.key_mem[6][58]$_DFFE_PN0P_  (.D(_02326_),
    .RN(net100),
    .CK(clknet_leaf_102_clk),
    .Q(\core.keymem.key_mem[6][58] ),
    .QN(_20278_));
 DFFR_X1 \core.keymem.key_mem[6][59]$_DFFE_PN0P_  (.D(_02327_),
    .RN(net100),
    .CK(clknet_leaf_20_clk),
    .Q(\core.keymem.key_mem[6][59] ),
    .QN(_20277_));
 DFFR_X1 \core.keymem.key_mem[6][5]$_DFFE_PN0P_  (.D(_02328_),
    .RN(net100),
    .CK(clknet_leaf_18_clk),
    .Q(\core.keymem.key_mem[6][5] ),
    .QN(_20276_));
 DFFR_X1 \core.keymem.key_mem[6][60]$_DFFE_PN0P_  (.D(_02329_),
    .RN(net89),
    .CK(clknet_leaf_24_clk),
    .Q(\core.keymem.key_mem[6][60] ),
    .QN(_20275_));
 DFFR_X1 \core.keymem.key_mem[6][61]$_DFFE_PN0P_  (.D(_02330_),
    .RN(net88),
    .CK(clknet_leaf_93_clk),
    .Q(\core.keymem.key_mem[6][61] ),
    .QN(_20274_));
 DFFR_X1 \core.keymem.key_mem[6][62]$_DFFE_PN0P_  (.D(_02331_),
    .RN(net100),
    .CK(clknet_leaf_99_clk),
    .Q(\core.keymem.key_mem[6][62] ),
    .QN(_20273_));
 DFFR_X1 \core.keymem.key_mem[6][63]$_DFFE_PN0P_  (.D(_02332_),
    .RN(net100),
    .CK(clknet_leaf_20_clk),
    .Q(\core.keymem.key_mem[6][63] ),
    .QN(_20272_));
 DFFR_X1 \core.keymem.key_mem[6][64]$_DFFE_PN0P_  (.D(_02333_),
    .RN(net82),
    .CK(clknet_leaf_14_clk),
    .Q(\core.keymem.key_mem[6][64] ),
    .QN(_20271_));
 DFFR_X1 \core.keymem.key_mem[6][65]$_DFFE_PN0P_  (.D(_02334_),
    .RN(net99),
    .CK(clknet_leaf_120_clk),
    .Q(\core.keymem.key_mem[6][65] ),
    .QN(_20270_));
 DFFR_X1 \core.keymem.key_mem[6][66]$_DFFE_PN0P_  (.D(_02335_),
    .RN(net100),
    .CK(clknet_leaf_16_clk),
    .Q(\core.keymem.key_mem[6][66] ),
    .QN(_20269_));
 DFFR_X1 \core.keymem.key_mem[6][67]$_DFFE_PN0P_  (.D(_02336_),
    .RN(net95),
    .CK(clknet_leaf_77_clk),
    .Q(\core.keymem.key_mem[6][67] ),
    .QN(_20268_));
 DFFR_X1 \core.keymem.key_mem[6][68]$_DFFE_PN0P_  (.D(_02337_),
    .RN(net99),
    .CK(clknet_leaf_118_clk),
    .Q(\core.keymem.key_mem[6][68] ),
    .QN(_20267_));
 DFFR_X1 \core.keymem.key_mem[6][69]$_DFFE_PN0P_  (.D(_02338_),
    .RN(net95),
    .CK(clknet_leaf_180_clk),
    .Q(\core.keymem.key_mem[6][69] ),
    .QN(_20266_));
 DFFR_X1 \core.keymem.key_mem[6][6]$_DFFE_PN0P_  (.D(_02339_),
    .RN(net89),
    .CK(clknet_leaf_94_clk),
    .Q(\core.keymem.key_mem[6][6] ),
    .QN(_20265_));
 DFFR_X1 \core.keymem.key_mem[6][70]$_DFFE_PN0P_  (.D(_02340_),
    .RN(net100),
    .CK(clknet_leaf_101_clk),
    .Q(\core.keymem.key_mem[6][70] ),
    .QN(_20264_));
 DFFR_X1 \core.keymem.key_mem[6][71]$_DFFE_PN0P_  (.D(_02341_),
    .RN(net99),
    .CK(clknet_leaf_75_clk),
    .Q(\core.keymem.key_mem[6][71] ),
    .QN(_20263_));
 DFFR_X1 \core.keymem.key_mem[6][72]$_DFFE_PN0P_  (.D(_02342_),
    .RN(net95),
    .CK(clknet_leaf_75_clk),
    .Q(\core.keymem.key_mem[6][72] ),
    .QN(_20262_));
 DFFR_X1 \core.keymem.key_mem[6][73]$_DFFE_PN0P_  (.D(_02343_),
    .RN(net97),
    .CK(clknet_leaf_147_clk),
    .Q(\core.keymem.key_mem[6][73] ),
    .QN(_20261_));
 DFFR_X1 \core.keymem.key_mem[6][74]$_DFFE_PN0P_  (.D(_02344_),
    .RN(net97),
    .CK(clknet_leaf_156_clk),
    .Q(\core.keymem.key_mem[6][74] ),
    .QN(_20260_));
 DFFR_X1 \core.keymem.key_mem[6][75]$_DFFE_PN0P_  (.D(_02345_),
    .RN(net97),
    .CK(clknet_leaf_153_clk),
    .Q(\core.keymem.key_mem[6][75] ),
    .QN(_20259_));
 DFFR_X1 \core.keymem.key_mem[6][76]$_DFFE_PN0P_  (.D(_02346_),
    .RN(net93),
    .CK(clknet_leaf_282_clk),
    .Q(\core.keymem.key_mem[6][76] ),
    .QN(_20258_));
 DFFR_X1 \core.keymem.key_mem[6][77]$_DFFE_PN0P_  (.D(_02347_),
    .RN(net97),
    .CK(clknet_leaf_159_clk),
    .Q(\core.keymem.key_mem[6][77] ),
    .QN(_20257_));
 DFFR_X1 \core.keymem.key_mem[6][78]$_DFFE_PN0P_  (.D(_02348_),
    .RN(net96),
    .CK(clknet_leaf_171_clk),
    .Q(\core.keymem.key_mem[6][78] ),
    .QN(_20256_));
 DFFR_X1 \core.keymem.key_mem[6][79]$_DFFE_PN0P_  (.D(_02349_),
    .RN(net96),
    .CK(clknet_leaf_227_clk),
    .Q(\core.keymem.key_mem[6][79] ),
    .QN(_20255_));
 DFFR_X1 \core.keymem.key_mem[6][7]$_DFFE_PN0P_  (.D(_02350_),
    .RN(net98),
    .CK(clknet_leaf_174_clk),
    .Q(\core.keymem.key_mem[6][7] ),
    .QN(_20254_));
 DFFR_X1 \core.keymem.key_mem[6][80]$_DFFE_PN0P_  (.D(_02351_),
    .RN(net97),
    .CK(clknet_leaf_158_clk),
    .Q(\core.keymem.key_mem[6][80] ),
    .QN(_20253_));
 DFFR_X1 \core.keymem.key_mem[6][81]$_DFFE_PN0P_  (.D(_02352_),
    .RN(net97),
    .CK(clknet_leaf_153_clk),
    .Q(\core.keymem.key_mem[6][81] ),
    .QN(_20252_));
 DFFR_X1 \core.keymem.key_mem[6][82]$_DFFE_PN0P_  (.D(_02353_),
    .RN(net98),
    .CK(clknet_leaf_169_clk),
    .Q(\core.keymem.key_mem[6][82] ),
    .QN(_20251_));
 DFFR_X1 \core.keymem.key_mem[6][83]$_DFFE_PN0P_  (.D(_02354_),
    .RN(net93),
    .CK(clknet_leaf_182_clk),
    .Q(\core.keymem.key_mem[6][83] ),
    .QN(_20250_));
 DFFR_X1 \core.keymem.key_mem[6][84]$_DFFE_PN0P_  (.D(_02355_),
    .RN(net95),
    .CK(clknet_leaf_182_clk),
    .Q(\core.keymem.key_mem[6][84] ),
    .QN(_20249_));
 DFFR_X1 \core.keymem.key_mem[6][85]$_DFFE_PN0P_  (.D(_02356_),
    .RN(net97),
    .CK(clknet_leaf_239_clk),
    .Q(\core.keymem.key_mem[6][85] ),
    .QN(_20248_));
 DFFR_X1 \core.keymem.key_mem[6][86]$_DFFE_PN0P_  (.D(_02357_),
    .RN(net97),
    .CK(clknet_leaf_159_clk),
    .Q(\core.keymem.key_mem[6][86] ),
    .QN(_20247_));
 DFFR_X1 \core.keymem.key_mem[6][87]$_DFFE_PN0P_  (.D(_02358_),
    .RN(net89),
    .CK(clknet_leaf_56_clk),
    .Q(\core.keymem.key_mem[6][87] ),
    .QN(_20246_));
 DFFR_X1 \core.keymem.key_mem[6][88]$_DFFE_PN0P_  (.D(_02359_),
    .RN(net93),
    .CK(clknet_leaf_282_clk),
    .Q(\core.keymem.key_mem[6][88] ),
    .QN(_20245_));
 DFFR_X1 \core.keymem.key_mem[6][89]$_DFFE_PN0P_  (.D(_02360_),
    .RN(net93),
    .CK(clknet_leaf_199_clk),
    .Q(\core.keymem.key_mem[6][89] ),
    .QN(_20244_));
 DFFR_X1 \core.keymem.key_mem[6][8]$_DFFE_PN0P_  (.D(_02361_),
    .RN(net93),
    .CK(clknet_leaf_281_clk),
    .Q(\core.keymem.key_mem[6][8] ),
    .QN(_20243_));
 DFFR_X1 \core.keymem.key_mem[6][90]$_DFFE_PN0P_  (.D(_02362_),
    .RN(net97),
    .CK(clknet_leaf_161_clk),
    .Q(\core.keymem.key_mem[6][90] ),
    .QN(_20242_));
 DFFR_X1 \core.keymem.key_mem[6][91]$_DFFE_PN0P_  (.D(_02363_),
    .RN(net93),
    .CK(clknet_leaf_184_clk),
    .Q(\core.keymem.key_mem[6][91] ),
    .QN(_20241_));
 DFFR_X1 \core.keymem.key_mem[6][92]$_DFFE_PN0P_  (.D(_02364_),
    .RN(net95),
    .CK(clknet_leaf_72_clk),
    .Q(\core.keymem.key_mem[6][92] ),
    .QN(_20240_));
 DFFR_X1 \core.keymem.key_mem[6][93]$_DFFE_PN0P_  (.D(_02365_),
    .RN(net97),
    .CK(clknet_leaf_162_clk),
    .Q(\core.keymem.key_mem[6][93] ),
    .QN(_20239_));
 DFFR_X1 \core.keymem.key_mem[6][94]$_DFFE_PN0P_  (.D(_02366_),
    .RN(net94),
    .CK(clknet_leaf_213_clk),
    .Q(\core.keymem.key_mem[6][94] ),
    .QN(_20238_));
 DFFR_X1 \core.keymem.key_mem[6][95]$_DFFE_PN0P_  (.D(_02367_),
    .RN(net96),
    .CK(clknet_leaf_244_clk),
    .Q(\core.keymem.key_mem[6][95] ),
    .QN(_20237_));
 DFFR_X1 \core.keymem.key_mem[6][96]$_DFFE_PN0P_  (.D(_02368_),
    .RN(net92),
    .CK(clknet_leaf_276_clk),
    .Q(\core.keymem.key_mem[6][96] ),
    .QN(_20236_));
 DFFR_X1 \core.keymem.key_mem[6][97]$_DFFE_PN0P_  (.D(_02369_),
    .RN(net95),
    .CK(clknet_leaf_194_clk),
    .Q(\core.keymem.key_mem[6][97] ),
    .QN(_20235_));
 DFFR_X1 \core.keymem.key_mem[6][98]$_DFFE_PN0P_  (.D(_02370_),
    .RN(net93),
    .CK(clknet_leaf_193_clk),
    .Q(\core.keymem.key_mem[6][98] ),
    .QN(_20234_));
 DFFR_X1 \core.keymem.key_mem[6][99]$_DFFE_PN0P_  (.D(_02371_),
    .RN(net92),
    .CK(clknet_leaf_202_clk),
    .Q(\core.keymem.key_mem[6][99] ),
    .QN(_20233_));
 DFFR_X1 \core.keymem.key_mem[6][9]$_DFFE_PN0P_  (.D(_02372_),
    .RN(net92),
    .CK(clknet_leaf_203_clk),
    .Q(\core.keymem.key_mem[6][9] ),
    .QN(_20232_));
 DFFR_X1 \core.keymem.key_mem[7][0]$_DFFE_PN0P_  (.D(_02373_),
    .RN(net96),
    .CK(clknet_leaf_248_clk),
    .Q(\core.keymem.key_mem[7][0] ),
    .QN(_20231_));
 DFFR_X1 \core.keymem.key_mem[7][100]$_DFFE_PN0P_  (.D(_02374_),
    .RN(net98),
    .CK(clknet_leaf_211_clk),
    .Q(\core.keymem.key_mem[7][100] ),
    .QN(_20230_));
 DFFR_X1 \core.keymem.key_mem[7][101]$_DFFE_PN0P_  (.D(_02375_),
    .RN(net94),
    .CK(clknet_leaf_218_clk),
    .Q(\core.keymem.key_mem[7][101] ),
    .QN(_20229_));
 DFFR_X1 \core.keymem.key_mem[7][102]$_DFFE_PN0P_  (.D(_02376_),
    .RN(net96),
    .CK(clknet_leaf_232_clk),
    .Q(\core.keymem.key_mem[7][102] ),
    .QN(_20228_));
 DFFR_X1 \core.keymem.key_mem[7][103]$_DFFE_PN0P_  (.D(_02377_),
    .RN(net96),
    .CK(clknet_leaf_224_clk),
    .Q(\core.keymem.key_mem[7][103] ),
    .QN(_20227_));
 DFFR_X1 \core.keymem.key_mem[7][104]$_DFFE_PN0P_  (.D(_02378_),
    .RN(net93),
    .CK(clknet_leaf_193_clk),
    .Q(\core.keymem.key_mem[7][104] ),
    .QN(_20226_));
 DFFR_X1 \core.keymem.key_mem[7][105]$_DFFE_PN0P_  (.D(_02379_),
    .RN(net96),
    .CK(clknet_leaf_246_clk),
    .Q(\core.keymem.key_mem[7][105] ),
    .QN(_20225_));
 DFFR_X1 \core.keymem.key_mem[7][106]$_DFFE_PN0P_  (.D(_02380_),
    .RN(net92),
    .CK(clknet_leaf_268_clk),
    .Q(\core.keymem.key_mem[7][106] ),
    .QN(_20224_));
 DFFR_X1 \core.keymem.key_mem[7][107]$_DFFE_PN0P_  (.D(_02381_),
    .RN(net92),
    .CK(clknet_leaf_267_clk),
    .Q(\core.keymem.key_mem[7][107] ),
    .QN(_20223_));
 DFFR_X1 \core.keymem.key_mem[7][108]$_DFFE_PN0P_  (.D(_02382_),
    .RN(net91),
    .CK(clknet_leaf_277_clk),
    .Q(\core.keymem.key_mem[7][108] ),
    .QN(_20222_));
 DFFR_X1 \core.keymem.key_mem[7][109]$_DFFE_PN0P_  (.D(_02383_),
    .RN(net94),
    .CK(clknet_leaf_258_clk),
    .Q(\core.keymem.key_mem[7][109] ),
    .QN(_20221_));
 DFFR_X1 \core.keymem.key_mem[7][10]$_DFFE_PN0P_  (.D(_02384_),
    .RN(net98),
    .CK(clknet_leaf_167_clk),
    .Q(\core.keymem.key_mem[7][10] ),
    .QN(_20220_));
 DFFR_X1 \core.keymem.key_mem[7][110]$_DFFE_PN0P_  (.D(_02385_),
    .RN(net96),
    .CK(clknet_leaf_249_clk),
    .Q(\core.keymem.key_mem[7][110] ),
    .QN(_20219_));
 DFFR_X1 \core.keymem.key_mem[7][111]$_DFFE_PN0P_  (.D(_02386_),
    .RN(net96),
    .CK(clknet_leaf_225_clk),
    .Q(\core.keymem.key_mem[7][111] ),
    .QN(_20218_));
 DFFR_X1 \core.keymem.key_mem[7][112]$_DFFE_PN0P_  (.D(_02387_),
    .RN(net94),
    .CK(clknet_leaf_260_clk),
    .Q(\core.keymem.key_mem[7][112] ),
    .QN(_20217_));
 DFFR_X1 \core.keymem.key_mem[7][113]$_DFFE_PN0P_  (.D(_02388_),
    .RN(net91),
    .CK(clknet_leaf_273_clk),
    .Q(\core.keymem.key_mem[7][113] ),
    .QN(_20216_));
 DFFR_X1 \core.keymem.key_mem[7][114]$_DFFE_PN0P_  (.D(_02389_),
    .RN(net91),
    .CK(clknet_leaf_279_clk),
    .Q(\core.keymem.key_mem[7][114] ),
    .QN(_20215_));
 DFFR_X1 \core.keymem.key_mem[7][115]$_DFFE_PN0P_  (.D(_02390_),
    .RN(net92),
    .CK(clknet_leaf_272_clk),
    .Q(\core.keymem.key_mem[7][115] ),
    .QN(_20214_));
 DFFR_X1 \core.keymem.key_mem[7][116]$_DFFE_PN0P_  (.D(_02391_),
    .RN(net94),
    .CK(clknet_leaf_215_clk),
    .Q(\core.keymem.key_mem[7][116] ),
    .QN(_20213_));
 DFFR_X1 \core.keymem.key_mem[7][117]$_DFFE_PN0P_  (.D(_02392_),
    .RN(net96),
    .CK(clknet_leaf_225_clk),
    .Q(\core.keymem.key_mem[7][117] ),
    .QN(_20212_));
 DFFR_X1 \core.keymem.key_mem[7][118]$_DFFE_PN0P_  (.D(_02393_),
    .RN(net96),
    .CK(clknet_leaf_243_clk),
    .Q(\core.keymem.key_mem[7][118] ),
    .QN(_20211_));
 DFFR_X1 \core.keymem.key_mem[7][119]$_DFFE_PN0P_  (.D(_02394_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[7][119] ),
    .QN(_20210_));
 DFFR_X1 \core.keymem.key_mem[7][11]$_DFFE_PN0P_  (.D(_02395_),
    .RN(net95),
    .CK(clknet_leaf_61_clk),
    .Q(\core.keymem.key_mem[7][11] ),
    .QN(_20209_));
 DFFR_X1 \core.keymem.key_mem[7][120]$_DFFE_PN0P_  (.D(_02396_),
    .RN(net94),
    .CK(clknet_leaf_215_clk),
    .Q(\core.keymem.key_mem[7][120] ),
    .QN(_20208_));
 DFFR_X1 \core.keymem.key_mem[7][121]$_DFFE_PN0P_  (.D(_02397_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[7][121] ),
    .QN(_20207_));
 DFFR_X1 \core.keymem.key_mem[7][122]$_DFFE_PN0P_  (.D(_02398_),
    .RN(net97),
    .CK(clknet_leaf_237_clk),
    .Q(\core.keymem.key_mem[7][122] ),
    .QN(_20206_));
 DFFR_X1 \core.keymem.key_mem[7][123]$_DFFE_PN0P_  (.D(_02399_),
    .RN(net93),
    .CK(clknet_leaf_198_clk),
    .Q(\core.keymem.key_mem[7][123] ),
    .QN(_20205_));
 DFFR_X1 \core.keymem.key_mem[7][124]$_DFFE_PN0P_  (.D(_02400_),
    .RN(net93),
    .CK(clknet_leaf_198_clk),
    .Q(\core.keymem.key_mem[7][124] ),
    .QN(_20204_));
 DFFR_X1 \core.keymem.key_mem[7][125]$_DFFE_PN0P_  (.D(_02401_),
    .RN(net97),
    .CK(clknet_leaf_231_clk),
    .Q(\core.keymem.key_mem[7][125] ),
    .QN(_20203_));
 DFFR_X1 \core.keymem.key_mem[7][126]$_DFFE_PN0P_  (.D(_02402_),
    .RN(net98),
    .CK(clknet_leaf_167_clk),
    .Q(\core.keymem.key_mem[7][126] ),
    .QN(_20202_));
 DFFR_X1 \core.keymem.key_mem[7][127]$_DFFE_PN0P_  (.D(_02403_),
    .RN(net97),
    .CK(clknet_leaf_243_clk),
    .Q(\core.keymem.key_mem[7][127] ),
    .QN(_20201_));
 DFFR_X1 \core.keymem.key_mem[7][12]$_DFFE_PN0P_  (.D(_02404_),
    .RN(net93),
    .CK(clknet_leaf_191_clk),
    .Q(\core.keymem.key_mem[7][12] ),
    .QN(_20200_));
 DFFR_X1 \core.keymem.key_mem[7][13]$_DFFE_PN0P_  (.D(_02405_),
    .RN(net87),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[7][13] ),
    .QN(_20199_));
 DFFR_X1 \core.keymem.key_mem[7][14]$_DFFE_PN0P_  (.D(_02406_),
    .RN(net94),
    .CK(clknet_leaf_211_clk),
    .Q(\core.keymem.key_mem[7][14] ),
    .QN(_20198_));
 DFFR_X1 \core.keymem.key_mem[7][15]$_DFFE_PN0P_  (.D(_02407_),
    .RN(net96),
    .CK(clknet_leaf_171_clk),
    .Q(\core.keymem.key_mem[7][15] ),
    .QN(_20197_));
 DFFR_X1 \core.keymem.key_mem[7][16]$_DFFE_PN0P_  (.D(_02408_),
    .RN(net87),
    .CK(clknet_leaf_33_clk),
    .Q(\core.keymem.key_mem[7][16] ),
    .QN(_20196_));
 DFFR_X1 \core.keymem.key_mem[7][17]$_DFFE_PN0P_  (.D(_02409_),
    .RN(net98),
    .CK(clknet_leaf_171_clk),
    .Q(\core.keymem.key_mem[7][17] ),
    .QN(_20195_));
 DFFR_X1 \core.keymem.key_mem[7][18]$_DFFE_PN0P_  (.D(_02410_),
    .RN(net89),
    .CK(clknet_leaf_26_clk),
    .Q(\core.keymem.key_mem[7][18] ),
    .QN(_20194_));
 DFFR_X1 \core.keymem.key_mem[7][19]$_DFFE_PN0P_  (.D(_02411_),
    .RN(net85),
    .CK(clknet_leaf_50_clk),
    .Q(\core.keymem.key_mem[7][19] ),
    .QN(_20193_));
 DFFR_X1 \core.keymem.key_mem[7][1]$_DFFE_PN0P_  (.D(_02412_),
    .RN(net89),
    .CK(clknet_leaf_26_clk),
    .Q(\core.keymem.key_mem[7][1] ),
    .QN(_20192_));
 DFFR_X1 \core.keymem.key_mem[7][20]$_DFFE_PN0P_  (.D(_02413_),
    .RN(net89),
    .CK(clknet_leaf_95_clk),
    .Q(\core.keymem.key_mem[7][20] ),
    .QN(_20191_));
 DFFR_X1 \core.keymem.key_mem[7][21]$_DFFE_PN0P_  (.D(_02414_),
    .RN(net89),
    .CK(clknet_leaf_69_clk),
    .Q(\core.keymem.key_mem[7][21] ),
    .QN(_20190_));
 DFFR_X1 \core.keymem.key_mem[7][22]$_DFFE_PN0P_  (.D(_02415_),
    .RN(net96),
    .CK(clknet_leaf_249_clk),
    .Q(\core.keymem.key_mem[7][22] ),
    .QN(_20189_));
 DFFR_X1 \core.keymem.key_mem[7][23]$_DFFE_PN0P_  (.D(_02416_),
    .RN(net89),
    .CK(clknet_leaf_55_clk),
    .Q(\core.keymem.key_mem[7][23] ),
    .QN(_20188_));
 DFFR_X1 \core.keymem.key_mem[7][24]$_DFFE_PN0P_  (.D(_02417_),
    .RN(net85),
    .CK(clknet_leaf_50_clk),
    .Q(\core.keymem.key_mem[7][24] ),
    .QN(_20187_));
 DFFR_X1 \core.keymem.key_mem[7][25]$_DFFE_PN0P_  (.D(_02418_),
    .RN(net85),
    .CK(clknet_leaf_48_clk),
    .Q(\core.keymem.key_mem[7][25] ),
    .QN(_20186_));
 DFFR_X1 \core.keymem.key_mem[7][26]$_DFFE_PN0P_  (.D(_02419_),
    .RN(net89),
    .CK(clknet_leaf_27_clk),
    .Q(\core.keymem.key_mem[7][26] ),
    .QN(_20185_));
 DFFR_X1 \core.keymem.key_mem[7][27]$_DFFE_PN0P_  (.D(_02420_),
    .RN(net16),
    .CK(clknet_leaf_151_clk),
    .Q(\core.keymem.key_mem[7][27] ),
    .QN(_20184_));
 DFFR_X1 \core.keymem.key_mem[7][28]$_DFFE_PN0P_  (.D(_02421_),
    .RN(net16),
    .CK(clknet_leaf_125_clk),
    .Q(\core.keymem.key_mem[7][28] ),
    .QN(_20183_));
 DFFR_X1 \core.keymem.key_mem[7][29]$_DFFE_PN0P_  (.D(_02422_),
    .RN(net16),
    .CK(clknet_leaf_149_clk),
    .Q(\core.keymem.key_mem[7][29] ),
    .QN(_20182_));
 DFFR_X1 \core.keymem.key_mem[7][2]$_DFFE_PN0P_  (.D(_02423_),
    .RN(net89),
    .CK(clknet_leaf_64_clk),
    .Q(\core.keymem.key_mem[7][2] ),
    .QN(_20181_));
 DFFR_X1 \core.keymem.key_mem[7][30]$_DFFE_PN0P_  (.D(_02424_),
    .RN(net98),
    .CK(clknet_leaf_144_clk),
    .Q(\core.keymem.key_mem[7][30] ),
    .QN(_20180_));
 DFFR_X1 \core.keymem.key_mem[7][31]$_DFFE_PN0P_  (.D(_02425_),
    .RN(net98),
    .CK(clknet_leaf_139_clk),
    .Q(\core.keymem.key_mem[7][31] ),
    .QN(_20179_));
 DFFR_X1 \core.keymem.key_mem[7][32]$_DFFE_PN0P_  (.D(_02426_),
    .RN(net99),
    .CK(clknet_leaf_116_clk),
    .Q(\core.keymem.key_mem[7][32] ),
    .QN(_20178_));
 DFFR_X1 \core.keymem.key_mem[7][33]$_DFFE_PN0P_  (.D(_02427_),
    .RN(net99),
    .CK(clknet_leaf_127_clk),
    .Q(\core.keymem.key_mem[7][33] ),
    .QN(_20177_));
 DFFR_X1 \core.keymem.key_mem[7][34]$_DFFE_PN0P_  (.D(_02428_),
    .RN(net16),
    .CK(clknet_leaf_136_clk),
    .Q(\core.keymem.key_mem[7][34] ),
    .QN(_20176_));
 DFFR_X1 \core.keymem.key_mem[7][35]$_DFFE_PN0P_  (.D(_02429_),
    .RN(net99),
    .CK(clknet_leaf_128_clk),
    .Q(\core.keymem.key_mem[7][35] ),
    .QN(_20175_));
 DFFR_X1 \core.keymem.key_mem[7][36]$_DFFE_PN0P_  (.D(_02430_),
    .RN(net88),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[7][36] ),
    .QN(_20174_));
 DFFR_X1 \core.keymem.key_mem[7][37]$_DFFE_PN0P_  (.D(_02431_),
    .RN(net89),
    .CK(clknet_leaf_85_clk),
    .Q(\core.keymem.key_mem[7][37] ),
    .QN(_20173_));
 DFFR_X1 \core.keymem.key_mem[7][38]$_DFFE_PN0P_  (.D(_02432_),
    .RN(net99),
    .CK(clknet_leaf_123_clk),
    .Q(\core.keymem.key_mem[7][38] ),
    .QN(_20172_));
 DFFR_X1 \core.keymem.key_mem[7][39]$_DFFE_PN0P_  (.D(_02433_),
    .RN(net99),
    .CK(clknet_leaf_86_clk),
    .Q(\core.keymem.key_mem[7][39] ),
    .QN(_20171_));
 DFFR_X1 \core.keymem.key_mem[7][3]$_DFFE_PN0P_  (.D(_02434_),
    .RN(net85),
    .CK(clknet_leaf_47_clk),
    .Q(\core.keymem.key_mem[7][3] ),
    .QN(_20170_));
 DFFR_X1 \core.keymem.key_mem[7][40]$_DFFE_PN0P_  (.D(_02435_),
    .RN(net85),
    .CK(clknet_leaf_30_clk),
    .Q(\core.keymem.key_mem[7][40] ),
    .QN(_20169_));
 DFFR_X1 \core.keymem.key_mem[7][41]$_DFFE_PN0P_  (.D(_02436_),
    .RN(net89),
    .CK(clknet_leaf_82_clk),
    .Q(\core.keymem.key_mem[7][41] ),
    .QN(_20168_));
 DFFR_X1 \core.keymem.key_mem[7][42]$_DFFE_PN0P_  (.D(_02437_),
    .RN(net100),
    .CK(clknet_leaf_109_clk),
    .Q(\core.keymem.key_mem[7][42] ),
    .QN(_20167_));
 DFFR_X1 \core.keymem.key_mem[7][43]$_DFFE_PN0P_  (.D(_02438_),
    .RN(net85),
    .CK(clknet_leaf_88_clk),
    .Q(\core.keymem.key_mem[7][43] ),
    .QN(_20166_));
 DFFR_X1 \core.keymem.key_mem[7][44]$_DFFE_PN0P_  (.D(_02439_),
    .RN(net100),
    .CK(clknet_leaf_105_clk),
    .Q(\core.keymem.key_mem[7][44] ),
    .QN(_20165_));
 DFFR_X1 \core.keymem.key_mem[7][45]$_DFFE_PN0P_  (.D(_02440_),
    .RN(net99),
    .CK(clknet_leaf_71_clk),
    .Q(\core.keymem.key_mem[7][45] ),
    .QN(_20164_));
 DFFR_X1 \core.keymem.key_mem[7][46]$_DFFE_PN0P_  (.D(_02441_),
    .RN(net99),
    .CK(clknet_leaf_86_clk),
    .Q(\core.keymem.key_mem[7][46] ),
    .QN(_20163_));
 DFFR_X1 \core.keymem.key_mem[7][47]$_DFFE_PN0P_  (.D(_02442_),
    .RN(net98),
    .CK(clknet_leaf_180_clk),
    .Q(\core.keymem.key_mem[7][47] ),
    .QN(_20162_));
 DFFR_X1 \core.keymem.key_mem[7][48]$_DFFE_PN0P_  (.D(_02443_),
    .RN(net95),
    .CK(clknet_leaf_119_clk),
    .Q(\core.keymem.key_mem[7][48] ),
    .QN(_20161_));
 DFFR_X1 \core.keymem.key_mem[7][49]$_DFFE_PN0P_  (.D(_02444_),
    .RN(net99),
    .CK(clknet_leaf_79_clk),
    .Q(\core.keymem.key_mem[7][49] ),
    .QN(_20160_));
 DFFR_X1 \core.keymem.key_mem[7][4]$_DFFE_PN0P_  (.D(_02445_),
    .RN(net100),
    .CK(clknet_leaf_105_clk),
    .Q(\core.keymem.key_mem[7][4] ),
    .QN(_20159_));
 DFFR_X1 \core.keymem.key_mem[7][50]$_DFFE_PN0P_  (.D(_02446_),
    .RN(net98),
    .CK(clknet_leaf_139_clk),
    .Q(\core.keymem.key_mem[7][50] ),
    .QN(_20158_));
 DFFR_X1 \core.keymem.key_mem[7][51]$_DFFE_PN0P_  (.D(_02447_),
    .RN(net100),
    .CK(clknet_leaf_129_clk),
    .Q(\core.keymem.key_mem[7][51] ),
    .QN(_20157_));
 DFFR_X1 \core.keymem.key_mem[7][52]$_DFFE_PN0P_  (.D(_02448_),
    .RN(net99),
    .CK(clknet_leaf_79_clk),
    .Q(\core.keymem.key_mem[7][52] ),
    .QN(_20156_));
 DFFR_X1 \core.keymem.key_mem[7][53]$_DFFE_PN0P_  (.D(_02449_),
    .RN(net98),
    .CK(clknet_leaf_176_clk),
    .Q(\core.keymem.key_mem[7][53] ),
    .QN(_20155_));
 DFFR_X1 \core.keymem.key_mem[7][54]$_DFFE_PN0P_  (.D(_02450_),
    .RN(net98),
    .CK(clknet_leaf_143_clk),
    .Q(\core.keymem.key_mem[7][54] ),
    .QN(_20154_));
 DFFR_X1 \core.keymem.key_mem[7][55]$_DFFE_PN0P_  (.D(_02451_),
    .RN(net16),
    .CK(clknet_leaf_135_clk),
    .Q(\core.keymem.key_mem[7][55] ),
    .QN(_20153_));
 DFFR_X1 \core.keymem.key_mem[7][56]$_DFFE_PN0P_  (.D(_02452_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[7][56] ),
    .QN(_20152_));
 DFFR_X1 \core.keymem.key_mem[7][57]$_DFFE_PN0P_  (.D(_02453_),
    .RN(net100),
    .CK(clknet_leaf_107_clk),
    .Q(\core.keymem.key_mem[7][57] ),
    .QN(_20151_));
 DFFR_X1 \core.keymem.key_mem[7][58]$_DFFE_PN0P_  (.D(_02454_),
    .RN(net100),
    .CK(clknet_leaf_107_clk),
    .Q(\core.keymem.key_mem[7][58] ),
    .QN(_20150_));
 DFFR_X1 \core.keymem.key_mem[7][59]$_DFFE_PN0P_  (.D(_02455_),
    .RN(net100),
    .CK(clknet_leaf_18_clk),
    .Q(\core.keymem.key_mem[7][59] ),
    .QN(_20149_));
 DFFR_X1 \core.keymem.key_mem[7][5]$_DFFE_PN0P_  (.D(_02456_),
    .RN(net100),
    .CK(clknet_leaf_20_clk),
    .Q(\core.keymem.key_mem[7][5] ),
    .QN(_20148_));
 DFFR_X1 \core.keymem.key_mem[7][60]$_DFFE_PN0P_  (.D(_02457_),
    .RN(net82),
    .CK(clknet_leaf_23_clk),
    .Q(\core.keymem.key_mem[7][60] ),
    .QN(_20147_));
 DFFR_X1 \core.keymem.key_mem[7][61]$_DFFE_PN0P_  (.D(_02458_),
    .RN(net89),
    .CK(clknet_leaf_94_clk),
    .Q(\core.keymem.key_mem[7][61] ),
    .QN(_20146_));
 DFFR_X1 \core.keymem.key_mem[7][62]$_DFFE_PN0P_  (.D(_02459_),
    .RN(net100),
    .CK(clknet_leaf_97_clk),
    .Q(\core.keymem.key_mem[7][62] ),
    .QN(_20145_));
 DFFR_X1 \core.keymem.key_mem[7][63]$_DFFE_PN0P_  (.D(_02460_),
    .RN(net100),
    .CK(clknet_leaf_95_clk),
    .Q(\core.keymem.key_mem[7][63] ),
    .QN(_20144_));
 DFFR_X1 \core.keymem.key_mem[7][64]$_DFFE_PN0P_  (.D(_02461_),
    .RN(net100),
    .CK(clknet_leaf_13_clk),
    .Q(\core.keymem.key_mem[7][64] ),
    .QN(_20143_));
 DFFR_X1 \core.keymem.key_mem[7][65]$_DFFE_PN0P_  (.D(_02462_),
    .RN(net98),
    .CK(clknet_leaf_140_clk),
    .Q(\core.keymem.key_mem[7][65] ),
    .QN(_20142_));
 DFFR_X1 \core.keymem.key_mem[7][66]$_DFFE_PN0P_  (.D(_02463_),
    .RN(net100),
    .CK(clknet_leaf_16_clk),
    .Q(\core.keymem.key_mem[7][66] ),
    .QN(_20141_));
 DFFR_X1 \core.keymem.key_mem[7][67]$_DFFE_PN0P_  (.D(_02464_),
    .RN(net95),
    .CK(clknet_leaf_79_clk),
    .Q(\core.keymem.key_mem[7][67] ),
    .QN(_20140_));
 DFFR_X1 \core.keymem.key_mem[7][68]$_DFFE_PN0P_  (.D(_02465_),
    .RN(net95),
    .CK(clknet_leaf_77_clk),
    .Q(\core.keymem.key_mem[7][68] ),
    .QN(_20139_));
 DFFR_X1 \core.keymem.key_mem[7][69]$_DFFE_PN0P_  (.D(_02466_),
    .RN(net98),
    .CK(clknet_leaf_177_clk),
    .Q(\core.keymem.key_mem[7][69] ),
    .QN(_20138_));
 DFFR_X1 \core.keymem.key_mem[7][6]$_DFFE_PN0P_  (.D(_02467_),
    .RN(net100),
    .CK(clknet_leaf_103_clk),
    .Q(\core.keymem.key_mem[7][6] ),
    .QN(_20137_));
 DFFR_X1 \core.keymem.key_mem[7][70]$_DFFE_PN0P_  (.D(_02468_),
    .RN(net100),
    .CK(clknet_leaf_98_clk),
    .Q(\core.keymem.key_mem[7][70] ),
    .QN(_20136_));
 DFFR_X1 \core.keymem.key_mem[7][71]$_DFFE_PN0P_  (.D(_02469_),
    .RN(net99),
    .CK(clknet_leaf_75_clk),
    .Q(\core.keymem.key_mem[7][71] ),
    .QN(_20135_));
 DFFR_X1 \core.keymem.key_mem[7][72]$_DFFE_PN0P_  (.D(_02470_),
    .RN(net95),
    .CK(clknet_leaf_75_clk),
    .Q(\core.keymem.key_mem[7][72] ),
    .QN(_20134_));
 DFFR_X1 \core.keymem.key_mem[7][73]$_DFFE_PN0P_  (.D(_02471_),
    .RN(net97),
    .CK(clknet_leaf_146_clk),
    .Q(\core.keymem.key_mem[7][73] ),
    .QN(_20133_));
 DFFR_X1 \core.keymem.key_mem[7][74]$_DFFE_PN0P_  (.D(_02472_),
    .RN(net97),
    .CK(clknet_leaf_155_clk),
    .Q(\core.keymem.key_mem[7][74] ),
    .QN(_20132_));
 DFFR_X1 \core.keymem.key_mem[7][75]$_DFFE_PN0P_  (.D(_02473_),
    .RN(net97),
    .CK(clknet_leaf_154_clk),
    .Q(\core.keymem.key_mem[7][75] ),
    .QN(_20131_));
 DFFR_X1 \core.keymem.key_mem[7][76]$_DFFE_PN0P_  (.D(_02474_),
    .RN(net93),
    .CK(clknet_leaf_283_clk),
    .Q(\core.keymem.key_mem[7][76] ),
    .QN(_20130_));
 DFFR_X1 \core.keymem.key_mem[7][77]$_DFFE_PN0P_  (.D(_02475_),
    .RN(net97),
    .CK(clknet_leaf_161_clk),
    .Q(\core.keymem.key_mem[7][77] ),
    .QN(_20129_));
 DFFR_X1 \core.keymem.key_mem[7][78]$_DFFE_PN0P_  (.D(_02476_),
    .RN(net96),
    .CK(clknet_leaf_171_clk),
    .Q(\core.keymem.key_mem[7][78] ),
    .QN(_20128_));
 DFFR_X1 \core.keymem.key_mem[7][79]$_DFFE_PN0P_  (.D(_02477_),
    .RN(net96),
    .CK(clknet_leaf_227_clk),
    .Q(\core.keymem.key_mem[7][79] ),
    .QN(_20127_));
 DFFR_X1 \core.keymem.key_mem[7][7]$_DFFE_PN0P_  (.D(_02478_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[7][7] ),
    .QN(_20126_));
 DFFR_X1 \core.keymem.key_mem[7][80]$_DFFE_PN0P_  (.D(_02479_),
    .RN(net97),
    .CK(clknet_leaf_159_clk),
    .Q(\core.keymem.key_mem[7][80] ),
    .QN(_20125_));
 DFFR_X1 \core.keymem.key_mem[7][81]$_DFFE_PN0P_  (.D(_02480_),
    .RN(net97),
    .CK(clknet_leaf_155_clk),
    .Q(\core.keymem.key_mem[7][81] ),
    .QN(_20124_));
 DFFR_X1 \core.keymem.key_mem[7][82]$_DFFE_PN0P_  (.D(_02481_),
    .RN(net98),
    .CK(clknet_leaf_174_clk),
    .Q(\core.keymem.key_mem[7][82] ),
    .QN(_20123_));
 DFFR_X1 \core.keymem.key_mem[7][83]$_DFFE_PN0P_  (.D(_02482_),
    .RN(net93),
    .CK(clknet_leaf_184_clk),
    .Q(\core.keymem.key_mem[7][83] ),
    .QN(_20122_));
 DFFR_X1 \core.keymem.key_mem[7][84]$_DFFE_PN0P_  (.D(_02483_),
    .RN(net95),
    .CK(clknet_leaf_181_clk),
    .Q(\core.keymem.key_mem[7][84] ),
    .QN(_20121_));
 DFFR_X1 \core.keymem.key_mem[7][85]$_DFFE_PN0P_  (.D(_02484_),
    .RN(net97),
    .CK(clknet_leaf_238_clk),
    .Q(\core.keymem.key_mem[7][85] ),
    .QN(_20120_));
 DFFR_X1 \core.keymem.key_mem[7][86]$_DFFE_PN0P_  (.D(_02485_),
    .RN(net98),
    .CK(clknet_leaf_166_clk),
    .Q(\core.keymem.key_mem[7][86] ),
    .QN(_20119_));
 DFFR_X1 \core.keymem.key_mem[7][87]$_DFFE_PN0P_  (.D(_02486_),
    .RN(net89),
    .CK(clknet_leaf_57_clk),
    .Q(\core.keymem.key_mem[7][87] ),
    .QN(_20118_));
 DFFR_X1 \core.keymem.key_mem[7][88]$_DFFE_PN0P_  (.D(_02487_),
    .RN(net93),
    .CK(clknet_leaf_281_clk),
    .Q(\core.keymem.key_mem[7][88] ),
    .QN(_20117_));
 DFFR_X1 \core.keymem.key_mem[7][89]$_DFFE_PN0P_  (.D(_02488_),
    .RN(net93),
    .CK(clknet_leaf_281_clk),
    .Q(\core.keymem.key_mem[7][89] ),
    .QN(_20116_));
 DFFR_X1 \core.keymem.key_mem[7][8]$_DFFE_PN0P_  (.D(_02489_),
    .RN(net93),
    .CK(clknet_leaf_282_clk),
    .Q(\core.keymem.key_mem[7][8] ),
    .QN(_20115_));
 DFFR_X1 \core.keymem.key_mem[7][90]$_DFFE_PN0P_  (.D(_02490_),
    .RN(net97),
    .CK(clknet_leaf_161_clk),
    .Q(\core.keymem.key_mem[7][90] ),
    .QN(_20114_));
 DFFR_X1 \core.keymem.key_mem[7][91]$_DFFE_PN0P_  (.D(_02491_),
    .RN(net95),
    .CK(clknet_leaf_185_clk),
    .Q(\core.keymem.key_mem[7][91] ),
    .QN(_20113_));
 DFFR_X1 \core.keymem.key_mem[7][92]$_DFFE_PN0P_  (.D(_02492_),
    .RN(net95),
    .CK(clknet_leaf_63_clk),
    .Q(\core.keymem.key_mem[7][92] ),
    .QN(_20112_));
 DFFR_X1 \core.keymem.key_mem[7][93]$_DFFE_PN0P_  (.D(_02493_),
    .RN(net97),
    .CK(clknet_leaf_236_clk),
    .Q(\core.keymem.key_mem[7][93] ),
    .QN(_20111_));
 DFFR_X1 \core.keymem.key_mem[7][94]$_DFFE_PN0P_  (.D(_02494_),
    .RN(net94),
    .CK(clknet_leaf_214_clk),
    .Q(\core.keymem.key_mem[7][94] ),
    .QN(_20110_));
 DFFR_X1 \core.keymem.key_mem[7][95]$_DFFE_PN0P_  (.D(_02495_),
    .RN(net96),
    .CK(clknet_leaf_242_clk),
    .Q(\core.keymem.key_mem[7][95] ),
    .QN(_20109_));
 DFFR_X1 \core.keymem.key_mem[7][96]$_DFFE_PN0P_  (.D(_02496_),
    .RN(net92),
    .CK(clknet_leaf_266_clk),
    .Q(\core.keymem.key_mem[7][96] ),
    .QN(_20108_));
 DFFR_X1 \core.keymem.key_mem[7][97]$_DFFE_PN0P_  (.D(_02497_),
    .RN(net95),
    .CK(clknet_leaf_183_clk),
    .Q(\core.keymem.key_mem[7][97] ),
    .QN(_20107_));
 DFFR_X1 \core.keymem.key_mem[7][98]$_DFFE_PN0P_  (.D(_02498_),
    .RN(net95),
    .CK(clknet_leaf_62_clk),
    .Q(\core.keymem.key_mem[7][98] ),
    .QN(_20106_));
 DFFR_X1 \core.keymem.key_mem[7][99]$_DFFE_PN0P_  (.D(_02499_),
    .RN(net92),
    .CK(clknet_leaf_197_clk),
    .Q(\core.keymem.key_mem[7][99] ),
    .QN(_20105_));
 DFFR_X1 \core.keymem.key_mem[7][9]$_DFFE_PN0P_  (.D(_02500_),
    .RN(net92),
    .CK(clknet_leaf_202_clk),
    .Q(\core.keymem.key_mem[7][9] ),
    .QN(_20104_));
 DFFR_X1 \core.keymem.key_mem[8][0]$_DFFE_PN0P_  (.D(_02501_),
    .RN(net96),
    .CK(clknet_leaf_247_clk),
    .Q(\core.keymem.key_mem[8][0] ),
    .QN(_20103_));
 DFFR_X1 \core.keymem.key_mem[8][100]$_DFFE_PN0P_  (.D(_02502_),
    .RN(net98),
    .CK(clknet_leaf_211_clk),
    .Q(\core.keymem.key_mem[8][100] ),
    .QN(_20102_));
 DFFR_X1 \core.keymem.key_mem[8][101]$_DFFE_PN0P_  (.D(_02503_),
    .RN(net94),
    .CK(clknet_leaf_219_clk),
    .Q(\core.keymem.key_mem[8][101] ),
    .QN(_20101_));
 DFFR_X1 \core.keymem.key_mem[8][102]$_DFFE_PN0P_  (.D(_02504_),
    .RN(net96),
    .CK(clknet_leaf_232_clk),
    .Q(\core.keymem.key_mem[8][102] ),
    .QN(_20100_));
 DFFR_X1 \core.keymem.key_mem[8][103]$_DFFE_PN0P_  (.D(_02505_),
    .RN(net96),
    .CK(clknet_leaf_224_clk),
    .Q(\core.keymem.key_mem[8][103] ),
    .QN(_20099_));
 DFFR_X1 \core.keymem.key_mem[8][104]$_DFFE_PN0P_  (.D(_02506_),
    .RN(net93),
    .CK(clknet_leaf_193_clk),
    .Q(\core.keymem.key_mem[8][104] ),
    .QN(_20098_));
 DFFR_X1 \core.keymem.key_mem[8][105]$_DFFE_PN0P_  (.D(_02507_),
    .RN(net96),
    .CK(clknet_leaf_246_clk),
    .Q(\core.keymem.key_mem[8][105] ),
    .QN(_20097_));
 DFFR_X1 \core.keymem.key_mem[8][106]$_DFFE_PN0P_  (.D(_02508_),
    .RN(net92),
    .CK(clknet_leaf_275_clk),
    .Q(\core.keymem.key_mem[8][106] ),
    .QN(_20096_));
 DFFR_X1 \core.keymem.key_mem[8][107]$_DFFE_PN0P_  (.D(_02509_),
    .RN(net92),
    .CK(clknet_leaf_275_clk),
    .Q(\core.keymem.key_mem[8][107] ),
    .QN(_20095_));
 DFFR_X1 \core.keymem.key_mem[8][108]$_DFFE_PN0P_  (.D(_02510_),
    .RN(net91),
    .CK(clknet_leaf_278_clk),
    .Q(\core.keymem.key_mem[8][108] ),
    .QN(_20094_));
 DFFR_X1 \core.keymem.key_mem[8][109]$_DFFE_PN0P_  (.D(_02511_),
    .RN(net94),
    .CK(clknet_leaf_269_clk),
    .Q(\core.keymem.key_mem[8][109] ),
    .QN(_20093_));
 DFFR_X1 \core.keymem.key_mem[8][10]$_DFFE_PN0P_  (.D(_02512_),
    .RN(net98),
    .CK(clknet_leaf_188_clk),
    .Q(\core.keymem.key_mem[8][10] ),
    .QN(_20092_));
 DFFR_X1 \core.keymem.key_mem[8][110]$_DFFE_PN0P_  (.D(_02513_),
    .RN(net96),
    .CK(clknet_leaf_221_clk),
    .Q(\core.keymem.key_mem[8][110] ),
    .QN(_20091_));
 DFFR_X1 \core.keymem.key_mem[8][111]$_DFFE_PN0P_  (.D(_02514_),
    .RN(net96),
    .CK(clknet_leaf_226_clk),
    .Q(\core.keymem.key_mem[8][111] ),
    .QN(_20090_));
 DFFR_X1 \core.keymem.key_mem[8][112]$_DFFE_PN0P_  (.D(_02515_),
    .RN(net94),
    .CK(clknet_leaf_261_clk),
    .Q(\core.keymem.key_mem[8][112] ),
    .QN(_20089_));
 DFFR_X1 \core.keymem.key_mem[8][113]$_DFFE_PN0P_  (.D(_02516_),
    .RN(net92),
    .CK(clknet_leaf_273_clk),
    .Q(\core.keymem.key_mem[8][113] ),
    .QN(_20088_));
 DFFR_X1 \core.keymem.key_mem[8][114]$_DFFE_PN0P_  (.D(_02517_),
    .RN(net91),
    .CK(clknet_leaf_279_clk),
    .Q(\core.keymem.key_mem[8][114] ),
    .QN(_20087_));
 DFFR_X1 \core.keymem.key_mem[8][115]$_DFFE_PN0P_  (.D(_02518_),
    .RN(net92),
    .CK(clknet_leaf_278_clk),
    .Q(\core.keymem.key_mem[8][115] ),
    .QN(_20086_));
 DFFR_X1 \core.keymem.key_mem[8][116]$_DFFE_PN0P_  (.D(_02519_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[8][116] ),
    .QN(_20085_));
 DFFR_X1 \core.keymem.key_mem[8][117]$_DFFE_PN0P_  (.D(_02520_),
    .RN(net96),
    .CK(clknet_leaf_222_clk),
    .Q(\core.keymem.key_mem[8][117] ),
    .QN(_20084_));
 DFFR_X1 \core.keymem.key_mem[8][118]$_DFFE_PN0P_  (.D(_02521_),
    .RN(net96),
    .CK(clknet_leaf_243_clk),
    .Q(\core.keymem.key_mem[8][118] ),
    .QN(_20083_));
 DFFR_X1 \core.keymem.key_mem[8][119]$_DFFE_PN0P_  (.D(_02522_),
    .RN(net94),
    .CK(clknet_leaf_217_clk),
    .Q(\core.keymem.key_mem[8][119] ),
    .QN(_20082_));
 DFFR_X1 \core.keymem.key_mem[8][11]$_DFFE_PN0P_  (.D(_02523_),
    .RN(net95),
    .CK(clknet_leaf_61_clk),
    .Q(\core.keymem.key_mem[8][11] ),
    .QN(_20081_));
 DFFR_X1 \core.keymem.key_mem[8][120]$_DFFE_PN0P_  (.D(_02524_),
    .RN(net93),
    .CK(clknet_leaf_206_clk),
    .Q(\core.keymem.key_mem[8][120] ),
    .QN(_20080_));
 DFFR_X1 \core.keymem.key_mem[8][121]$_DFFE_PN0P_  (.D(_02525_),
    .RN(net94),
    .CK(clknet_leaf_216_clk),
    .Q(\core.keymem.key_mem[8][121] ),
    .QN(_20079_));
 DFFR_X1 \core.keymem.key_mem[8][122]$_DFFE_PN0P_  (.D(_02526_),
    .RN(net97),
    .CK(clknet_leaf_160_clk),
    .Q(\core.keymem.key_mem[8][122] ),
    .QN(_20078_));
 DFFR_X1 \core.keymem.key_mem[8][123]$_DFFE_PN0P_  (.D(_02527_),
    .RN(net93),
    .CK(clknet_leaf_195_clk),
    .Q(\core.keymem.key_mem[8][123] ),
    .QN(_20077_));
 DFFR_X1 \core.keymem.key_mem[8][124]$_DFFE_PN0P_  (.D(_02528_),
    .RN(net93),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[8][124] ),
    .QN(_20076_));
 DFFR_X1 \core.keymem.key_mem[8][125]$_DFFE_PN0P_  (.D(_02529_),
    .RN(net97),
    .CK(clknet_leaf_231_clk),
    .Q(\core.keymem.key_mem[8][125] ),
    .QN(_20075_));
 DFFR_X1 \core.keymem.key_mem[8][126]$_DFFE_PN0P_  (.D(_02530_),
    .RN(net98),
    .CK(clknet_leaf_168_clk),
    .Q(\core.keymem.key_mem[8][126] ),
    .QN(_20074_));
 DFFR_X1 \core.keymem.key_mem[8][127]$_DFFE_PN0P_  (.D(_02531_),
    .RN(net97),
    .CK(clknet_leaf_235_clk),
    .Q(\core.keymem.key_mem[8][127] ),
    .QN(_20073_));
 DFFR_X1 \core.keymem.key_mem[8][12]$_DFFE_PN0P_  (.D(_02532_),
    .RN(net93),
    .CK(clknet_leaf_206_clk),
    .Q(\core.keymem.key_mem[8][12] ),
    .QN(_20072_));
 DFFR_X1 \core.keymem.key_mem[8][13]$_DFFE_PN0P_  (.D(_02533_),
    .RN(net87),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[8][13] ),
    .QN(_20071_));
 DFFR_X1 \core.keymem.key_mem[8][14]$_DFFE_PN0P_  (.D(_02534_),
    .RN(net94),
    .CK(clknet_leaf_211_clk),
    .Q(\core.keymem.key_mem[8][14] ),
    .QN(_20070_));
 DFFR_X1 \core.keymem.key_mem[8][15]$_DFFE_PN0P_  (.D(_02535_),
    .RN(net96),
    .CK(clknet_leaf_165_clk),
    .Q(\core.keymem.key_mem[8][15] ),
    .QN(_20069_));
 DFFR_X1 \core.keymem.key_mem[8][16]$_DFFE_PN0P_  (.D(_02536_),
    .RN(net89),
    .CK(clknet_leaf_34_clk),
    .Q(\core.keymem.key_mem[8][16] ),
    .QN(_20068_));
 DFFR_X1 \core.keymem.key_mem[8][17]$_DFFE_PN0P_  (.D(_02537_),
    .RN(net98),
    .CK(clknet_leaf_168_clk),
    .Q(\core.keymem.key_mem[8][17] ),
    .QN(_20067_));
 DFFR_X1 \core.keymem.key_mem[8][18]$_DFFE_PN0P_  (.D(_02538_),
    .RN(net82),
    .CK(clknet_leaf_35_clk),
    .Q(\core.keymem.key_mem[8][18] ),
    .QN(_20066_));
 DFFR_X1 \core.keymem.key_mem[8][19]$_DFFE_PN0P_  (.D(_02539_),
    .RN(net89),
    .CK(clknet_leaf_64_clk),
    .Q(\core.keymem.key_mem[8][19] ),
    .QN(_20065_));
 DFFR_X1 \core.keymem.key_mem[8][1]$_DFFE_PN0P_  (.D(_02540_),
    .RN(net89),
    .CK(clknet_leaf_26_clk),
    .Q(\core.keymem.key_mem[8][1] ),
    .QN(_20064_));
 DFFR_X1 \core.keymem.key_mem[8][20]$_DFFE_PN0P_  (.D(_02541_),
    .RN(net89),
    .CK(clknet_leaf_95_clk),
    .Q(\core.keymem.key_mem[8][20] ),
    .QN(_20063_));
 DFFR_X1 \core.keymem.key_mem[8][21]$_DFFE_PN0P_  (.D(_02542_),
    .RN(net85),
    .CK(clknet_leaf_67_clk),
    .Q(\core.keymem.key_mem[8][21] ),
    .QN(_20062_));
 DFFR_X1 \core.keymem.key_mem[8][22]$_DFFE_PN0P_  (.D(_02543_),
    .RN(net96),
    .CK(clknet_leaf_222_clk),
    .Q(\core.keymem.key_mem[8][22] ),
    .QN(_20061_));
 DFFR_X1 \core.keymem.key_mem[8][23]$_DFFE_PN0P_  (.D(_02544_),
    .RN(net89),
    .CK(clknet_leaf_56_clk),
    .Q(\core.keymem.key_mem[8][23] ),
    .QN(_20060_));
 DFFR_X1 \core.keymem.key_mem[8][24]$_DFFE_PN0P_  (.D(_02545_),
    .RN(net85),
    .CK(clknet_leaf_49_clk),
    .Q(\core.keymem.key_mem[8][24] ),
    .QN(_20059_));
 DFFR_X1 \core.keymem.key_mem[8][25]$_DFFE_PN0P_  (.D(_02546_),
    .RN(net85),
    .CK(clknet_leaf_50_clk),
    .Q(\core.keymem.key_mem[8][25] ),
    .QN(_20058_));
 DFFR_X1 \core.keymem.key_mem[8][26]$_DFFE_PN0P_  (.D(_02547_),
    .RN(net89),
    .CK(clknet_leaf_91_clk),
    .Q(\core.keymem.key_mem[8][26] ),
    .QN(_20057_));
 DFFR_X1 \core.keymem.key_mem[8][27]$_DFFE_PN0P_  (.D(_02548_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[8][27] ),
    .QN(_20056_));
 DFFR_X1 \core.keymem.key_mem[8][28]$_DFFE_PN0P_  (.D(_02549_),
    .RN(net16),
    .CK(clknet_leaf_125_clk),
    .Q(\core.keymem.key_mem[8][28] ),
    .QN(_20055_));
 DFFR_X1 \core.keymem.key_mem[8][29]$_DFFE_PN0P_  (.D(_02550_),
    .RN(net16),
    .CK(clknet_leaf_149_clk),
    .Q(\core.keymem.key_mem[8][29] ),
    .QN(_20054_));
 DFFR_X1 \core.keymem.key_mem[8][2]$_DFFE_PN0P_  (.D(_02551_),
    .RN(net95),
    .CK(clknet_leaf_62_clk),
    .Q(\core.keymem.key_mem[8][2] ),
    .QN(_20053_));
 DFFR_X1 \core.keymem.key_mem[8][30]$_DFFE_PN0P_  (.D(_02552_),
    .RN(net98),
    .CK(clknet_leaf_144_clk),
    .Q(\core.keymem.key_mem[8][30] ),
    .QN(_20052_));
 DFFR_X1 \core.keymem.key_mem[8][31]$_DFFE_PN0P_  (.D(_02553_),
    .RN(net16),
    .CK(clknet_leaf_138_clk),
    .Q(\core.keymem.key_mem[8][31] ),
    .QN(_20051_));
 DFFR_X1 \core.keymem.key_mem[8][32]$_DFFE_PN0P_  (.D(_02554_),
    .RN(net100),
    .CK(clknet_leaf_116_clk),
    .Q(\core.keymem.key_mem[8][32] ),
    .QN(_20050_));
 DFFR_X1 \core.keymem.key_mem[8][33]$_DFFE_PN0P_  (.D(_02555_),
    .RN(net99),
    .CK(clknet_leaf_111_clk),
    .Q(\core.keymem.key_mem[8][33] ),
    .QN(_20049_));
 DFFR_X1 \core.keymem.key_mem[8][34]$_DFFE_PN0P_  (.D(_02556_),
    .RN(net16),
    .CK(clknet_leaf_136_clk),
    .Q(\core.keymem.key_mem[8][34] ),
    .QN(_20048_));
 DFFR_X1 \core.keymem.key_mem[8][35]$_DFFE_PN0P_  (.D(_02557_),
    .RN(net99),
    .CK(clknet_leaf_122_clk),
    .Q(\core.keymem.key_mem[8][35] ),
    .QN(_20047_));
 DFFR_X1 \core.keymem.key_mem[8][36]$_DFFE_PN0P_  (.D(_02558_),
    .RN(net88),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[8][36] ),
    .QN(_20046_));
 DFFR_X1 \core.keymem.key_mem[8][37]$_DFFE_PN0P_  (.D(_02559_),
    .RN(net89),
    .CK(clknet_leaf_85_clk),
    .Q(\core.keymem.key_mem[8][37] ),
    .QN(_20045_));
 DFFR_X1 \core.keymem.key_mem[8][38]$_DFFE_PN0P_  (.D(_02560_),
    .RN(net99),
    .CK(clknet_leaf_123_clk),
    .Q(\core.keymem.key_mem[8][38] ),
    .QN(_20044_));
 DFFR_X1 \core.keymem.key_mem[8][39]$_DFFE_PN0P_  (.D(_02561_),
    .RN(net89),
    .CK(clknet_leaf_85_clk),
    .Q(\core.keymem.key_mem[8][39] ),
    .QN(_20043_));
 DFFR_X1 \core.keymem.key_mem[8][3]$_DFFE_PN0P_  (.D(_02562_),
    .RN(net85),
    .CK(clknet_leaf_30_clk),
    .Q(\core.keymem.key_mem[8][3] ),
    .QN(_20042_));
 DFFR_X1 \core.keymem.key_mem[8][40]$_DFFE_PN0P_  (.D(_02563_),
    .RN(net85),
    .CK(clknet_leaf_30_clk),
    .Q(\core.keymem.key_mem[8][40] ),
    .QN(_20041_));
 DFFR_X1 \core.keymem.key_mem[8][41]$_DFFE_PN0P_  (.D(_02564_),
    .RN(net89),
    .CK(clknet_leaf_115_clk),
    .Q(\core.keymem.key_mem[8][41] ),
    .QN(_20040_));
 DFFR_X1 \core.keymem.key_mem[8][42]$_DFFE_PN0P_  (.D(_02565_),
    .RN(net100),
    .CK(clknet_leaf_110_clk),
    .Q(\core.keymem.key_mem[8][42] ),
    .QN(_20039_));
 DFFR_X1 \core.keymem.key_mem[8][43]$_DFFE_PN0P_  (.D(_02566_),
    .RN(net85),
    .CK(clknet_leaf_47_clk),
    .Q(\core.keymem.key_mem[8][43] ),
    .QN(_20038_));
 DFFR_X1 \core.keymem.key_mem[8][44]$_DFFE_PN0P_  (.D(_02567_),
    .RN(net100),
    .CK(clknet_leaf_114_clk),
    .Q(\core.keymem.key_mem[8][44] ),
    .QN(_20037_));
 DFFR_X1 \core.keymem.key_mem[8][45]$_DFFE_PN0P_  (.D(_02568_),
    .RN(net99),
    .CK(clknet_leaf_69_clk),
    .Q(\core.keymem.key_mem[8][45] ),
    .QN(_20036_));
 DFFR_X1 \core.keymem.key_mem[8][46]$_DFFE_PN0P_  (.D(_02569_),
    .RN(net99),
    .CK(clknet_leaf_79_clk),
    .Q(\core.keymem.key_mem[8][46] ),
    .QN(_20035_));
 DFFR_X1 \core.keymem.key_mem[8][47]$_DFFE_PN0P_  (.D(_02570_),
    .RN(net98),
    .CK(clknet_leaf_175_clk),
    .Q(\core.keymem.key_mem[8][47] ),
    .QN(_20034_));
 DFFR_X1 \core.keymem.key_mem[8][48]$_DFFE_PN0P_  (.D(_02571_),
    .RN(net95),
    .CK(clknet_leaf_119_clk),
    .Q(\core.keymem.key_mem[8][48] ),
    .QN(_20033_));
 DFFR_X1 \core.keymem.key_mem[8][49]$_DFFE_PN0P_  (.D(_02572_),
    .RN(net99),
    .CK(clknet_leaf_78_clk),
    .Q(\core.keymem.key_mem[8][49] ),
    .QN(_20032_));
 DFFR_X1 \core.keymem.key_mem[8][4]$_DFFE_PN0P_  (.D(_02573_),
    .RN(net100),
    .CK(clknet_leaf_105_clk),
    .Q(\core.keymem.key_mem[8][4] ),
    .QN(_20031_));
 DFFR_X1 \core.keymem.key_mem[8][50]$_DFFE_PN0P_  (.D(_02574_),
    .RN(net98),
    .CK(clknet_leaf_137_clk),
    .Q(\core.keymem.key_mem[8][50] ),
    .QN(_20030_));
 DFFR_X1 \core.keymem.key_mem[8][51]$_DFFE_PN0P_  (.D(_02575_),
    .RN(net100),
    .CK(clknet_leaf_129_clk),
    .Q(\core.keymem.key_mem[8][51] ),
    .QN(_20029_));
 DFFR_X1 \core.keymem.key_mem[8][52]$_DFFE_PN0P_  (.D(_02576_),
    .RN(net99),
    .CK(clknet_leaf_79_clk),
    .Q(\core.keymem.key_mem[8][52] ),
    .QN(_20028_));
 DFFR_X1 \core.keymem.key_mem[8][53]$_DFFE_PN0P_  (.D(_02577_),
    .RN(net98),
    .CK(clknet_leaf_175_clk),
    .Q(\core.keymem.key_mem[8][53] ),
    .QN(_20027_));
 DFFR_X1 \core.keymem.key_mem[8][54]$_DFFE_PN0P_  (.D(_02578_),
    .RN(net98),
    .CK(clknet_leaf_142_clk),
    .Q(\core.keymem.key_mem[8][54] ),
    .QN(_20026_));
 DFFR_X1 \core.keymem.key_mem[8][55]$_DFFE_PN0P_  (.D(_02579_),
    .RN(net16),
    .CK(clknet_leaf_136_clk),
    .Q(\core.keymem.key_mem[8][55] ),
    .QN(_20025_));
 DFFR_X1 \core.keymem.key_mem[8][56]$_DFFE_PN0P_  (.D(_02580_),
    .RN(net16),
    .CK(clknet_leaf_134_clk),
    .Q(\core.keymem.key_mem[8][56] ),
    .QN(_20024_));
 DFFR_X1 \core.keymem.key_mem[8][57]$_DFFE_PN0P_  (.D(_02581_),
    .RN(net100),
    .CK(clknet_leaf_110_clk),
    .Q(\core.keymem.key_mem[8][57] ),
    .QN(_20023_));
 DFFR_X1 \core.keymem.key_mem[8][58]$_DFFE_PN0P_  (.D(_02582_),
    .RN(net100),
    .CK(clknet_leaf_106_clk),
    .Q(\core.keymem.key_mem[8][58] ),
    .QN(_20022_));
 DFFR_X1 \core.keymem.key_mem[8][59]$_DFFE_PN0P_  (.D(_02583_),
    .RN(net100),
    .CK(clknet_leaf_17_clk),
    .Q(\core.keymem.key_mem[8][59] ),
    .QN(_20021_));
 DFFR_X1 \core.keymem.key_mem[8][5]$_DFFE_PN0P_  (.D(_02584_),
    .RN(net100),
    .CK(clknet_leaf_18_clk),
    .Q(\core.keymem.key_mem[8][5] ),
    .QN(_20020_));
 DFFR_X1 \core.keymem.key_mem[8][60]$_DFFE_PN0P_  (.D(_02585_),
    .RN(net82),
    .CK(clknet_leaf_13_clk),
    .Q(\core.keymem.key_mem[8][60] ),
    .QN(_20019_));
 DFFR_X1 \core.keymem.key_mem[8][61]$_DFFE_PN0P_  (.D(_02586_),
    .RN(net88),
    .CK(clknet_leaf_94_clk),
    .Q(\core.keymem.key_mem[8][61] ),
    .QN(_20018_));
 DFFR_X1 \core.keymem.key_mem[8][62]$_DFFE_PN0P_  (.D(_02587_),
    .RN(net100),
    .CK(clknet_leaf_99_clk),
    .Q(\core.keymem.key_mem[8][62] ),
    .QN(_20017_));
 DFFR_X1 \core.keymem.key_mem[8][63]$_DFFE_PN0P_  (.D(_02588_),
    .RN(net100),
    .CK(clknet_leaf_20_clk),
    .Q(\core.keymem.key_mem[8][63] ),
    .QN(_20016_));
 DFFR_X1 \core.keymem.key_mem[8][64]$_DFFE_PN0P_  (.D(_02589_),
    .RN(net82),
    .CK(clknet_leaf_13_clk),
    .Q(\core.keymem.key_mem[8][64] ),
    .QN(_20015_));
 DFFR_X1 \core.keymem.key_mem[8][65]$_DFFE_PN0P_  (.D(_02590_),
    .RN(net99),
    .CK(clknet_leaf_120_clk),
    .Q(\core.keymem.key_mem[8][65] ),
    .QN(_20014_));
 DFFR_X1 \core.keymem.key_mem[8][66]$_DFFE_PN0P_  (.D(_02591_),
    .RN(net100),
    .CK(clknet_leaf_16_clk),
    .Q(\core.keymem.key_mem[8][66] ),
    .QN(_20013_));
 DFFR_X1 \core.keymem.key_mem[8][67]$_DFFE_PN0P_  (.D(_02592_),
    .RN(net99),
    .CK(clknet_leaf_74_clk),
    .Q(\core.keymem.key_mem[8][67] ),
    .QN(_20012_));
 DFFR_X1 \core.keymem.key_mem[8][68]$_DFFE_PN0P_  (.D(_02593_),
    .RN(net95),
    .CK(clknet_leaf_78_clk),
    .Q(\core.keymem.key_mem[8][68] ),
    .QN(_20011_));
 DFFR_X1 \core.keymem.key_mem[8][69]$_DFFE_PN0P_  (.D(_02594_),
    .RN(net98),
    .CK(clknet_leaf_177_clk),
    .Q(\core.keymem.key_mem[8][69] ),
    .QN(_20010_));
 DFFR_X1 \core.keymem.key_mem[8][6]$_DFFE_PN0P_  (.D(_02595_),
    .RN(net100),
    .CK(clknet_leaf_101_clk),
    .Q(\core.keymem.key_mem[8][6] ),
    .QN(_20009_));
 DFFR_X1 \core.keymem.key_mem[8][70]$_DFFE_PN0P_  (.D(_02596_),
    .RN(net100),
    .CK(clknet_leaf_100_clk),
    .Q(\core.keymem.key_mem[8][70] ),
    .QN(_20008_));
 DFFR_X1 \core.keymem.key_mem[8][71]$_DFFE_PN0P_  (.D(_02597_),
    .RN(net99),
    .CK(clknet_leaf_75_clk),
    .Q(\core.keymem.key_mem[8][71] ),
    .QN(_20007_));
 DFFR_X1 \core.keymem.key_mem[8][72]$_DFFE_PN0P_  (.D(_02598_),
    .RN(net95),
    .CK(clknet_leaf_73_clk),
    .Q(\core.keymem.key_mem[8][72] ),
    .QN(_20006_));
 DFFR_X1 \core.keymem.key_mem[8][73]$_DFFE_PN0P_  (.D(_02599_),
    .RN(net97),
    .CK(clknet_leaf_146_clk),
    .Q(\core.keymem.key_mem[8][73] ),
    .QN(_20005_));
 DFFR_X1 \core.keymem.key_mem[8][74]$_DFFE_PN0P_  (.D(_02600_),
    .RN(net97),
    .CK(clknet_leaf_154_clk),
    .Q(\core.keymem.key_mem[8][74] ),
    .QN(_20004_));
 DFFR_X1 \core.keymem.key_mem[8][75]$_DFFE_PN0P_  (.D(_02601_),
    .RN(net97),
    .CK(clknet_leaf_154_clk),
    .Q(\core.keymem.key_mem[8][75] ),
    .QN(_20003_));
 DFFR_X1 \core.keymem.key_mem[8][76]$_DFFE_PN0P_  (.D(_02602_),
    .RN(net93),
    .CK(clknet_leaf_377_clk),
    .Q(\core.keymem.key_mem[8][76] ),
    .QN(_20002_));
 DFFR_X1 \core.keymem.key_mem[8][77]$_DFFE_PN0P_  (.D(_02603_),
    .RN(net97),
    .CK(clknet_leaf_160_clk),
    .Q(\core.keymem.key_mem[8][77] ),
    .QN(_20001_));
 DFFR_X1 \core.keymem.key_mem[8][78]$_DFFE_PN0P_  (.D(_02604_),
    .RN(net97),
    .CK(clknet_leaf_172_clk),
    .Q(\core.keymem.key_mem[8][78] ),
    .QN(_20000_));
 DFFR_X1 \core.keymem.key_mem[8][79]$_DFFE_PN0P_  (.D(_02605_),
    .RN(net98),
    .CK(clknet_leaf_230_clk),
    .Q(\core.keymem.key_mem[8][79] ),
    .QN(_19999_));
 DFFR_X1 \core.keymem.key_mem[8][7]$_DFFE_PN0P_  (.D(_02606_),
    .RN(net98),
    .CK(clknet_leaf_175_clk),
    .Q(\core.keymem.key_mem[8][7] ),
    .QN(_19998_));
 DFFR_X1 \core.keymem.key_mem[8][80]$_DFFE_PN0P_  (.D(_02607_),
    .RN(net97),
    .CK(clknet_leaf_159_clk),
    .Q(\core.keymem.key_mem[8][80] ),
    .QN(_19997_));
 DFFR_X1 \core.keymem.key_mem[8][81]$_DFFE_PN0P_  (.D(_02608_),
    .RN(net97),
    .CK(clknet_leaf_155_clk),
    .Q(\core.keymem.key_mem[8][81] ),
    .QN(_19996_));
 DFFR_X1 \core.keymem.key_mem[8][82]$_DFFE_PN0P_  (.D(_02609_),
    .RN(net98),
    .CK(clknet_leaf_174_clk),
    .Q(\core.keymem.key_mem[8][82] ),
    .QN(_19995_));
 DFFR_X2 \core.keymem.key_mem[8][83]$_DFFE_PN0P_  (.D(_02610_),
    .RN(net95),
    .CK(clknet_leaf_181_clk),
    .Q(\core.keymem.key_mem[8][83] ),
    .QN(_19994_));
 DFFR_X1 \core.keymem.key_mem[8][84]$_DFFE_PN0P_  (.D(_02611_),
    .RN(net95),
    .CK(clknet_leaf_181_clk),
    .Q(\core.keymem.key_mem[8][84] ),
    .QN(_19993_));
 DFFR_X1 \core.keymem.key_mem[8][85]$_DFFE_PN0P_  (.D(_02612_),
    .RN(net97),
    .CK(clknet_leaf_237_clk),
    .Q(\core.keymem.key_mem[8][85] ),
    .QN(_19992_));
 DFFR_X1 \core.keymem.key_mem[8][86]$_DFFE_PN0P_  (.D(_02613_),
    .RN(net97),
    .CK(clknet_leaf_162_clk),
    .Q(\core.keymem.key_mem[8][86] ),
    .QN(_19991_));
 DFFR_X1 \core.keymem.key_mem[8][87]$_DFFE_PN0P_  (.D(_02614_),
    .RN(net89),
    .CK(clknet_leaf_56_clk),
    .Q(\core.keymem.key_mem[8][87] ),
    .QN(_19990_));
 DFFR_X1 \core.keymem.key_mem[8][88]$_DFFE_PN0P_  (.D(_02615_),
    .RN(net93),
    .CK(clknet_leaf_282_clk),
    .Q(\core.keymem.key_mem[8][88] ),
    .QN(_19989_));
 DFFR_X1 \core.keymem.key_mem[8][89]$_DFFE_PN0P_  (.D(_02616_),
    .RN(net93),
    .CK(clknet_leaf_281_clk),
    .Q(\core.keymem.key_mem[8][89] ),
    .QN(_19988_));
 DFFR_X1 \core.keymem.key_mem[8][8]$_DFFE_PN0P_  (.D(_02617_),
    .RN(net93),
    .CK(clknet_leaf_282_clk),
    .Q(\core.keymem.key_mem[8][8] ),
    .QN(_19987_));
 DFFR_X1 \core.keymem.key_mem[8][90]$_DFFE_PN0P_  (.D(_02618_),
    .RN(net97),
    .CK(clknet_leaf_162_clk),
    .Q(\core.keymem.key_mem[8][90] ),
    .QN(_19986_));
 DFFR_X1 \core.keymem.key_mem[8][91]$_DFFE_PN0P_  (.D(_02619_),
    .RN(net95),
    .CK(clknet_leaf_181_clk),
    .Q(\core.keymem.key_mem[8][91] ),
    .QN(_19985_));
 DFFR_X1 \core.keymem.key_mem[8][92]$_DFFE_PN0P_  (.D(_02620_),
    .RN(net95),
    .CK(clknet_leaf_63_clk),
    .Q(\core.keymem.key_mem[8][92] ),
    .QN(_19984_));
 DFFR_X1 \core.keymem.key_mem[8][93]$_DFFE_PN0P_  (.D(_02621_),
    .RN(net94),
    .CK(clknet_leaf_189_clk),
    .Q(\core.keymem.key_mem[8][93] ),
    .QN(_19983_));
 DFFR_X1 \core.keymem.key_mem[8][94]$_DFFE_PN0P_  (.D(_02622_),
    .RN(net94),
    .CK(clknet_leaf_214_clk),
    .Q(\core.keymem.key_mem[8][94] ),
    .QN(_19982_));
 DFFR_X1 \core.keymem.key_mem[8][95]$_DFFE_PN0P_  (.D(_02623_),
    .RN(net96),
    .CK(clknet_leaf_234_clk),
    .Q(\core.keymem.key_mem[8][95] ),
    .QN(_19981_));
 DFFR_X1 \core.keymem.key_mem[8][96]$_DFFE_PN0P_  (.D(_02624_),
    .RN(net92),
    .CK(clknet_leaf_204_clk),
    .Q(\core.keymem.key_mem[8][96] ),
    .QN(_19980_));
 DFFR_X1 \core.keymem.key_mem[8][97]$_DFFE_PN0P_  (.D(_02625_),
    .RN(net95),
    .CK(clknet_leaf_62_clk),
    .Q(\core.keymem.key_mem[8][97] ),
    .QN(_19979_));
 DFFR_X1 \core.keymem.key_mem[8][98]$_DFFE_PN0P_  (.D(_02626_),
    .RN(net95),
    .CK(clknet_leaf_62_clk),
    .Q(\core.keymem.key_mem[8][98] ),
    .QN(_19978_));
 DFFR_X1 \core.keymem.key_mem[8][99]$_DFFE_PN0P_  (.D(_02627_),
    .RN(net92),
    .CK(clknet_leaf_202_clk),
    .Q(\core.keymem.key_mem[8][99] ),
    .QN(_19977_));
 DFFR_X1 \core.keymem.key_mem[8][9]$_DFFE_PN0P_  (.D(_02628_),
    .RN(net92),
    .CK(clknet_leaf_202_clk),
    .Q(\core.keymem.key_mem[8][9] ),
    .QN(_19976_));
 DFFR_X1 \core.keymem.key_mem[9][0]$_DFFE_PN0P_  (.D(_02629_),
    .RN(net94),
    .CK(clknet_leaf_220_clk),
    .Q(\core.keymem.key_mem[9][0] ),
    .QN(_19975_));
 DFFR_X1 \core.keymem.key_mem[9][100]$_DFFE_PN0P_  (.D(_02630_),
    .RN(net94),
    .CK(clknet_leaf_209_clk),
    .Q(\core.keymem.key_mem[9][100] ),
    .QN(_19974_));
 DFFR_X1 \core.keymem.key_mem[9][101]$_DFFE_PN0P_  (.D(_02631_),
    .RN(net94),
    .CK(clknet_leaf_218_clk),
    .Q(\core.keymem.key_mem[9][101] ),
    .QN(_19973_));
 DFFR_X1 \core.keymem.key_mem[9][102]$_DFFE_PN0P_  (.D(_02632_),
    .RN(net96),
    .CK(clknet_leaf_231_clk),
    .Q(\core.keymem.key_mem[9][102] ),
    .QN(_19972_));
 DFFR_X1 \core.keymem.key_mem[9][103]$_DFFE_PN0P_  (.D(_02633_),
    .RN(net96),
    .CK(clknet_leaf_224_clk),
    .Q(\core.keymem.key_mem[9][103] ),
    .QN(_19971_));
 DFFR_X1 \core.keymem.key_mem[9][104]$_DFFE_PN0P_  (.D(_02634_),
    .RN(net93),
    .CK(clknet_leaf_196_clk),
    .Q(\core.keymem.key_mem[9][104] ),
    .QN(_19970_));
 DFFR_X1 \core.keymem.key_mem[9][105]$_DFFE_PN0P_  (.D(_02635_),
    .RN(net96),
    .CK(clknet_leaf_249_clk),
    .Q(\core.keymem.key_mem[9][105] ),
    .QN(_19969_));
 DFFR_X1 \core.keymem.key_mem[9][106]$_DFFE_PN0P_  (.D(_02636_),
    .RN(net92),
    .CK(clknet_leaf_268_clk),
    .Q(\core.keymem.key_mem[9][106] ),
    .QN(_19968_));
 DFFR_X1 \core.keymem.key_mem[9][107]$_DFFE_PN0P_  (.D(_02637_),
    .RN(net92),
    .CK(clknet_leaf_272_clk),
    .Q(\core.keymem.key_mem[9][107] ),
    .QN(_19967_));
 DFFR_X1 \core.keymem.key_mem[9][108]$_DFFE_PN0P_  (.D(_02638_),
    .RN(net92),
    .CK(clknet_leaf_203_clk),
    .Q(\core.keymem.key_mem[9][108] ),
    .QN(_19966_));
 DFFR_X1 \core.keymem.key_mem[9][109]$_DFFE_PN0P_  (.D(_02639_),
    .RN(net92),
    .CK(clknet_leaf_269_clk),
    .Q(\core.keymem.key_mem[9][109] ),
    .QN(_19965_));
 DFFR_X1 \core.keymem.key_mem[9][10]$_DFFE_PN0P_  (.D(_02640_),
    .RN(net95),
    .CK(clknet_leaf_187_clk),
    .Q(\core.keymem.key_mem[9][10] ),
    .QN(_19964_));
 DFFR_X1 \core.keymem.key_mem[9][110]$_DFFE_PN0P_  (.D(_02641_),
    .RN(net96),
    .CK(clknet_leaf_249_clk),
    .Q(\core.keymem.key_mem[9][110] ),
    .QN(_19963_));
 DFFR_X1 \core.keymem.key_mem[9][111]$_DFFE_PN0P_  (.D(_02642_),
    .RN(net96),
    .CK(clknet_leaf_227_clk),
    .Q(\core.keymem.key_mem[9][111] ),
    .QN(_19962_));
 DFFR_X1 \core.keymem.key_mem[9][112]$_DFFE_PN0P_  (.D(_02643_),
    .RN(net94),
    .CK(clknet_leaf_263_clk),
    .Q(\core.keymem.key_mem[9][112] ),
    .QN(_19961_));
 DFFR_X1 \core.keymem.key_mem[9][113]$_DFFE_PN0P_  (.D(_02644_),
    .RN(net91),
    .CK(clknet_leaf_288_clk),
    .Q(\core.keymem.key_mem[9][113] ),
    .QN(_19960_));
 DFFR_X1 \core.keymem.key_mem[9][114]$_DFFE_PN0P_  (.D(_02645_),
    .RN(net91),
    .CK(clknet_leaf_288_clk),
    .Q(\core.keymem.key_mem[9][114] ),
    .QN(_19959_));
 DFFR_X1 \core.keymem.key_mem[9][115]$_DFFE_PN0P_  (.D(_02646_),
    .RN(net92),
    .CK(clknet_leaf_276_clk),
    .Q(\core.keymem.key_mem[9][115] ),
    .QN(_19958_));
 DFFR_X1 \core.keymem.key_mem[9][116]$_DFFE_PN0P_  (.D(_02647_),
    .RN(net92),
    .CK(clknet_leaf_265_clk),
    .Q(\core.keymem.key_mem[9][116] ),
    .QN(_19957_));
 DFFR_X1 \core.keymem.key_mem[9][117]$_DFFE_PN0P_  (.D(_02648_),
    .RN(net96),
    .CK(clknet_leaf_226_clk),
    .Q(\core.keymem.key_mem[9][117] ),
    .QN(_19956_));
 DFFR_X1 \core.keymem.key_mem[9][118]$_DFFE_PN0P_  (.D(_02649_),
    .RN(net97),
    .CK(clknet_leaf_235_clk),
    .Q(\core.keymem.key_mem[9][118] ),
    .QN(_19955_));
 DFFR_X1 \core.keymem.key_mem[9][119]$_DFFE_PN0P_  (.D(_02650_),
    .RN(net94),
    .CK(clknet_leaf_220_clk),
    .Q(\core.keymem.key_mem[9][119] ),
    .QN(_19954_));
 DFFR_X1 \core.keymem.key_mem[9][11]$_DFFE_PN0P_  (.D(_02651_),
    .RN(net95),
    .CK(clknet_leaf_59_clk),
    .Q(\core.keymem.key_mem[9][11] ),
    .QN(_19953_));
 DFFR_X1 \core.keymem.key_mem[9][120]$_DFFE_PN0P_  (.D(_02652_),
    .RN(net94),
    .CK(clknet_leaf_204_clk),
    .Q(\core.keymem.key_mem[9][120] ),
    .QN(_19952_));
 DFFR_X1 \core.keymem.key_mem[9][121]$_DFFE_PN0P_  (.D(_02653_),
    .RN(net92),
    .CK(clknet_leaf_265_clk),
    .Q(\core.keymem.key_mem[9][121] ),
    .QN(_19951_));
 DFFR_X1 \core.keymem.key_mem[9][122]$_DFFE_PN0P_  (.D(_02654_),
    .RN(net97),
    .CK(clknet_leaf_235_clk),
    .Q(\core.keymem.key_mem[9][122] ),
    .QN(_19950_));
 DFFR_X1 \core.keymem.key_mem[9][123]$_DFFE_PN0P_  (.D(_02655_),
    .RN(net93),
    .CK(clknet_leaf_195_clk),
    .Q(\core.keymem.key_mem[9][123] ),
    .QN(_19949_));
 DFFR_X1 \core.keymem.key_mem[9][124]$_DFFE_PN0P_  (.D(_02656_),
    .RN(net93),
    .CK(clknet_leaf_58_clk),
    .Q(\core.keymem.key_mem[9][124] ),
    .QN(_19948_));
 DFFR_X1 \core.keymem.key_mem[9][125]$_DFFE_PN0P_  (.D(_02657_),
    .RN(net97),
    .CK(clknet_leaf_231_clk),
    .Q(\core.keymem.key_mem[9][125] ),
    .QN(_19947_));
 DFFR_X1 \core.keymem.key_mem[9][126]$_DFFE_PN0P_  (.D(_02658_),
    .RN(net95),
    .CK(clknet_leaf_190_clk),
    .Q(\core.keymem.key_mem[9][126] ),
    .QN(_19946_));
 DFFR_X1 \core.keymem.key_mem[9][127]$_DFFE_PN0P_  (.D(_02659_),
    .RN(net97),
    .CK(clknet_leaf_235_clk),
    .Q(\core.keymem.key_mem[9][127] ),
    .QN(_19945_));
 DFFR_X1 \core.keymem.key_mem[9][12]$_DFFE_PN0P_  (.D(_02660_),
    .RN(net93),
    .CK(clknet_leaf_191_clk),
    .Q(\core.keymem.key_mem[9][12] ),
    .QN(_19944_));
 DFFR_X1 \core.keymem.key_mem[9][13]$_DFFE_PN0P_  (.D(_02661_),
    .RN(net87),
    .CK(clknet_leaf_32_clk),
    .Q(\core.keymem.key_mem[9][13] ),
    .QN(_19943_));
 DFFR_X1 \core.keymem.key_mem[9][14]$_DFFE_PN0P_  (.D(_02662_),
    .RN(net94),
    .CK(clknet_leaf_208_clk),
    .Q(\core.keymem.key_mem[9][14] ),
    .QN(_19942_));
 DFFR_X1 \core.keymem.key_mem[9][15]$_DFFE_PN0P_  (.D(_02663_),
    .RN(net98),
    .CK(clknet_leaf_229_clk),
    .Q(\core.keymem.key_mem[9][15] ),
    .QN(_19941_));
 DFFR_X1 \core.keymem.key_mem[9][16]$_DFFE_PN0P_  (.D(_02664_),
    .RN(net87),
    .CK(clknet_leaf_32_clk),
    .Q(\core.keymem.key_mem[9][16] ),
    .QN(_19940_));
 DFFR_X1 \core.keymem.key_mem[9][17]$_DFFE_PN0P_  (.D(_02665_),
    .RN(net95),
    .CK(clknet_leaf_185_clk),
    .Q(\core.keymem.key_mem[9][17] ),
    .QN(_19939_));
 DFFR_X1 \core.keymem.key_mem[9][18]$_DFFE_PN0P_  (.D(_02666_),
    .RN(net89),
    .CK(clknet_leaf_34_clk),
    .Q(\core.keymem.key_mem[9][18] ),
    .QN(_19938_));
 DFFR_X1 \core.keymem.key_mem[9][19]$_DFFE_PN0P_  (.D(_02667_),
    .RN(net85),
    .CK(clknet_leaf_50_clk),
    .Q(\core.keymem.key_mem[9][19] ),
    .QN(_19937_));
 DFFR_X1 \core.keymem.key_mem[9][1]$_DFFE_PN0P_  (.D(_02668_),
    .RN(net89),
    .CK(clknet_leaf_25_clk),
    .Q(\core.keymem.key_mem[9][1] ),
    .QN(_19936_));
 DFFR_X1 \core.keymem.key_mem[9][20]$_DFFE_PN0P_  (.D(_02669_),
    .RN(net82),
    .CK(clknet_leaf_23_clk),
    .Q(\core.keymem.key_mem[9][20] ),
    .QN(_19935_));
 DFFR_X1 \core.keymem.key_mem[9][21]$_DFFE_PN0P_  (.D(_02670_),
    .RN(net85),
    .CK(clknet_leaf_67_clk),
    .Q(\core.keymem.key_mem[9][21] ),
    .QN(_19934_));
 DFFR_X1 \core.keymem.key_mem[9][22]$_DFFE_PN0P_  (.D(_02671_),
    .RN(net96),
    .CK(clknet_leaf_221_clk),
    .Q(\core.keymem.key_mem[9][22] ),
    .QN(_19933_));
 DFFR_X1 \core.keymem.key_mem[9][23]$_DFFE_PN0P_  (.D(_02672_),
    .RN(net89),
    .CK(clknet_leaf_379_clk),
    .Q(\core.keymem.key_mem[9][23] ),
    .QN(_19932_));
 DFFR_X1 \core.keymem.key_mem[9][24]$_DFFE_PN0P_  (.D(_02673_),
    .RN(net85),
    .CK(clknet_leaf_49_clk),
    .Q(\core.keymem.key_mem[9][24] ),
    .QN(_19931_));
 DFFR_X1 \core.keymem.key_mem[9][25]$_DFFE_PN0P_  (.D(_02674_),
    .RN(net85),
    .CK(clknet_leaf_50_clk),
    .Q(\core.keymem.key_mem[9][25] ),
    .QN(_19930_));
 DFFR_X1 \core.keymem.key_mem[9][26]$_DFFE_PN0P_  (.D(_02675_),
    .RN(net89),
    .CK(clknet_leaf_21_clk),
    .Q(\core.keymem.key_mem[9][26] ),
    .QN(_19929_));
 DFFR_X1 \core.keymem.key_mem[9][27]$_DFFE_PN0P_  (.D(_02676_),
    .RN(net16),
    .CK(clknet_leaf_150_clk),
    .Q(\core.keymem.key_mem[9][27] ),
    .QN(_19928_));
 DFFR_X1 \core.keymem.key_mem[9][28]$_DFFE_PN0P_  (.D(_02677_),
    .RN(net16),
    .CK(clknet_leaf_125_clk),
    .Q(\core.keymem.key_mem[9][28] ),
    .QN(_19927_));
 DFFR_X1 \core.keymem.key_mem[9][29]$_DFFE_PN0P_  (.D(_02678_),
    .RN(net16),
    .CK(clknet_leaf_133_clk),
    .Q(\core.keymem.key_mem[9][29] ),
    .QN(_19926_));
 DFFR_X1 \core.keymem.key_mem[9][2]$_DFFE_PN0P_  (.D(_02679_),
    .RN(net89),
    .CK(clknet_leaf_64_clk),
    .Q(\core.keymem.key_mem[9][2] ),
    .QN(_19925_));
 DFFR_X1 \core.keymem.key_mem[9][30]$_DFFE_PN0P_  (.D(_02680_),
    .RN(net98),
    .CK(clknet_leaf_149_clk),
    .Q(\core.keymem.key_mem[9][30] ),
    .QN(_19924_));
 DFFR_X1 \core.keymem.key_mem[9][31]$_DFFE_PN0P_  (.D(_02681_),
    .RN(net16),
    .CK(clknet_leaf_138_clk),
    .Q(\core.keymem.key_mem[9][31] ),
    .QN(_19923_));
 DFFR_X1 \core.keymem.key_mem[9][32]$_DFFE_PN0P_  (.D(_02682_),
    .RN(net100),
    .CK(clknet_leaf_113_clk),
    .Q(\core.keymem.key_mem[9][32] ),
    .QN(_19922_));
 DFFR_X1 \core.keymem.key_mem[9][33]$_DFFE_PN0P_  (.D(_02683_),
    .RN(net99),
    .CK(clknet_leaf_112_clk),
    .Q(\core.keymem.key_mem[9][33] ),
    .QN(_19921_));
 DFFR_X1 \core.keymem.key_mem[9][34]$_DFFE_PN0P_  (.D(_02684_),
    .RN(net16),
    .CK(clknet_leaf_135_clk),
    .Q(\core.keymem.key_mem[9][34] ),
    .QN(_19920_));
 DFFR_X1 \core.keymem.key_mem[9][35]$_DFFE_PN0P_  (.D(_02685_),
    .RN(net99),
    .CK(clknet_leaf_112_clk),
    .Q(\core.keymem.key_mem[9][35] ),
    .QN(_19919_));
 DFFR_X1 \core.keymem.key_mem[9][36]$_DFFE_PN0P_  (.D(_02686_),
    .RN(net87),
    .CK(clknet_leaf_29_clk),
    .Q(\core.keymem.key_mem[9][36] ),
    .QN(_19918_));
 DFFR_X1 \core.keymem.key_mem[9][37]$_DFFE_PN0P_  (.D(_02687_),
    .RN(net89),
    .CK(clknet_leaf_85_clk),
    .Q(\core.keymem.key_mem[9][37] ),
    .QN(_19917_));
 DFFR_X1 \core.keymem.key_mem[9][38]$_DFFE_PN0P_  (.D(_02688_),
    .RN(net99),
    .CK(clknet_leaf_122_clk),
    .Q(\core.keymem.key_mem[9][38] ),
    .QN(_19916_));
 DFFR_X1 \core.keymem.key_mem[9][39]$_DFFE_PN0P_  (.D(_02689_),
    .RN(net99),
    .CK(clknet_leaf_86_clk),
    .Q(\core.keymem.key_mem[9][39] ),
    .QN(_19915_));
 DFFR_X1 \core.keymem.key_mem[9][3]$_DFFE_PN0P_  (.D(_02690_),
    .RN(net85),
    .CK(clknet_leaf_30_clk),
    .Q(\core.keymem.key_mem[9][3] ),
    .QN(_19914_));
 DFFR_X1 \core.keymem.key_mem[9][40]$_DFFE_PN0P_  (.D(_02691_),
    .RN(net85),
    .CK(clknet_leaf_89_clk),
    .Q(\core.keymem.key_mem[9][40] ),
    .QN(_19913_));
 DFFR_X1 \core.keymem.key_mem[9][41]$_DFFE_PN0P_  (.D(_02692_),
    .RN(net100),
    .CK(clknet_leaf_115_clk),
    .Q(\core.keymem.key_mem[9][41] ),
    .QN(_19912_));
 DFFR_X1 \core.keymem.key_mem[9][42]$_DFFE_PN0P_  (.D(_02693_),
    .RN(net100),
    .CK(clknet_leaf_110_clk),
    .Q(\core.keymem.key_mem[9][42] ),
    .QN(_19911_));
 DFFR_X1 \core.keymem.key_mem[9][43]$_DFFE_PN0P_  (.D(_02694_),
    .RN(net85),
    .CK(clknet_leaf_68_clk),
    .Q(\core.keymem.key_mem[9][43] ),
    .QN(_19910_));
 DFFR_X1 \core.keymem.key_mem[9][44]$_DFFE_PN0P_  (.D(_02695_),
    .RN(net89),
    .CK(clknet_leaf_114_clk),
    .Q(\core.keymem.key_mem[9][44] ),
    .QN(_19909_));
 DFFR_X1 \core.keymem.key_mem[9][45]$_DFFE_PN0P_  (.D(_02696_),
    .RN(net89),
    .CK(clknet_leaf_69_clk),
    .Q(\core.keymem.key_mem[9][45] ),
    .QN(_19908_));
 DFFR_X1 \core.keymem.key_mem[9][46]$_DFFE_PN0P_  (.D(_02697_),
    .RN(net99),
    .CK(clknet_leaf_80_clk),
    .Q(\core.keymem.key_mem[9][46] ),
    .QN(_19907_));
 DFFR_X2 \core.keymem.key_mem[9][47]$_DFFE_PN0P_  (.D(_02698_),
    .RN(net98),
    .CK(clknet_leaf_175_clk),
    .Q(\core.keymem.key_mem[9][47] ),
    .QN(_19906_));
 DFFR_X1 \core.keymem.key_mem[9][48]$_DFFE_PN0P_  (.D(_02699_),
    .RN(net95),
    .CK(clknet_leaf_120_clk),
    .Q(\core.keymem.key_mem[9][48] ),
    .QN(_19905_));
 DFFR_X1 \core.keymem.key_mem[9][49]$_DFFE_PN0P_  (.D(_02700_),
    .RN(net99),
    .CK(clknet_leaf_78_clk),
    .Q(\core.keymem.key_mem[9][49] ),
    .QN(_19904_));
 DFFR_X1 \core.keymem.key_mem[9][4]$_DFFE_PN0P_  (.D(_02701_),
    .RN(net100),
    .CK(clknet_leaf_104_clk),
    .Q(\core.keymem.key_mem[9][4] ),
    .QN(_19903_));
 DFFR_X1 \core.keymem.key_mem[9][50]$_DFFE_PN0P_  (.D(_02702_),
    .RN(net98),
    .CK(clknet_leaf_139_clk),
    .Q(\core.keymem.key_mem[9][50] ),
    .QN(_19902_));
 DFFR_X1 \core.keymem.key_mem[9][51]$_DFFE_PN0P_  (.D(_02703_),
    .RN(net99),
    .CK(clknet_leaf_129_clk),
    .Q(\core.keymem.key_mem[9][51] ),
    .QN(_19901_));
 DFFR_X1 \core.keymem.key_mem[9][52]$_DFFE_PN0P_  (.D(_02704_),
    .RN(net99),
    .CK(clknet_leaf_80_clk),
    .Q(\core.keymem.key_mem[9][52] ),
    .QN(_19900_));
 DFFR_X2 \core.keymem.key_mem[9][53]$_DFFE_PN0P_  (.D(_02705_),
    .RN(net98),
    .CK(clknet_leaf_176_clk),
    .Q(\core.keymem.key_mem[9][53] ),
    .QN(_19899_));
 DFFR_X1 \core.keymem.key_mem[9][54]$_DFFE_PN0P_  (.D(_02706_),
    .RN(net98),
    .CK(clknet_leaf_141_clk),
    .Q(\core.keymem.key_mem[9][54] ),
    .QN(_19898_));
 DFFR_X1 \core.keymem.key_mem[9][55]$_DFFE_PN0P_  (.D(_02707_),
    .RN(net16),
    .CK(clknet_leaf_135_clk),
    .Q(\core.keymem.key_mem[9][55] ),
    .QN(_19897_));
 DFFR_X1 \core.keymem.key_mem[9][56]$_DFFE_PN0P_  (.D(_02708_),
    .RN(net98),
    .CK(clknet_leaf_148_clk),
    .Q(\core.keymem.key_mem[9][56] ),
    .QN(_19896_));
 DFFR_X1 \core.keymem.key_mem[9][57]$_DFFE_PN0P_  (.D(_02709_),
    .RN(net100),
    .CK(clknet_leaf_110_clk),
    .Q(\core.keymem.key_mem[9][57] ),
    .QN(_19895_));
 DFFR_X1 \core.keymem.key_mem[9][58]$_DFFE_PN0P_  (.D(_02710_),
    .RN(net100),
    .CK(clknet_leaf_103_clk),
    .Q(\core.keymem.key_mem[9][58] ),
    .QN(_19894_));
 DFFR_X1 \core.keymem.key_mem[9][59]$_DFFE_PN0P_  (.D(_02711_),
    .RN(net82),
    .CK(clknet_leaf_23_clk),
    .Q(\core.keymem.key_mem[9][59] ),
    .QN(_19893_));
 DFFR_X1 \core.keymem.key_mem[9][5]$_DFFE_PN0P_  (.D(_02712_),
    .RN(net100),
    .CK(clknet_leaf_18_clk),
    .Q(\core.keymem.key_mem[9][5] ),
    .QN(_19892_));
 DFFR_X1 \core.keymem.key_mem[9][60]$_DFFE_PN0P_  (.D(_02713_),
    .RN(net82),
    .CK(clknet_leaf_24_clk),
    .Q(\core.keymem.key_mem[9][60] ),
    .QN(_19891_));
 DFFR_X1 \core.keymem.key_mem[9][61]$_DFFE_PN0P_  (.D(_02714_),
    .RN(net88),
    .CK(clknet_leaf_93_clk),
    .Q(\core.keymem.key_mem[9][61] ),
    .QN(_19890_));
 DFFR_X1 \core.keymem.key_mem[9][62]$_DFFE_PN0P_  (.D(_02715_),
    .RN(net100),
    .CK(clknet_leaf_99_clk),
    .Q(\core.keymem.key_mem[9][62] ),
    .QN(_19889_));
 DFFR_X1 \core.keymem.key_mem[9][63]$_DFFE_PN0P_  (.D(_02716_),
    .RN(net100),
    .CK(clknet_leaf_21_clk),
    .Q(\core.keymem.key_mem[9][63] ),
    .QN(_19888_));
 DFFR_X1 \core.keymem.key_mem[9][64]$_DFFE_PN0P_  (.D(_02717_),
    .RN(net82),
    .CK(clknet_leaf_14_clk),
    .Q(\core.keymem.key_mem[9][64] ),
    .QN(_19887_));
 DFFR_X1 \core.keymem.key_mem[9][65]$_DFFE_PN0P_  (.D(_02718_),
    .RN(net99),
    .CK(clknet_leaf_120_clk),
    .Q(\core.keymem.key_mem[9][65] ),
    .QN(_19886_));
 DFFR_X1 \core.keymem.key_mem[9][66]$_DFFE_PN0P_  (.D(_02719_),
    .RN(net100),
    .CK(clknet_leaf_16_clk),
    .Q(\core.keymem.key_mem[9][66] ),
    .QN(_19885_));
 DFFR_X1 \core.keymem.key_mem[9][67]$_DFFE_PN0P_  (.D(_02720_),
    .RN(net99),
    .CK(clknet_leaf_79_clk),
    .Q(\core.keymem.key_mem[9][67] ),
    .QN(_19884_));
 DFFR_X1 \core.keymem.key_mem[9][68]$_DFFE_PN0P_  (.D(_02721_),
    .RN(net95),
    .CK(clknet_leaf_118_clk),
    .Q(\core.keymem.key_mem[9][68] ),
    .QN(_19883_));
 DFFR_X1 \core.keymem.key_mem[9][69]$_DFFE_PN0P_  (.D(_02722_),
    .RN(net98),
    .CK(clknet_leaf_178_clk),
    .Q(\core.keymem.key_mem[9][69] ),
    .QN(_19882_));
 DFFR_X1 \core.keymem.key_mem[9][6]$_DFFE_PN0P_  (.D(_02723_),
    .RN(net100),
    .CK(clknet_leaf_95_clk),
    .Q(\core.keymem.key_mem[9][6] ),
    .QN(_19881_));
 DFFR_X1 \core.keymem.key_mem[9][70]$_DFFE_PN0P_  (.D(_02724_),
    .RN(net100),
    .CK(clknet_leaf_100_clk),
    .Q(\core.keymem.key_mem[9][70] ),
    .QN(_19880_));
 DFFR_X1 \core.keymem.key_mem[9][71]$_DFFE_PN0P_  (.D(_02725_),
    .RN(net99),
    .CK(clknet_leaf_74_clk),
    .Q(\core.keymem.key_mem[9][71] ),
    .QN(_19879_));
 DFFR_X1 \core.keymem.key_mem[9][72]$_DFFE_PN0P_  (.D(_02726_),
    .RN(net95),
    .CK(clknet_leaf_75_clk),
    .Q(\core.keymem.key_mem[9][72] ),
    .QN(_19878_));
 DFFR_X1 \core.keymem.key_mem[9][73]$_DFFE_PN0P_  (.D(_02727_),
    .RN(net97),
    .CK(clknet_leaf_147_clk),
    .Q(\core.keymem.key_mem[9][73] ),
    .QN(_19877_));
 DFFR_X1 \core.keymem.key_mem[9][74]$_DFFE_PN0P_  (.D(_02728_),
    .RN(net97),
    .CK(clknet_leaf_163_clk),
    .Q(\core.keymem.key_mem[9][74] ),
    .QN(_19876_));
 DFFR_X1 \core.keymem.key_mem[9][75]$_DFFE_PN0P_  (.D(_02729_),
    .RN(net97),
    .CK(clknet_leaf_154_clk),
    .Q(\core.keymem.key_mem[9][75] ),
    .QN(_19875_));
 DFFR_X1 \core.keymem.key_mem[9][76]$_DFFE_PN0P_  (.D(_02730_),
    .RN(net93),
    .CK(clknet_leaf_376_clk),
    .Q(\core.keymem.key_mem[9][76] ),
    .QN(_19874_));
 DFFR_X1 \core.keymem.key_mem[9][77]$_DFFE_PN0P_  (.D(_02731_),
    .RN(net97),
    .CK(clknet_leaf_161_clk),
    .Q(\core.keymem.key_mem[9][77] ),
    .QN(_19873_));
 DFFR_X1 \core.keymem.key_mem[9][78]$_DFFE_PN0P_  (.D(_02732_),
    .RN(net98),
    .CK(clknet_leaf_170_clk),
    .Q(\core.keymem.key_mem[9][78] ),
    .QN(_19872_));
 DFFR_X1 \core.keymem.key_mem[9][79]$_DFFE_PN0P_  (.D(_02733_),
    .RN(net98),
    .CK(clknet_leaf_229_clk),
    .Q(\core.keymem.key_mem[9][79] ),
    .QN(_19871_));
 DFFR_X1 \core.keymem.key_mem[9][7]$_DFFE_PN0P_  (.D(_02734_),
    .RN(net98),
    .CK(clknet_leaf_173_clk),
    .Q(\core.keymem.key_mem[9][7] ),
    .QN(_19870_));
 DFFR_X1 \core.keymem.key_mem[9][80]$_DFFE_PN0P_  (.D(_02735_),
    .RN(net97),
    .CK(clknet_leaf_160_clk),
    .Q(\core.keymem.key_mem[9][80] ),
    .QN(_19869_));
 DFFR_X1 \core.keymem.key_mem[9][81]$_DFFE_PN0P_  (.D(_02736_),
    .RN(net96),
    .CK(clknet_leaf_164_clk),
    .Q(\core.keymem.key_mem[9][81] ),
    .QN(_19868_));
 DFFR_X1 \core.keymem.key_mem[9][82]$_DFFE_PN0P_  (.D(_02737_),
    .RN(net98),
    .CK(clknet_leaf_180_clk),
    .Q(\core.keymem.key_mem[9][82] ),
    .QN(_19867_));
 DFFR_X1 \core.keymem.key_mem[9][83]$_DFFE_PN0P_  (.D(_02738_),
    .RN(net95),
    .CK(clknet_leaf_182_clk),
    .Q(\core.keymem.key_mem[9][83] ),
    .QN(_19866_));
 DFFR_X1 \core.keymem.key_mem[9][84]$_DFFE_PN0P_  (.D(_02739_),
    .RN(net95),
    .CK(clknet_leaf_182_clk),
    .Q(\core.keymem.key_mem[9][84] ),
    .QN(_19865_));
 DFFR_X1 \core.keymem.key_mem[9][85]$_DFFE_PN0P_  (.D(_02740_),
    .RN(net97),
    .CK(clknet_leaf_237_clk),
    .Q(\core.keymem.key_mem[9][85] ),
    .QN(_19864_));
 DFFR_X1 \core.keymem.key_mem[9][86]$_DFFE_PN0P_  (.D(_02741_),
    .RN(net95),
    .CK(clknet_leaf_209_clk),
    .Q(\core.keymem.key_mem[9][86] ),
    .QN(_19863_));
 DFFR_X1 \core.keymem.key_mem[9][87]$_DFFE_PN0P_  (.D(_02742_),
    .RN(net89),
    .CK(clknet_leaf_378_clk),
    .Q(\core.keymem.key_mem[9][87] ),
    .QN(_19862_));
 DFFR_X1 \core.keymem.key_mem[9][88]$_DFFE_PN0P_  (.D(_02743_),
    .RN(net93),
    .CK(clknet_leaf_280_clk),
    .Q(\core.keymem.key_mem[9][88] ),
    .QN(_19861_));
 DFFR_X1 \core.keymem.key_mem[9][89]$_DFFE_PN0P_  (.D(_02744_),
    .RN(net93),
    .CK(clknet_leaf_200_clk),
    .Q(\core.keymem.key_mem[9][89] ),
    .QN(_19860_));
 DFFR_X1 \core.keymem.key_mem[9][8]$_DFFE_PN0P_  (.D(_02745_),
    .RN(net89),
    .CK(clknet_leaf_378_clk),
    .Q(\core.keymem.key_mem[9][8] ),
    .QN(_19859_));
 DFFR_X1 \core.keymem.key_mem[9][90]$_DFFE_PN0P_  (.D(_02746_),
    .RN(net97),
    .CK(clknet_leaf_163_clk),
    .Q(\core.keymem.key_mem[9][90] ),
    .QN(_19858_));
 DFFR_X1 \core.keymem.key_mem[9][91]$_DFFE_PN0P_  (.D(_02747_),
    .RN(net95),
    .CK(clknet_leaf_182_clk),
    .Q(\core.keymem.key_mem[9][91] ),
    .QN(_19857_));
 DFFR_X1 \core.keymem.key_mem[9][92]$_DFFE_PN0P_  (.D(_02748_),
    .RN(net95),
    .CK(clknet_leaf_63_clk),
    .Q(\core.keymem.key_mem[9][92] ),
    .QN(_19856_));
 DFFR_X1 \core.keymem.key_mem[9][93]$_DFFE_PN0P_  (.D(_02749_),
    .RN(net98),
    .CK(clknet_leaf_188_clk),
    .Q(\core.keymem.key_mem[9][93] ),
    .QN(_19855_));
 DFFR_X1 \core.keymem.key_mem[9][94]$_DFFE_PN0P_  (.D(_02750_),
    .RN(net94),
    .CK(clknet_leaf_214_clk),
    .Q(\core.keymem.key_mem[9][94] ),
    .QN(_19854_));
 DFFR_X1 \core.keymem.key_mem[9][95]$_DFFE_PN0P_  (.D(_02751_),
    .RN(net96),
    .CK(clknet_leaf_234_clk),
    .Q(\core.keymem.key_mem[9][95] ),
    .QN(_19853_));
 DFFR_X1 \core.keymem.key_mem[9][96]$_DFFE_PN0P_  (.D(_02752_),
    .RN(net92),
    .CK(clknet_leaf_204_clk),
    .Q(\core.keymem.key_mem[9][96] ),
    .QN(_19852_));
 DFFR_X1 \core.keymem.key_mem[9][97]$_DFFE_PN0P_  (.D(_02753_),
    .RN(net95),
    .CK(clknet_leaf_72_clk),
    .Q(\core.keymem.key_mem[9][97] ),
    .QN(_19851_));
 DFFR_X1 \core.keymem.key_mem[9][98]$_DFFE_PN0P_  (.D(_02754_),
    .RN(net95),
    .CK(clknet_leaf_63_clk),
    .Q(\core.keymem.key_mem[9][98] ),
    .QN(_19850_));
 DFFR_X1 \core.keymem.key_mem[9][99]$_DFFE_PN0P_  (.D(_02755_),
    .RN(net92),
    .CK(clknet_leaf_197_clk),
    .Q(\core.keymem.key_mem[9][99] ),
    .QN(_19849_));
 DFFR_X1 \core.keymem.key_mem[9][9]$_DFFE_PN0P_  (.D(_02756_),
    .RN(net92),
    .CK(clknet_leaf_202_clk),
    .Q(\core.keymem.key_mem[9][9] ),
    .QN(_21959_));
 DFFS_X1 \core.keymem.key_mem_ctrl_reg[0]$_DFF_PN1_  (.D(_00013_),
    .SN(net88),
    .CK(clknet_leaf_42_clk),
    .Q(\core.keymem.key_mem_ctrl_reg[0] ),
    .QN(_00320_));
 DFFR_X2 \core.keymem.key_mem_ctrl_reg[1]$_DFF_PN0_  (.D(_00014_),
    .RN(net88),
    .CK(clknet_leaf_41_clk),
    .Q(\core.keymem.key_mem_ctrl_reg[1] ),
    .QN(_00318_));
 DFFR_X1 \core.keymem.key_mem_ctrl_reg[2]$_DFF_PN0_  (.D(_00004_),
    .RN(net88),
    .CK(clknet_leaf_42_clk),
    .Q(\core.keymem.key_mem_ctrl_reg[2] ),
    .QN(_00326_));
 DFFR_X1 \core.keymem.key_mem_ctrl_reg[3]$_DFF_PN0_  (.D(_00005_),
    .RN(net88),
    .CK(clknet_leaf_42_clk),
    .Q(\core.keymem.key_mem_ctrl_reg[3] ),
    .QN(_19848_));
 DFFR_X1 \core.keymem.prev_key0_reg[0]$_DFFE_PN0P_  (.D(_02757_),
    .RN(net88),
    .CK(clknet_leaf_399_clk),
    .Q(\core.keymem.prev_key0_reg[0] ),
    .QN(_19847_));
 DFFR_X2 \core.keymem.prev_key0_reg[100]$_DFFE_PN0P_  (.D(_02758_),
    .RN(net82),
    .CK(clknet_leaf_8_clk),
    .Q(\core.keymem.prev_key0_reg[100] ),
    .QN(_19846_));
 DFFR_X1 \core.keymem.prev_key0_reg[101]$_DFFE_PN0P_  (.D(_02759_),
    .RN(net82),
    .CK(clknet_leaf_5_clk),
    .Q(\core.keymem.prev_key0_reg[101] ),
    .QN(_19845_));
 DFFR_X1 \core.keymem.prev_key0_reg[102]$_DFFE_PN0P_  (.D(_02760_),
    .RN(net82),
    .CK(clknet_leaf_423_clk),
    .Q(\core.keymem.prev_key0_reg[102] ),
    .QN(_19844_));
 DFFR_X1 \core.keymem.prev_key0_reg[103]$_DFFE_PN0P_  (.D(_02761_),
    .RN(net82),
    .CK(clknet_leaf_423_clk),
    .Q(\core.keymem.prev_key0_reg[103] ),
    .QN(_19843_));
 DFFR_X1 \core.keymem.prev_key0_reg[104]$_DFFE_PN0P_  (.D(_02762_),
    .RN(net86),
    .CK(clknet_leaf_407_clk),
    .Q(\core.keymem.prev_key0_reg[104] ),
    .QN(_19842_));
 DFFR_X2 \core.keymem.prev_key0_reg[105]$_DFFE_PN0P_  (.D(_02763_),
    .RN(net84),
    .CK(clknet_leaf_352_clk),
    .Q(\core.keymem.prev_key0_reg[105] ),
    .QN(_19841_));
 DFFR_X1 \core.keymem.prev_key0_reg[106]$_DFFE_PN0P_  (.D(_02764_),
    .RN(net86),
    .CK(clknet_leaf_406_clk),
    .Q(\core.keymem.prev_key0_reg[106] ),
    .QN(_19840_));
 DFFR_X1 \core.keymem.prev_key0_reg[107]$_DFFE_PN0P_  (.D(_02765_),
    .RN(net86),
    .CK(clknet_leaf_388_clk),
    .Q(\core.keymem.prev_key0_reg[107] ),
    .QN(_19839_));
 DFFR_X1 \core.keymem.prev_key0_reg[108]$_DFFE_PN0P_  (.D(_02766_),
    .RN(net86),
    .CK(clknet_leaf_345_clk),
    .Q(\core.keymem.prev_key0_reg[108] ),
    .QN(_19838_));
 DFFR_X1 \core.keymem.prev_key0_reg[109]$_DFFE_PN0P_  (.D(_02767_),
    .RN(net88),
    .CK(clknet_leaf_399_clk),
    .Q(\core.keymem.prev_key0_reg[109] ),
    .QN(_19837_));
 DFFR_X1 \core.keymem.prev_key0_reg[10]$_DFFE_PN0P_  (.D(_02768_),
    .RN(net86),
    .CK(clknet_leaf_407_clk),
    .Q(\core.keymem.prev_key0_reg[10] ),
    .QN(_19836_));
 DFFR_X1 \core.keymem.prev_key0_reg[110]$_DFFE_PN0P_  (.D(_02769_),
    .RN(net86),
    .CK(clknet_leaf_348_clk),
    .Q(\core.keymem.prev_key0_reg[110] ),
    .QN(_19835_));
 DFFR_X1 \core.keymem.prev_key0_reg[111]$_DFFE_PN0P_  (.D(_02770_),
    .RN(net86),
    .CK(clknet_leaf_345_clk),
    .Q(\core.keymem.prev_key0_reg[111] ),
    .QN(_19834_));
 DFFR_X2 \core.keymem.prev_key0_reg[112]$_DFFE_PN0P_  (.D(_02771_),
    .RN(net84),
    .CK(clknet_leaf_353_clk),
    .Q(\core.keymem.prev_key0_reg[112] ),
    .QN(_19833_));
 DFFR_X2 \core.keymem.prev_key0_reg[113]$_DFFE_PN0P_  (.D(_02772_),
    .RN(net84),
    .CK(clknet_leaf_353_clk),
    .Q(\core.keymem.prev_key0_reg[113] ),
    .QN(_19832_));
 DFFR_X1 \core.keymem.prev_key0_reg[114]$_DFFE_PN0P_  (.D(_02773_),
    .RN(net86),
    .CK(clknet_leaf_408_clk),
    .Q(\core.keymem.prev_key0_reg[114] ),
    .QN(_19831_));
 DFFR_X1 \core.keymem.prev_key0_reg[115]$_DFFE_PN0P_  (.D(_02774_),
    .RN(net86),
    .CK(clknet_leaf_345_clk),
    .Q(\core.keymem.prev_key0_reg[115] ),
    .QN(_19830_));
 DFFR_X1 \core.keymem.prev_key0_reg[116]$_DFFE_PN0P_  (.D(_02775_),
    .RN(net86),
    .CK(clknet_leaf_345_clk),
    .Q(\core.keymem.prev_key0_reg[116] ),
    .QN(_19829_));
 DFFR_X2 \core.keymem.prev_key0_reg[117]$_DFFE_PN0P_  (.D(_02776_),
    .RN(net86),
    .CK(clknet_leaf_348_clk),
    .Q(\core.keymem.prev_key0_reg[117] ),
    .QN(_19828_));
 DFFR_X1 \core.keymem.prev_key0_reg[118]$_DFFE_PN0P_  (.D(_02777_),
    .RN(net86),
    .CK(clknet_leaf_346_clk),
    .Q(\core.keymem.prev_key0_reg[118] ),
    .QN(_19827_));
 DFFR_X1 \core.keymem.prev_key0_reg[119]$_DFFE_PN0P_  (.D(_02778_),
    .RN(net86),
    .CK(clknet_leaf_345_clk),
    .Q(\core.keymem.prev_key0_reg[119] ),
    .QN(_19826_));
 DFFR_X1 \core.keymem.prev_key0_reg[11]$_DFFE_PN0P_  (.D(_02779_),
    .RN(net86),
    .CK(clknet_leaf_398_clk),
    .Q(\core.keymem.prev_key0_reg[11] ),
    .QN(_19825_));
 DFFR_X1 \core.keymem.prev_key0_reg[120]$_DFFE_PN0P_  (.D(_02780_),
    .RN(net86),
    .CK(clknet_leaf_406_clk),
    .Q(\core.keymem.prev_key0_reg[120] ),
    .QN(_19824_));
 DFFR_X1 \core.keymem.prev_key0_reg[121]$_DFFE_PN0P_  (.D(_02781_),
    .RN(net86),
    .CK(clknet_leaf_410_clk),
    .Q(\core.keymem.prev_key0_reg[121] ),
    .QN(_19823_));
 DFFR_X1 \core.keymem.prev_key0_reg[122]$_DFFE_PN0P_  (.D(_02782_),
    .RN(net87),
    .CK(clknet_leaf_409_clk),
    .Q(\core.keymem.prev_key0_reg[122] ),
    .QN(_19822_));
 DFFR_X1 \core.keymem.prev_key0_reg[123]$_DFFE_PN0P_  (.D(_02783_),
    .RN(net82),
    .CK(clknet_leaf_422_clk),
    .Q(\core.keymem.prev_key0_reg[123] ),
    .QN(_19821_));
 DFFR_X1 \core.keymem.prev_key0_reg[124]$_DFFE_PN0P_  (.D(_02784_),
    .RN(net82),
    .CK(clknet_leaf_423_clk),
    .Q(\core.keymem.prev_key0_reg[124] ),
    .QN(_19820_));
 DFFR_X1 \core.keymem.prev_key0_reg[125]$_DFFE_PN0P_  (.D(_02785_),
    .RN(net87),
    .CK(clknet_leaf_416_clk),
    .Q(\core.keymem.prev_key0_reg[125] ),
    .QN(_19819_));
 DFFR_X1 \core.keymem.prev_key0_reg[126]$_DFFE_PN0P_  (.D(_02786_),
    .RN(net82),
    .CK(clknet_leaf_411_clk),
    .Q(\core.keymem.prev_key0_reg[126] ),
    .QN(_19818_));
 DFFR_X1 \core.keymem.prev_key0_reg[127]$_DFFE_PN0P_  (.D(_02787_),
    .RN(net82),
    .CK(clknet_leaf_421_clk),
    .Q(\core.keymem.prev_key0_reg[127] ),
    .QN(_19817_));
 DFFR_X1 \core.keymem.prev_key0_reg[12]$_DFFE_PN0P_  (.D(_02788_),
    .RN(net86),
    .CK(clknet_leaf_404_clk),
    .Q(\core.keymem.prev_key0_reg[12] ),
    .QN(_19816_));
 DFFR_X1 \core.keymem.prev_key0_reg[13]$_DFFE_PN0P_  (.D(_02789_),
    .RN(net86),
    .CK(clknet_leaf_392_clk),
    .Q(\core.keymem.prev_key0_reg[13] ),
    .QN(_19815_));
 DFFR_X1 \core.keymem.prev_key0_reg[14]$_DFFE_PN0P_  (.D(_02790_),
    .RN(net86),
    .CK(clknet_leaf_347_clk),
    .Q(\core.keymem.prev_key0_reg[14] ),
    .QN(_19814_));
 DFFR_X1 \core.keymem.prev_key0_reg[15]$_DFFE_PN0P_  (.D(_02791_),
    .RN(net86),
    .CK(clknet_leaf_346_clk),
    .Q(\core.keymem.prev_key0_reg[15] ),
    .QN(_19813_));
 DFFR_X1 \core.keymem.prev_key0_reg[16]$_DFFE_PN0P_  (.D(_02792_),
    .RN(net84),
    .CK(clknet_leaf_351_clk),
    .Q(\core.keymem.prev_key0_reg[16] ),
    .QN(_19812_));
 DFFR_X1 \core.keymem.prev_key0_reg[17]$_DFFE_PN0P_  (.D(_02793_),
    .RN(net84),
    .CK(clknet_leaf_367_clk),
    .Q(\core.keymem.prev_key0_reg[17] ),
    .QN(_19811_));
 DFFR_X1 \core.keymem.prev_key0_reg[18]$_DFFE_PN0P_  (.D(_02794_),
    .RN(net86),
    .CK(clknet_leaf_409_clk),
    .Q(\core.keymem.prev_key0_reg[18] ),
    .QN(_19810_));
 DFFR_X1 \core.keymem.prev_key0_reg[19]$_DFFE_PN0P_  (.D(_02795_),
    .RN(net86),
    .CK(clknet_leaf_395_clk),
    .Q(\core.keymem.prev_key0_reg[19] ),
    .QN(_19809_));
 DFFR_X1 \core.keymem.prev_key0_reg[1]$_DFFE_PN0P_  (.D(_02796_),
    .RN(net87),
    .CK(clknet_leaf_394_clk),
    .Q(\core.keymem.prev_key0_reg[1] ),
    .QN(_19808_));
 DFFR_X1 \core.keymem.prev_key0_reg[20]$_DFFE_PN0P_  (.D(_02797_),
    .RN(net86),
    .CK(clknet_leaf_405_clk),
    .Q(\core.keymem.prev_key0_reg[20] ),
    .QN(_19807_));
 DFFR_X1 \core.keymem.prev_key0_reg[21]$_DFFE_PN0P_  (.D(_02798_),
    .RN(net86),
    .CK(clknet_leaf_404_clk),
    .Q(\core.keymem.prev_key0_reg[21] ),
    .QN(_19806_));
 DFFR_X2 \core.keymem.prev_key0_reg[22]$_DFFE_PN0P_  (.D(_02799_),
    .RN(net86),
    .CK(clknet_leaf_405_clk),
    .Q(\core.keymem.prev_key0_reg[22] ),
    .QN(_19805_));
 DFFR_X1 \core.keymem.prev_key0_reg[23]$_DFFE_PN0P_  (.D(_02800_),
    .RN(net86),
    .CK(clknet_leaf_405_clk),
    .Q(\core.keymem.prev_key0_reg[23] ),
    .QN(_19804_));
 DFFR_X1 \core.keymem.prev_key0_reg[24]$_DFFE_PN0P_  (.D(_02801_),
    .RN(net86),
    .CK(clknet_leaf_414_clk),
    .Q(\core.keymem.prev_key0_reg[24] ),
    .QN(_19803_));
 DFFR_X1 \core.keymem.prev_key0_reg[25]$_DFFE_PN0P_  (.D(_02802_),
    .RN(net86),
    .CK(clknet_leaf_409_clk),
    .Q(\core.keymem.prev_key0_reg[25] ),
    .QN(_19802_));
 DFFR_X1 \core.keymem.prev_key0_reg[26]$_DFFE_PN0P_  (.D(_02803_),
    .RN(net87),
    .CK(clknet_leaf_411_clk),
    .Q(\core.keymem.prev_key0_reg[26] ),
    .QN(_19801_));
 DFFR_X1 \core.keymem.prev_key0_reg[27]$_DFFE_PN0P_  (.D(_02804_),
    .RN(net87),
    .CK(clknet_leaf_411_clk),
    .Q(\core.keymem.prev_key0_reg[27] ),
    .QN(_19800_));
 DFFR_X1 \core.keymem.prev_key0_reg[28]$_DFFE_PN0P_  (.D(_02805_),
    .RN(net82),
    .CK(clknet_leaf_38_clk),
    .Q(\core.keymem.prev_key0_reg[28] ),
    .QN(_19799_));
 DFFR_X1 \core.keymem.prev_key0_reg[29]$_DFFE_PN0P_  (.D(_02806_),
    .RN(net82),
    .CK(clknet_leaf_421_clk),
    .Q(\core.keymem.prev_key0_reg[29] ),
    .QN(_19798_));
 DFFR_X1 \core.keymem.prev_key0_reg[2]$_DFFE_PN0P_  (.D(_02807_),
    .RN(net87),
    .CK(clknet_leaf_413_clk),
    .Q(\core.keymem.prev_key0_reg[2] ),
    .QN(_19797_));
 DFFR_X1 \core.keymem.prev_key0_reg[30]$_DFFE_PN0P_  (.D(_02808_),
    .RN(net87),
    .CK(clknet_leaf_421_clk),
    .Q(\core.keymem.prev_key0_reg[30] ),
    .QN(_19796_));
 DFFR_X1 \core.keymem.prev_key0_reg[31]$_DFFE_PN0P_  (.D(_02809_),
    .RN(net82),
    .CK(clknet_leaf_421_clk),
    .Q(\core.keymem.prev_key0_reg[31] ),
    .QN(_19795_));
 DFFR_X1 \core.keymem.prev_key0_reg[32]$_DFFE_PN0P_  (.D(_02810_),
    .RN(net88),
    .CK(clknet_leaf_386_clk),
    .Q(\core.keymem.prev_key0_reg[32] ),
    .QN(_19794_));
 DFFR_X1 \core.keymem.prev_key0_reg[33]$_DFFE_PN0P_  (.D(_02811_),
    .RN(net87),
    .CK(clknet_leaf_40_clk),
    .Q(\core.keymem.prev_key0_reg[33] ),
    .QN(_19793_));
 DFFR_X1 \core.keymem.prev_key0_reg[34]$_DFFE_PN0P_  (.D(_02812_),
    .RN(net82),
    .CK(clknet_leaf_424_clk),
    .Q(\core.keymem.prev_key0_reg[34] ),
    .QN(_19792_));
 DFFR_X1 \core.keymem.prev_key0_reg[35]$_DFFE_PN0P_  (.D(_02813_),
    .RN(net82),
    .CK(clknet_leaf_424_clk),
    .Q(\core.keymem.prev_key0_reg[35] ),
    .QN(_19791_));
 DFFR_X1 \core.keymem.prev_key0_reg[36]$_DFFE_PN0P_  (.D(_02814_),
    .RN(net82),
    .CK(clknet_leaf_8_clk),
    .Q(\core.keymem.prev_key0_reg[36] ),
    .QN(_19790_));
 DFFR_X1 \core.keymem.prev_key0_reg[37]$_DFFE_PN0P_  (.D(_02815_),
    .RN(net82),
    .CK(clknet_leaf_5_clk),
    .Q(\core.keymem.prev_key0_reg[37] ),
    .QN(_19789_));
 DFFR_X1 \core.keymem.prev_key0_reg[38]$_DFFE_PN0P_  (.D(_02816_),
    .RN(net82),
    .CK(clknet_leaf_423_clk),
    .Q(\core.keymem.prev_key0_reg[38] ),
    .QN(_19788_));
 DFFR_X1 \core.keymem.prev_key0_reg[39]$_DFFE_PN0P_  (.D(_02817_),
    .RN(net82),
    .CK(clknet_leaf_422_clk),
    .Q(\core.keymem.prev_key0_reg[39] ),
    .QN(_19787_));
 DFFR_X1 \core.keymem.prev_key0_reg[3]$_DFFE_PN0P_  (.D(_02818_),
    .RN(net82),
    .CK(clknet_leaf_420_clk),
    .Q(\core.keymem.prev_key0_reg[3] ),
    .QN(_19786_));
 DFFR_X1 \core.keymem.prev_key0_reg[40]$_DFFE_PN0P_  (.D(_02819_),
    .RN(net86),
    .CK(clknet_leaf_408_clk),
    .Q(\core.keymem.prev_key0_reg[40] ),
    .QN(_19785_));
 DFFR_X1 \core.keymem.prev_key0_reg[41]$_DFFE_PN0P_  (.D(_02820_),
    .RN(net86),
    .CK(clknet_leaf_393_clk),
    .Q(\core.keymem.prev_key0_reg[41] ),
    .QN(_19784_));
 DFFR_X1 \core.keymem.prev_key0_reg[42]$_DFFE_PN0P_  (.D(_02821_),
    .RN(net86),
    .CK(clknet_leaf_407_clk),
    .Q(\core.keymem.prev_key0_reg[42] ),
    .QN(_19783_));
 DFFR_X1 \core.keymem.prev_key0_reg[43]$_DFFE_PN0P_  (.D(_02822_),
    .RN(net88),
    .CK(clknet_leaf_388_clk),
    .Q(\core.keymem.prev_key0_reg[43] ),
    .QN(_19782_));
 DFFR_X1 \core.keymem.prev_key0_reg[44]$_DFFE_PN0P_  (.D(_02823_),
    .RN(net86),
    .CK(clknet_leaf_406_clk),
    .Q(\core.keymem.prev_key0_reg[44] ),
    .QN(_19781_));
 DFFR_X1 \core.keymem.prev_key0_reg[45]$_DFFE_PN0P_  (.D(_02824_),
    .RN(net86),
    .CK(clknet_leaf_392_clk),
    .Q(\core.keymem.prev_key0_reg[45] ),
    .QN(_19780_));
 DFFR_X1 \core.keymem.prev_key0_reg[46]$_DFFE_PN0P_  (.D(_02825_),
    .RN(net86),
    .CK(clknet_leaf_404_clk),
    .Q(\core.keymem.prev_key0_reg[46] ),
    .QN(_19779_));
 DFFR_X2 \core.keymem.prev_key0_reg[47]$_DFFE_PN0P_  (.D(_02826_),
    .RN(net84),
    .CK(clknet_leaf_386_clk),
    .Q(\core.keymem.prev_key0_reg[47] ),
    .QN(_19778_));
 DFFR_X1 \core.keymem.prev_key0_reg[48]$_DFFE_PN0P_  (.D(_02827_),
    .RN(net84),
    .CK(clknet_leaf_351_clk),
    .Q(\core.keymem.prev_key0_reg[48] ),
    .QN(_19777_));
 DFFR_X2 \core.keymem.prev_key0_reg[49]$_DFFE_PN0P_  (.D(_02828_),
    .RN(net88),
    .CK(clknet_leaf_387_clk),
    .Q(\core.keymem.prev_key0_reg[49] ),
    .QN(_19776_));
 DFFR_X1 \core.keymem.prev_key0_reg[4]$_DFFE_PN0P_  (.D(_02829_),
    .RN(net82),
    .CK(clknet_leaf_7_clk),
    .Q(\core.keymem.prev_key0_reg[4] ),
    .QN(_19775_));
 DFFR_X1 \core.keymem.prev_key0_reg[50]$_DFFE_PN0P_  (.D(_02830_),
    .RN(net87),
    .CK(clknet_leaf_409_clk),
    .Q(\core.keymem.prev_key0_reg[50] ),
    .QN(_19774_));
 DFFR_X1 \core.keymem.prev_key0_reg[51]$_DFFE_PN0P_  (.D(_02831_),
    .RN(net87),
    .CK(clknet_leaf_6_clk),
    .Q(\core.keymem.prev_key0_reg[51] ),
    .QN(_19773_));
 DFFR_X1 \core.keymem.prev_key0_reg[52]$_DFFE_PN0P_  (.D(_02832_),
    .RN(net86),
    .CK(clknet_leaf_405_clk),
    .Q(\core.keymem.prev_key0_reg[52] ),
    .QN(_19772_));
 DFFR_X2 \core.keymem.prev_key0_reg[53]$_DFFE_PN0P_  (.D(_02833_),
    .RN(net86),
    .CK(clknet_leaf_404_clk),
    .Q(\core.keymem.prev_key0_reg[53] ),
    .QN(_19771_));
 DFFR_X1 \core.keymem.prev_key0_reg[54]$_DFFE_PN0P_  (.D(_02834_),
    .RN(net86),
    .CK(clknet_leaf_404_clk),
    .Q(\core.keymem.prev_key0_reg[54] ),
    .QN(_19770_));
 DFFR_X1 \core.keymem.prev_key0_reg[55]$_DFFE_PN0P_  (.D(_02835_),
    .RN(net86),
    .CK(clknet_leaf_406_clk),
    .Q(\core.keymem.prev_key0_reg[55] ),
    .QN(_19769_));
 DFFR_X2 \core.keymem.prev_key0_reg[56]$_DFFE_PN0P_  (.D(_02836_),
    .RN(net87),
    .CK(clknet_leaf_415_clk),
    .Q(\core.keymem.prev_key0_reg[56] ),
    .QN(_19768_));
 DFFR_X1 \core.keymem.prev_key0_reg[57]$_DFFE_PN0P_  (.D(_02837_),
    .RN(net86),
    .CK(clknet_leaf_407_clk),
    .Q(\core.keymem.prev_key0_reg[57] ),
    .QN(_19767_));
 DFFR_X2 \core.keymem.prev_key0_reg[58]$_DFFE_PN0P_  (.D(_02838_),
    .RN(net87),
    .CK(clknet_leaf_413_clk),
    .Q(\core.keymem.prev_key0_reg[58] ),
    .QN(_19766_));
 DFFR_X1 \core.keymem.prev_key0_reg[59]$_DFFE_PN0P_  (.D(_02839_),
    .RN(net82),
    .CK(clknet_leaf_412_clk),
    .Q(\core.keymem.prev_key0_reg[59] ),
    .QN(_19765_));
 DFFR_X1 \core.keymem.prev_key0_reg[5]$_DFFE_PN0P_  (.D(_02840_),
    .RN(net82),
    .CK(clknet_leaf_5_clk),
    .Q(\core.keymem.prev_key0_reg[5] ),
    .QN(_19764_));
 DFFR_X1 \core.keymem.prev_key0_reg[60]$_DFFE_PN0P_  (.D(_02841_),
    .RN(net82),
    .CK(clknet_leaf_7_clk),
    .Q(\core.keymem.prev_key0_reg[60] ),
    .QN(_19763_));
 DFFR_X1 \core.keymem.prev_key0_reg[61]$_DFFE_PN0P_  (.D(_02842_),
    .RN(net87),
    .CK(clknet_leaf_417_clk),
    .Q(\core.keymem.prev_key0_reg[61] ),
    .QN(_19762_));
 DFFR_X1 \core.keymem.prev_key0_reg[62]$_DFFE_PN0P_  (.D(_02843_),
    .RN(net87),
    .CK(clknet_leaf_417_clk),
    .Q(\core.keymem.prev_key0_reg[62] ),
    .QN(_19761_));
 DFFR_X1 \core.keymem.prev_key0_reg[63]$_DFFE_PN0P_  (.D(_02844_),
    .RN(net82),
    .CK(clknet_leaf_420_clk),
    .Q(\core.keymem.prev_key0_reg[63] ),
    .QN(_19760_));
 DFFR_X1 \core.keymem.prev_key0_reg[64]$_DFFE_PN0P_  (.D(_02845_),
    .RN(net84),
    .CK(clknet_leaf_386_clk),
    .Q(\core.keymem.prev_key0_reg[64] ),
    .QN(_19759_));
 DFFR_X1 \core.keymem.prev_key0_reg[65]$_DFFE_PN0P_  (.D(_02846_),
    .RN(net87),
    .CK(clknet_leaf_39_clk),
    .Q(\core.keymem.prev_key0_reg[65] ),
    .QN(_19758_));
 DFFR_X1 \core.keymem.prev_key0_reg[66]$_DFFE_PN0P_  (.D(_02847_),
    .RN(net82),
    .CK(clknet_leaf_424_clk),
    .Q(\core.keymem.prev_key0_reg[66] ),
    .QN(_19757_));
 DFFR_X1 \core.keymem.prev_key0_reg[67]$_DFFE_PN0P_  (.D(_02848_),
    .RN(net82),
    .CK(clknet_leaf_420_clk),
    .Q(\core.keymem.prev_key0_reg[67] ),
    .QN(_19756_));
 DFFR_X1 \core.keymem.prev_key0_reg[68]$_DFFE_PN0P_  (.D(_02849_),
    .RN(net82),
    .CK(clknet_leaf_8_clk),
    .Q(\core.keymem.prev_key0_reg[68] ),
    .QN(_19755_));
 DFFR_X1 \core.keymem.prev_key0_reg[69]$_DFFE_PN0P_  (.D(_02850_),
    .RN(net82),
    .CK(clknet_leaf_5_clk),
    .Q(\core.keymem.prev_key0_reg[69] ),
    .QN(_19754_));
 DFFR_X1 \core.keymem.prev_key0_reg[6]$_DFFE_PN0P_  (.D(_02851_),
    .RN(net82),
    .CK(clknet_leaf_422_clk),
    .Q(\core.keymem.prev_key0_reg[6] ),
    .QN(_19753_));
 DFFR_X1 \core.keymem.prev_key0_reg[70]$_DFFE_PN0P_  (.D(_02852_),
    .RN(net82),
    .CK(clknet_leaf_423_clk),
    .Q(\core.keymem.prev_key0_reg[70] ),
    .QN(_19752_));
 DFFR_X1 \core.keymem.prev_key0_reg[71]$_DFFE_PN0P_  (.D(_02853_),
    .RN(net82),
    .CK(clknet_leaf_423_clk),
    .Q(\core.keymem.prev_key0_reg[71] ),
    .QN(_19751_));
 DFFR_X1 \core.keymem.prev_key0_reg[72]$_DFFE_PN0P_  (.D(_02854_),
    .RN(net86),
    .CK(clknet_leaf_408_clk),
    .Q(\core.keymem.prev_key0_reg[72] ),
    .QN(_19750_));
 DFFR_X2 \core.keymem.prev_key0_reg[73]$_DFFE_PN0P_  (.D(_02855_),
    .RN(net86),
    .CK(clknet_leaf_393_clk),
    .Q(\core.keymem.prev_key0_reg[73] ),
    .QN(_19749_));
 DFFR_X1 \core.keymem.prev_key0_reg[74]$_DFFE_PN0P_  (.D(_02856_),
    .RN(net86),
    .CK(clknet_leaf_407_clk),
    .Q(\core.keymem.prev_key0_reg[74] ),
    .QN(_19748_));
 DFFR_X1 \core.keymem.prev_key0_reg[75]$_DFFE_PN0P_  (.D(_02857_),
    .RN(net86),
    .CK(clknet_leaf_388_clk),
    .Q(\core.keymem.prev_key0_reg[75] ),
    .QN(_19747_));
 DFFR_X1 \core.keymem.prev_key0_reg[76]$_DFFE_PN0P_  (.D(_02858_),
    .RN(net86),
    .CK(clknet_leaf_346_clk),
    .Q(\core.keymem.prev_key0_reg[76] ),
    .QN(_19746_));
 DFFR_X1 \core.keymem.prev_key0_reg[77]$_DFFE_PN0P_  (.D(_02859_),
    .RN(net86),
    .CK(clknet_leaf_395_clk),
    .Q(\core.keymem.prev_key0_reg[77] ),
    .QN(_19745_));
 DFFR_X1 \core.keymem.prev_key0_reg[78]$_DFFE_PN0P_  (.D(_02860_),
    .RN(net86),
    .CK(clknet_leaf_347_clk),
    .Q(\core.keymem.prev_key0_reg[78] ),
    .QN(_19744_));
 DFFR_X1 \core.keymem.prev_key0_reg[79]$_DFFE_PN0P_  (.D(_02861_),
    .RN(net85),
    .CK(clknet_leaf_367_clk),
    .Q(\core.keymem.prev_key0_reg[79] ),
    .QN(_19743_));
 DFFR_X1 \core.keymem.prev_key0_reg[7]$_DFFE_PN0P_  (.D(_02862_),
    .RN(net82),
    .CK(clknet_leaf_422_clk),
    .Q(\core.keymem.prev_key0_reg[7] ),
    .QN(_19742_));
 DFFR_X1 \core.keymem.prev_key0_reg[80]$_DFFE_PN0P_  (.D(_02863_),
    .RN(net84),
    .CK(clknet_leaf_352_clk),
    .Q(\core.keymem.prev_key0_reg[80] ),
    .QN(_19741_));
 DFFR_X1 \core.keymem.prev_key0_reg[81]$_DFFE_PN0P_  (.D(_02864_),
    .RN(net85),
    .CK(clknet_leaf_367_clk),
    .Q(\core.keymem.prev_key0_reg[81] ),
    .QN(_19740_));
 DFFR_X1 \core.keymem.prev_key0_reg[82]$_DFFE_PN0P_  (.D(_02865_),
    .RN(net86),
    .CK(clknet_leaf_409_clk),
    .Q(\core.keymem.prev_key0_reg[82] ),
    .QN(_19739_));
 DFFR_X2 \core.keymem.prev_key0_reg[83]$_DFFE_PN0P_  (.D(_02866_),
    .RN(net86),
    .CK(clknet_leaf_395_clk),
    .Q(\core.keymem.prev_key0_reg[83] ),
    .QN(_19738_));
 DFFR_X1 \core.keymem.prev_key0_reg[84]$_DFFE_PN0P_  (.D(_02867_),
    .RN(net86),
    .CK(clknet_leaf_346_clk),
    .Q(\core.keymem.prev_key0_reg[84] ),
    .QN(_19737_));
 DFFR_X1 \core.keymem.prev_key0_reg[85]$_DFFE_PN0P_  (.D(_02868_),
    .RN(net86),
    .CK(clknet_leaf_347_clk),
    .Q(\core.keymem.prev_key0_reg[85] ),
    .QN(_19736_));
 DFFR_X1 \core.keymem.prev_key0_reg[86]$_DFFE_PN0P_  (.D(_02869_),
    .RN(net86),
    .CK(clknet_leaf_346_clk),
    .Q(\core.keymem.prev_key0_reg[86] ),
    .QN(_19735_));
 DFFR_X1 \core.keymem.prev_key0_reg[87]$_DFFE_PN0P_  (.D(_02870_),
    .RN(net86),
    .CK(clknet_leaf_346_clk),
    .Q(\core.keymem.prev_key0_reg[87] ),
    .QN(_19734_));
 DFFR_X1 \core.keymem.prev_key0_reg[88]$_DFFE_PN0P_  (.D(_02871_),
    .RN(net86),
    .CK(clknet_leaf_402_clk),
    .Q(\core.keymem.prev_key0_reg[88] ),
    .QN(_19733_));
 DFFR_X1 \core.keymem.prev_key0_reg[89]$_DFFE_PN0P_  (.D(_02872_),
    .RN(net86),
    .CK(clknet_leaf_407_clk),
    .Q(\core.keymem.prev_key0_reg[89] ),
    .QN(_19732_));
 DFFR_X1 \core.keymem.prev_key0_reg[8]$_DFFE_PN0P_  (.D(_02873_),
    .RN(net86),
    .CK(clknet_leaf_402_clk),
    .Q(\core.keymem.prev_key0_reg[8] ),
    .QN(_19731_));
 DFFR_X1 \core.keymem.prev_key0_reg[90]$_DFFE_PN0P_  (.D(_02874_),
    .RN(net87),
    .CK(clknet_leaf_414_clk),
    .Q(\core.keymem.prev_key0_reg[90] ),
    .QN(_19730_));
 DFFR_X1 \core.keymem.prev_key0_reg[91]$_DFFE_PN0P_  (.D(_02875_),
    .RN(net82),
    .CK(clknet_leaf_422_clk),
    .Q(\core.keymem.prev_key0_reg[91] ),
    .QN(_19729_));
 DFFR_X1 \core.keymem.prev_key0_reg[92]$_DFFE_PN0P_  (.D(_02876_),
    .RN(net82),
    .CK(clknet_leaf_423_clk),
    .Q(\core.keymem.prev_key0_reg[92] ),
    .QN(_19728_));
 DFFR_X1 \core.keymem.prev_key0_reg[93]$_DFFE_PN0P_  (.D(_02877_),
    .RN(net87),
    .CK(clknet_leaf_417_clk),
    .Q(\core.keymem.prev_key0_reg[93] ),
    .QN(_19727_));
 DFFR_X1 \core.keymem.prev_key0_reg[94]$_DFFE_PN0P_  (.D(_02878_),
    .RN(net82),
    .CK(clknet_leaf_411_clk),
    .Q(\core.keymem.prev_key0_reg[94] ),
    .QN(_19726_));
 DFFR_X1 \core.keymem.prev_key0_reg[95]$_DFFE_PN0P_  (.D(_02879_),
    .RN(net82),
    .CK(clknet_leaf_422_clk),
    .Q(\core.keymem.prev_key0_reg[95] ),
    .QN(_19725_));
 DFFR_X1 \core.keymem.prev_key0_reg[96]$_DFFE_PN0P_  (.D(_02880_),
    .RN(net88),
    .CK(clknet_leaf_387_clk),
    .Q(\core.keymem.prev_key0_reg[96] ),
    .QN(_19724_));
 DFFR_X1 \core.keymem.prev_key0_reg[97]$_DFFE_PN0P_  (.D(_02881_),
    .RN(net87),
    .CK(clknet_leaf_39_clk),
    .Q(\core.keymem.prev_key0_reg[97] ),
    .QN(_19723_));
 DFFR_X1 \core.keymem.prev_key0_reg[98]$_DFFE_PN0P_  (.D(_02882_),
    .RN(net82),
    .CK(clknet_leaf_424_clk),
    .Q(\core.keymem.prev_key0_reg[98] ),
    .QN(_19722_));
 DFFR_X1 \core.keymem.prev_key0_reg[99]$_DFFE_PN0P_  (.D(_02883_),
    .RN(net82),
    .CK(clknet_leaf_424_clk),
    .Q(\core.keymem.prev_key0_reg[99] ),
    .QN(_19721_));
 DFFR_X1 \core.keymem.prev_key0_reg[9]$_DFFE_PN0P_  (.D(_02884_),
    .RN(net86),
    .CK(clknet_leaf_398_clk),
    .Q(\core.keymem.prev_key0_reg[9] ),
    .QN(_19720_));
 DFFR_X1 \core.keymem.prev_key1_reg[0]$_DFFE_PN0P_  (.D(_02885_),
    .RN(net86),
    .CK(clknet_leaf_405_clk),
    .Q(\core.keymem.prev_key1_reg[0] ),
    .QN(_19719_));
 DFFR_X1 \core.keymem.prev_key1_reg[100]$_DFFE_PN0P_  (.D(_02886_),
    .RN(net82),
    .CK(clknet_leaf_7_clk),
    .Q(\core.keymem.prev_key1_reg[100] ),
    .QN(_00128_));
 DFFR_X1 \core.keymem.prev_key1_reg[101]$_DFFE_PN0P_  (.D(_02887_),
    .RN(net82),
    .CK(clknet_leaf_6_clk),
    .Q(\core.keymem.prev_key1_reg[101] ),
    .QN(_00377_));
 DFFR_X1 \core.keymem.prev_key1_reg[102]$_DFFE_PN0P_  (.D(_02888_),
    .RN(net82),
    .CK(clknet_leaf_419_clk),
    .Q(\core.keymem.prev_key1_reg[102] ),
    .QN(_00379_));
 DFFR_X1 \core.keymem.prev_key1_reg[103]$_DFFE_PN0P_  (.D(_02889_),
    .RN(net82),
    .CK(clknet_leaf_419_clk),
    .Q(\core.keymem.prev_key1_reg[103] ),
    .QN(_00132_));
 DFFR_X1 \core.keymem.prev_key1_reg[104]$_DFFE_PN0P_  (.D(_02890_),
    .RN(net86),
    .CK(clknet_leaf_397_clk),
    .Q(\core.keymem.prev_key1_reg[104] ),
    .QN(_19718_));
 DFFR_X1 \core.keymem.prev_key1_reg[105]$_DFFE_PN0P_  (.D(_02891_),
    .RN(net84),
    .CK(clknet_leaf_352_clk),
    .Q(\core.keymem.prev_key1_reg[105] ),
    .QN(_19717_));
 DFFR_X1 \core.keymem.prev_key1_reg[106]$_DFFE_PN0P_  (.D(_02892_),
    .RN(net86),
    .CK(clknet_leaf_397_clk),
    .Q(\core.keymem.prev_key1_reg[106] ),
    .QN(_00136_));
 DFFR_X1 \core.keymem.prev_key1_reg[107]$_DFFE_PN0P_  (.D(_02893_),
    .RN(net84),
    .CK(clknet_leaf_352_clk),
    .Q(\core.keymem.prev_key1_reg[107] ),
    .QN(_00138_));
 DFFR_X1 \core.keymem.prev_key1_reg[108]$_DFFE_PN0P_  (.D(_02894_),
    .RN(net84),
    .CK(clknet_leaf_353_clk),
    .Q(\core.keymem.prev_key1_reg[108] ),
    .QN(_00140_));
 DFFR_X1 \core.keymem.prev_key1_reg[109]$_DFFE_PN0P_  (.D(_02895_),
    .RN(net88),
    .CK(clknet_leaf_399_clk),
    .Q(\core.keymem.prev_key1_reg[109] ),
    .QN(_19716_));
 DFFR_X1 \core.keymem.prev_key1_reg[10]$_DFFE_PN0P_  (.D(_02896_),
    .RN(net86),
    .CK(clknet_leaf_398_clk),
    .Q(\core.keymem.prev_key1_reg[10] ),
    .QN(_00398_));
 DFFR_X1 \core.keymem.prev_key1_reg[110]$_DFFE_PN0P_  (.D(_02897_),
    .RN(net84),
    .CK(clknet_leaf_350_clk),
    .Q(\core.keymem.prev_key1_reg[110] ),
    .QN(_19715_));
 DFFR_X1 \core.keymem.prev_key1_reg[111]$_DFFE_PN0P_  (.D(_02898_),
    .RN(net85),
    .CK(clknet_leaf_366_clk),
    .Q(\core.keymem.prev_key1_reg[111] ),
    .QN(_00144_));
 DFFR_X1 \core.keymem.prev_key1_reg[112]$_DFFE_PN0P_  (.D(_02899_),
    .RN(net84),
    .CK(clknet_leaf_352_clk),
    .Q(\core.keymem.prev_key1_reg[112] ),
    .QN(_19714_));
 DFFR_X1 \core.keymem.prev_key1_reg[113]$_DFFE_PN0P_  (.D(_02900_),
    .RN(net84),
    .CK(clknet_leaf_352_clk),
    .Q(\core.keymem.prev_key1_reg[113] ),
    .QN(_19713_));
 DFFR_X1 \core.keymem.prev_key1_reg[114]$_DFFE_PN0P_  (.D(_02901_),
    .RN(net86),
    .CK(clknet_leaf_396_clk),
    .Q(\core.keymem.prev_key1_reg[114] ),
    .QN(_00148_));
 DFFR_X2 \core.keymem.prev_key1_reg[115]$_DFFE_PN0P_  (.D(_02902_),
    .RN(net84),
    .CK(clknet_leaf_350_clk),
    .Q(\core.keymem.prev_key1_reg[115] ),
    .QN(_00150_));
 DFFR_X1 \core.keymem.prev_key1_reg[116]$_DFFE_PN0P_  (.D(_02903_),
    .RN(net84),
    .CK(clknet_leaf_349_clk),
    .Q(\core.keymem.prev_key1_reg[116] ),
    .QN(_00152_));
 DFFR_X1 \core.keymem.prev_key1_reg[117]$_DFFE_PN0P_  (.D(_02904_),
    .RN(net86),
    .CK(clknet_leaf_347_clk),
    .Q(\core.keymem.prev_key1_reg[117] ),
    .QN(_19712_));
 DFFR_X1 \core.keymem.prev_key1_reg[118]$_DFFE_PN0P_  (.D(_02905_),
    .RN(net86),
    .CK(clknet_leaf_347_clk),
    .Q(\core.keymem.prev_key1_reg[118] ),
    .QN(_19711_));
 DFFR_X1 \core.keymem.prev_key1_reg[119]$_DFFE_PN0P_  (.D(_02906_),
    .RN(net84),
    .CK(clknet_leaf_349_clk),
    .Q(\core.keymem.prev_key1_reg[119] ),
    .QN(_00156_));
 DFFR_X2 \core.keymem.prev_key1_reg[11]$_DFFE_PN0P_  (.D(_02907_),
    .RN(net88),
    .CK(clknet_leaf_387_clk),
    .Q(\core.keymem.prev_key1_reg[11] ),
    .QN(_00401_));
 DFFR_X1 \core.keymem.prev_key1_reg[120]$_DFFE_PN0P_  (.D(_02908_),
    .RN(net86),
    .CK(clknet_leaf_402_clk),
    .Q(\core.keymem.prev_key1_reg[120] ),
    .QN(_00018_));
 DFFR_X1 \core.keymem.prev_key1_reg[121]$_DFFE_PN0P_  (.D(_02909_),
    .RN(net86),
    .CK(clknet_leaf_415_clk),
    .Q(\core.keymem.prev_key1_reg[121] ),
    .QN(_00021_));
 DFFR_X1 \core.keymem.prev_key1_reg[122]$_DFFE_PN0P_  (.D(_02910_),
    .RN(net87),
    .CK(clknet_leaf_415_clk),
    .Q(\core.keymem.prev_key1_reg[122] ),
    .QN(_00024_));
 DFFR_X1 \core.keymem.prev_key1_reg[123]$_DFFE_PN0P_  (.D(_02911_),
    .RN(net87),
    .CK(clknet_leaf_412_clk),
    .Q(\core.keymem.prev_key1_reg[123] ),
    .QN(_00027_));
 DFFR_X1 \core.keymem.prev_key1_reg[124]$_DFFE_PN0P_  (.D(_02912_),
    .RN(net87),
    .CK(clknet_leaf_7_clk),
    .Q(\core.keymem.prev_key1_reg[124] ),
    .QN(_00030_));
 DFFR_X1 \core.keymem.prev_key1_reg[125]$_DFFE_PN0P_  (.D(_02913_),
    .RN(net87),
    .CK(clknet_leaf_416_clk),
    .Q(\core.keymem.prev_key1_reg[125] ),
    .QN(_00033_));
 DFFR_X1 \core.keymem.prev_key1_reg[126]$_DFFE_PN0P_  (.D(_02914_),
    .RN(net82),
    .CK(clknet_leaf_418_clk),
    .Q(\core.keymem.prev_key1_reg[126] ),
    .QN(_00036_));
 DFFR_X1 \core.keymem.prev_key1_reg[127]$_DFFE_PN0P_  (.D(_02915_),
    .RN(net82),
    .CK(clknet_leaf_420_clk),
    .Q(\core.keymem.prev_key1_reg[127] ),
    .QN(_00039_));
 DFFR_X1 \core.keymem.prev_key1_reg[12]$_DFFE_PN0P_  (.D(_02916_),
    .RN(net86),
    .CK(clknet_leaf_399_clk),
    .Q(\core.keymem.prev_key1_reg[12] ),
    .QN(_19710_));
 DFFR_X2 \core.keymem.prev_key1_reg[13]$_DFFE_PN0P_  (.D(_02917_),
    .RN(net86),
    .CK(clknet_leaf_392_clk),
    .Q(\core.keymem.prev_key1_reg[13] ),
    .QN(_00384_));
 DFFR_X2 \core.keymem.prev_key1_reg[14]$_DFFE_PN0P_  (.D(_02918_),
    .RN(net86),
    .CK(clknet_leaf_346_clk),
    .Q(\core.keymem.prev_key1_reg[14] ),
    .QN(_00387_));
 DFFR_X2 \core.keymem.prev_key1_reg[15]$_DFFE_PN0P_  (.D(_02919_),
    .RN(net86),
    .CK(clknet_leaf_405_clk),
    .Q(\core.keymem.prev_key1_reg[15] ),
    .QN(_00390_));
 DFFR_X1 \core.keymem.prev_key1_reg[16]$_DFFE_PN0P_  (.D(_02920_),
    .RN(net84),
    .CK(clknet_leaf_353_clk),
    .Q(\core.keymem.prev_key1_reg[16] ),
    .QN(_19709_));
 DFFR_X1 \core.keymem.prev_key1_reg[17]$_DFFE_PN0P_  (.D(_02921_),
    .RN(net88),
    .CK(clknet_leaf_387_clk),
    .Q(\core.keymem.prev_key1_reg[17] ),
    .QN(_00425_));
 DFFR_X1 \core.keymem.prev_key1_reg[18]$_DFFE_PN0P_  (.D(_02922_),
    .RN(net86),
    .CK(clknet_leaf_392_clk),
    .Q(\core.keymem.prev_key1_reg[18] ),
    .QN(_00428_));
 DFFR_X1 \core.keymem.prev_key1_reg[19]$_DFFE_PN0P_  (.D(_02923_),
    .RN(net86),
    .CK(clknet_leaf_393_clk),
    .Q(\core.keymem.prev_key1_reg[19] ),
    .QN(_00431_));
 DFFR_X1 \core.keymem.prev_key1_reg[1]$_DFFE_PN0P_  (.D(_02924_),
    .RN(net86),
    .CK(clknet_leaf_393_clk),
    .Q(\core.keymem.prev_key1_reg[1] ),
    .QN(_00362_));
 DFFR_X1 \core.keymem.prev_key1_reg[20]$_DFFE_PN0P_  (.D(_02925_),
    .RN(net86),
    .CK(clknet_leaf_401_clk),
    .Q(\core.keymem.prev_key1_reg[20] ),
    .QN(_19708_));
 DFFR_X2 \core.keymem.prev_key1_reg[21]$_DFFE_PN0P_  (.D(_02926_),
    .RN(net86),
    .CK(clknet_leaf_401_clk),
    .Q(\core.keymem.prev_key1_reg[21] ),
    .QN(_00414_));
 DFFR_X2 \core.keymem.prev_key1_reg[22]$_DFFE_PN0P_  (.D(_02927_),
    .RN(net86),
    .CK(clknet_leaf_405_clk),
    .Q(\core.keymem.prev_key1_reg[22] ),
    .QN(_00417_));
 DFFR_X2 \core.keymem.prev_key1_reg[23]$_DFFE_PN0P_  (.D(_02928_),
    .RN(net86),
    .CK(clknet_leaf_406_clk),
    .Q(\core.keymem.prev_key1_reg[23] ),
    .QN(_00420_));
 DFFR_X1 \core.keymem.prev_key1_reg[24]$_DFFE_PN0P_  (.D(_02929_),
    .RN(net86),
    .CK(clknet_leaf_414_clk),
    .Q(\core.keymem.prev_key1_reg[24] ),
    .QN(_19707_));
 DFFR_X1 \core.keymem.prev_key1_reg[25]$_DFFE_PN0P_  (.D(_02930_),
    .RN(net86),
    .CK(clknet_leaf_415_clk),
    .Q(\core.keymem.prev_key1_reg[25] ),
    .QN(_00342_));
 DFFR_X1 \core.keymem.prev_key1_reg[26]$_DFFE_PN0P_  (.D(_02931_),
    .RN(net87),
    .CK(clknet_leaf_416_clk),
    .Q(\core.keymem.prev_key1_reg[26] ),
    .QN(_00345_));
 DFFR_X1 \core.keymem.prev_key1_reg[27]$_DFFE_PN0P_  (.D(_02932_),
    .RN(net87),
    .CK(clknet_leaf_412_clk),
    .Q(\core.keymem.prev_key1_reg[27] ),
    .QN(_00346_));
 DFFR_X1 \core.keymem.prev_key1_reg[28]$_DFFE_PN0P_  (.D(_02933_),
    .RN(net82),
    .CK(clknet_leaf_420_clk),
    .Q(\core.keymem.prev_key1_reg[28] ),
    .QN(_19706_));
 DFFR_X2 \core.keymem.prev_key1_reg[29]$_DFFE_PN0P_  (.D(_02934_),
    .RN(net82),
    .CK(clknet_leaf_421_clk),
    .Q(\core.keymem.prev_key1_reg[29] ),
    .QN(_00332_));
 DFFR_X1 \core.keymem.prev_key1_reg[2]$_DFFE_PN0P_  (.D(_02935_),
    .RN(net87),
    .CK(clknet_leaf_395_clk),
    .Q(\core.keymem.prev_key1_reg[2] ),
    .QN(_00365_));
 DFFR_X2 \core.keymem.prev_key1_reg[30]$_DFFE_PN0P_  (.D(_02936_),
    .RN(net82),
    .CK(clknet_leaf_411_clk),
    .Q(\core.keymem.prev_key1_reg[30] ),
    .QN(_00335_));
 DFFR_X2 \core.keymem.prev_key1_reg[31]$_DFFE_PN0P_  (.D(_02937_),
    .RN(net82),
    .CK(clknet_leaf_421_clk),
    .Q(\core.keymem.prev_key1_reg[31] ),
    .QN(_00338_));
 DFFR_X1 \core.keymem.prev_key1_reg[32]$_DFFE_PN0P_  (.D(_02938_),
    .RN(net88),
    .CK(clknet_leaf_386_clk),
    .Q(\core.keymem.prev_key1_reg[32] ),
    .QN(_19705_));
 DFFR_X1 \core.keymem.prev_key1_reg[33]$_DFFE_PN0P_  (.D(_02939_),
    .RN(net87),
    .CK(clknet_leaf_38_clk),
    .Q(\core.keymem.prev_key1_reg[33] ),
    .QN(_19704_));
 DFFR_X1 \core.keymem.prev_key1_reg[34]$_DFFE_PN0P_  (.D(_02940_),
    .RN(net82),
    .CK(clknet_leaf_5_clk),
    .Q(\core.keymem.prev_key1_reg[34] ),
    .QN(_19703_));
 DFFR_X1 \core.keymem.prev_key1_reg[35]$_DFFE_PN0P_  (.D(_02941_),
    .RN(net82),
    .CK(clknet_leaf_3_clk),
    .Q(\core.keymem.prev_key1_reg[35] ),
    .QN(_19702_));
 DFFR_X1 \core.keymem.prev_key1_reg[36]$_DFFE_PN0P_  (.D(_02942_),
    .RN(net82),
    .CK(clknet_leaf_9_clk),
    .Q(\core.keymem.prev_key1_reg[36] ),
    .QN(_19701_));
 DFFR_X1 \core.keymem.prev_key1_reg[37]$_DFFE_PN0P_  (.D(_02943_),
    .RN(net82),
    .CK(clknet_leaf_8_clk),
    .Q(\core.keymem.prev_key1_reg[37] ),
    .QN(_19700_));
 DFFR_X1 \core.keymem.prev_key1_reg[38]$_DFFE_PN0P_  (.D(_02944_),
    .RN(net82),
    .CK(clknet_leaf_4_clk),
    .Q(\core.keymem.prev_key1_reg[38] ),
    .QN(_19699_));
 DFFR_X1 \core.keymem.prev_key1_reg[39]$_DFFE_PN0P_  (.D(_02945_),
    .RN(net82),
    .CK(clknet_leaf_418_clk),
    .Q(\core.keymem.prev_key1_reg[39] ),
    .QN(_19698_));
 DFFR_X1 \core.keymem.prev_key1_reg[3]$_DFFE_PN0P_  (.D(_02946_),
    .RN(net82),
    .CK(clknet_leaf_418_clk),
    .Q(\core.keymem.prev_key1_reg[3] ),
    .QN(_00368_));
 DFFR_X1 \core.keymem.prev_key1_reg[40]$_DFFE_PN0P_  (.D(_02947_),
    .RN(net86),
    .CK(clknet_leaf_396_clk),
    .Q(\core.keymem.prev_key1_reg[40] ),
    .QN(_19697_));
 DFFR_X1 \core.keymem.prev_key1_reg[41]$_DFFE_PN0P_  (.D(_02948_),
    .RN(net86),
    .CK(clknet_leaf_39_clk),
    .Q(\core.keymem.prev_key1_reg[41] ),
    .QN(_19696_));
 DFFR_X2 \core.keymem.prev_key1_reg[42]$_DFFE_PN0P_  (.D(_02949_),
    .RN(net86),
    .CK(clknet_leaf_398_clk),
    .Q(\core.keymem.prev_key1_reg[42] ),
    .QN(_19695_));
 DFFR_X1 \core.keymem.prev_key1_reg[43]$_DFFE_PN0P_  (.D(_02950_),
    .RN(net88),
    .CK(clknet_leaf_388_clk),
    .Q(\core.keymem.prev_key1_reg[43] ),
    .QN(_19694_));
 DFFR_X2 \core.keymem.prev_key1_reg[44]$_DFFE_PN0P_  (.D(_02951_),
    .RN(net88),
    .CK(clknet_leaf_399_clk),
    .Q(\core.keymem.prev_key1_reg[44] ),
    .QN(_19693_));
 DFFR_X1 \core.keymem.prev_key1_reg[45]$_DFFE_PN0P_  (.D(_02952_),
    .RN(net86),
    .CK(clknet_leaf_391_clk),
    .Q(\core.keymem.prev_key1_reg[45] ),
    .QN(_19692_));
 DFFR_X1 \core.keymem.prev_key1_reg[46]$_DFFE_PN0P_  (.D(_02953_),
    .RN(net84),
    .CK(clknet_leaf_350_clk),
    .Q(\core.keymem.prev_key1_reg[46] ),
    .QN(_19691_));
 DFFR_X1 \core.keymem.prev_key1_reg[47]$_DFFE_PN0P_  (.D(_02954_),
    .RN(net84),
    .CK(clknet_leaf_386_clk),
    .Q(\core.keymem.prev_key1_reg[47] ),
    .QN(_19690_));
 DFFR_X1 \core.keymem.prev_key1_reg[48]$_DFFE_PN0P_  (.D(_02955_),
    .RN(net88),
    .CK(clknet_leaf_351_clk),
    .Q(\core.keymem.prev_key1_reg[48] ),
    .QN(_19689_));
 DFFR_X1 \core.keymem.prev_key1_reg[49]$_DFFE_PN0P_  (.D(_02956_),
    .RN(net88),
    .CK(clknet_leaf_387_clk),
    .Q(\core.keymem.prev_key1_reg[49] ),
    .QN(_19688_));
 DFFR_X1 \core.keymem.prev_key1_reg[4]$_DFFE_PN0P_  (.D(_02957_),
    .RN(net82),
    .CK(clknet_leaf_7_clk),
    .Q(\core.keymem.prev_key1_reg[4] ),
    .QN(_19687_));
 DFFR_X1 \core.keymem.prev_key1_reg[50]$_DFFE_PN0P_  (.D(_02958_),
    .RN(net86),
    .CK(clknet_leaf_395_clk),
    .Q(\core.keymem.prev_key1_reg[50] ),
    .QN(_19686_));
 DFFR_X1 \core.keymem.prev_key1_reg[51]$_DFFE_PN0P_  (.D(_02959_),
    .RN(net87),
    .CK(clknet_leaf_6_clk),
    .Q(\core.keymem.prev_key1_reg[51] ),
    .QN(_19685_));
 DFFR_X1 \core.keymem.prev_key1_reg[52]$_DFFE_PN0P_  (.D(_02960_),
    .RN(net86),
    .CK(clknet_leaf_401_clk),
    .Q(\core.keymem.prev_key1_reg[52] ),
    .QN(_19684_));
 DFFR_X1 \core.keymem.prev_key1_reg[53]$_DFFE_PN0P_  (.D(_02961_),
    .RN(net86),
    .CK(clknet_leaf_400_clk),
    .Q(\core.keymem.prev_key1_reg[53] ),
    .QN(_19683_));
 DFFR_X1 \core.keymem.prev_key1_reg[54]$_DFFE_PN0P_  (.D(_02962_),
    .RN(net86),
    .CK(clknet_leaf_401_clk),
    .Q(\core.keymem.prev_key1_reg[54] ),
    .QN(_19682_));
 DFFR_X1 \core.keymem.prev_key1_reg[55]$_DFFE_PN0P_  (.D(_02963_),
    .RN(net86),
    .CK(clknet_leaf_401_clk),
    .Q(\core.keymem.prev_key1_reg[55] ),
    .QN(_19681_));
 DFFR_X1 \core.keymem.prev_key1_reg[56]$_DFFE_PN0P_  (.D(_02964_),
    .RN(net86),
    .CK(clknet_leaf_396_clk),
    .Q(\core.keymem.prev_key1_reg[56] ),
    .QN(_19680_));
 DFFR_X1 \core.keymem.prev_key1_reg[57]$_DFFE_PN0P_  (.D(_02965_),
    .RN(net86),
    .CK(clknet_leaf_396_clk),
    .Q(\core.keymem.prev_key1_reg[57] ),
    .QN(_19679_));
 DFFR_X1 \core.keymem.prev_key1_reg[58]$_DFFE_PN0P_  (.D(_02966_),
    .RN(net87),
    .CK(clknet_leaf_416_clk),
    .Q(\core.keymem.prev_key1_reg[58] ),
    .QN(_19678_));
 DFFR_X1 \core.keymem.prev_key1_reg[59]$_DFFE_PN0P_  (.D(_02967_),
    .RN(net87),
    .CK(clknet_leaf_416_clk),
    .Q(\core.keymem.prev_key1_reg[59] ),
    .QN(_19677_));
 DFFR_X1 \core.keymem.prev_key1_reg[5]$_DFFE_PN0P_  (.D(_02968_),
    .RN(net82),
    .CK(clknet_leaf_5_clk),
    .Q(\core.keymem.prev_key1_reg[5] ),
    .QN(_00351_));
 DFFR_X1 \core.keymem.prev_key1_reg[60]$_DFFE_PN0P_  (.D(_02969_),
    .RN(net87),
    .CK(clknet_leaf_38_clk),
    .Q(\core.keymem.prev_key1_reg[60] ),
    .QN(_19676_));
 DFFR_X1 \core.keymem.prev_key1_reg[61]$_DFFE_PN0P_  (.D(_02970_),
    .RN(net87),
    .CK(clknet_leaf_6_clk),
    .Q(\core.keymem.prev_key1_reg[61] ),
    .QN(_19675_));
 DFFR_X1 \core.keymem.prev_key1_reg[62]$_DFFE_PN0P_  (.D(_02971_),
    .RN(net87),
    .CK(clknet_leaf_417_clk),
    .Q(\core.keymem.prev_key1_reg[62] ),
    .QN(_19674_));
 DFFR_X1 \core.keymem.prev_key1_reg[63]$_DFFE_PN0P_  (.D(_02972_),
    .RN(net82),
    .CK(clknet_leaf_418_clk),
    .Q(\core.keymem.prev_key1_reg[63] ),
    .QN(_19673_));
 DFFR_X1 \core.keymem.prev_key1_reg[64]$_DFFE_PN0P_  (.D(_02973_),
    .RN(net84),
    .CK(clknet_leaf_386_clk),
    .Q(\core.keymem.prev_key1_reg[64] ),
    .QN(_19672_));
 DFFR_X1 \core.keymem.prev_key1_reg[65]$_DFFE_PN0P_  (.D(_02974_),
    .RN(net87),
    .CK(clknet_leaf_38_clk),
    .Q(\core.keymem.prev_key1_reg[65] ),
    .QN(_19671_));
 DFFR_X1 \core.keymem.prev_key1_reg[66]$_DFFE_PN0P_  (.D(_02975_),
    .RN(net82),
    .CK(clknet_leaf_5_clk),
    .Q(\core.keymem.prev_key1_reg[66] ),
    .QN(_19670_));
 DFFR_X1 \core.keymem.prev_key1_reg[67]$_DFFE_PN0P_  (.D(_02976_),
    .RN(net82),
    .CK(clknet_leaf_419_clk),
    .Q(\core.keymem.prev_key1_reg[67] ),
    .QN(_19669_));
 DFFR_X1 \core.keymem.prev_key1_reg[68]$_DFFE_PN0P_  (.D(_02977_),
    .RN(net82),
    .CK(clknet_leaf_8_clk),
    .Q(\core.keymem.prev_key1_reg[68] ),
    .QN(_19668_));
 DFFR_X1 \core.keymem.prev_key1_reg[69]$_DFFE_PN0P_  (.D(_02978_),
    .RN(net82),
    .CK(clknet_leaf_7_clk),
    .Q(\core.keymem.prev_key1_reg[69] ),
    .QN(_19667_));
 DFFR_X2 \core.keymem.prev_key1_reg[6]$_DFFE_PN0P_  (.D(_02979_),
    .RN(net86),
    .CK(clknet_leaf_406_clk),
    .Q(\core.keymem.prev_key1_reg[6] ),
    .QN(_00354_));
 DFFR_X1 \core.keymem.prev_key1_reg[70]$_DFFE_PN0P_  (.D(_02980_),
    .RN(net82),
    .CK(clknet_leaf_4_clk),
    .Q(\core.keymem.prev_key1_reg[70] ),
    .QN(_19666_));
 DFFR_X1 \core.keymem.prev_key1_reg[71]$_DFFE_PN0P_  (.D(_02981_),
    .RN(net82),
    .CK(clknet_leaf_418_clk),
    .Q(\core.keymem.prev_key1_reg[71] ),
    .QN(_19665_));
 DFFR_X1 \core.keymem.prev_key1_reg[72]$_DFFE_PN0P_  (.D(_02982_),
    .RN(net86),
    .CK(clknet_leaf_397_clk),
    .Q(\core.keymem.prev_key1_reg[72] ),
    .QN(_19664_));
 DFFR_X1 \core.keymem.prev_key1_reg[73]$_DFFE_PN0P_  (.D(_02983_),
    .RN(net86),
    .CK(clknet_leaf_391_clk),
    .Q(\core.keymem.prev_key1_reg[73] ),
    .QN(_19663_));
 DFFR_X1 \core.keymem.prev_key1_reg[74]$_DFFE_PN0P_  (.D(_02984_),
    .RN(net86),
    .CK(clknet_leaf_398_clk),
    .Q(\core.keymem.prev_key1_reg[74] ),
    .QN(_19662_));
 DFFR_X1 \core.keymem.prev_key1_reg[75]$_DFFE_PN0P_  (.D(_02985_),
    .RN(net86),
    .CK(clknet_leaf_388_clk),
    .Q(\core.keymem.prev_key1_reg[75] ),
    .QN(_19661_));
 DFFR_X1 \core.keymem.prev_key1_reg[76]$_DFFE_PN0P_  (.D(_02986_),
    .RN(net84),
    .CK(clknet_leaf_353_clk),
    .Q(\core.keymem.prev_key1_reg[76] ),
    .QN(_19660_));
 DFFR_X1 \core.keymem.prev_key1_reg[77]$_DFFE_PN0P_  (.D(_02987_),
    .RN(net88),
    .CK(clknet_leaf_392_clk),
    .Q(\core.keymem.prev_key1_reg[77] ),
    .QN(_19659_));
 DFFR_X1 \core.keymem.prev_key1_reg[78]$_DFFE_PN0P_  (.D(_02988_),
    .RN(net84),
    .CK(clknet_leaf_351_clk),
    .Q(\core.keymem.prev_key1_reg[78] ),
    .QN(_19658_));
 DFFR_X1 \core.keymem.prev_key1_reg[79]$_DFFE_PN0P_  (.D(_02989_),
    .RN(net85),
    .CK(clknet_leaf_367_clk),
    .Q(\core.keymem.prev_key1_reg[79] ),
    .QN(_19657_));
 DFFR_X2 \core.keymem.prev_key1_reg[7]$_DFFE_PN0P_  (.D(_02990_),
    .RN(net86),
    .CK(clknet_leaf_415_clk),
    .Q(\core.keymem.prev_key1_reg[7] ),
    .QN(_00357_));
 DFFR_X1 \core.keymem.prev_key1_reg[80]$_DFFE_PN0P_  (.D(_02991_),
    .RN(net84),
    .CK(clknet_leaf_367_clk),
    .Q(\core.keymem.prev_key1_reg[80] ),
    .QN(_19656_));
 DFFR_X1 \core.keymem.prev_key1_reg[81]$_DFFE_PN0P_  (.D(_02992_),
    .RN(net85),
    .CK(clknet_leaf_367_clk),
    .Q(\core.keymem.prev_key1_reg[81] ),
    .QN(_19655_));
 DFFR_X1 \core.keymem.prev_key1_reg[82]$_DFFE_PN0P_  (.D(_02993_),
    .RN(net86),
    .CK(clknet_leaf_396_clk),
    .Q(\core.keymem.prev_key1_reg[82] ),
    .QN(_19654_));
 DFFR_X1 \core.keymem.prev_key1_reg[83]$_DFFE_PN0P_  (.D(_02994_),
    .RN(net86),
    .CK(clknet_leaf_396_clk),
    .Q(\core.keymem.prev_key1_reg[83] ),
    .QN(_19653_));
 DFFR_X1 \core.keymem.prev_key1_reg[84]$_DFFE_PN0P_  (.D(_02995_),
    .RN(net84),
    .CK(clknet_leaf_350_clk),
    .Q(\core.keymem.prev_key1_reg[84] ),
    .QN(_19652_));
 DFFR_X1 \core.keymem.prev_key1_reg[85]$_DFFE_PN0P_  (.D(_02996_),
    .RN(net84),
    .CK(clknet_leaf_351_clk),
    .Q(\core.keymem.prev_key1_reg[85] ),
    .QN(_19651_));
 DFFR_X1 \core.keymem.prev_key1_reg[86]$_DFFE_PN0P_  (.D(_02997_),
    .RN(net86),
    .CK(clknet_leaf_347_clk),
    .Q(\core.keymem.prev_key1_reg[86] ),
    .QN(_19650_));
 DFFR_X1 \core.keymem.prev_key1_reg[87]$_DFFE_PN0P_  (.D(_02998_),
    .RN(net84),
    .CK(clknet_leaf_350_clk),
    .Q(\core.keymem.prev_key1_reg[87] ),
    .QN(_19649_));
 DFFR_X1 \core.keymem.prev_key1_reg[88]$_DFFE_PN0P_  (.D(_02999_),
    .RN(net86),
    .CK(clknet_leaf_397_clk),
    .Q(\core.keymem.prev_key1_reg[88] ),
    .QN(_19648_));
 DFFR_X1 \core.keymem.prev_key1_reg[89]$_DFFE_PN0P_  (.D(_03000_),
    .RN(net86),
    .CK(clknet_leaf_397_clk),
    .Q(\core.keymem.prev_key1_reg[89] ),
    .QN(_19647_));
 DFFR_X1 \core.keymem.prev_key1_reg[8]$_DFFE_PN0P_  (.D(_03001_),
    .RN(net86),
    .CK(clknet_leaf_407_clk),
    .Q(\core.keymem.prev_key1_reg[8] ),
    .QN(_19646_));
 DFFR_X1 \core.keymem.prev_key1_reg[90]$_DFFE_PN0P_  (.D(_03002_),
    .RN(net87),
    .CK(clknet_leaf_416_clk),
    .Q(\core.keymem.prev_key1_reg[90] ),
    .QN(_19645_));
 DFFR_X1 \core.keymem.prev_key1_reg[91]$_DFFE_PN0P_  (.D(_03003_),
    .RN(net87),
    .CK(clknet_leaf_417_clk),
    .Q(\core.keymem.prev_key1_reg[91] ),
    .QN(_19644_));
 DFFR_X1 \core.keymem.prev_key1_reg[92]$_DFFE_PN0P_  (.D(_03004_),
    .RN(net87),
    .CK(clknet_leaf_38_clk),
    .Q(\core.keymem.prev_key1_reg[92] ),
    .QN(_19643_));
 DFFR_X1 \core.keymem.prev_key1_reg[93]$_DFFE_PN0P_  (.D(_03005_),
    .RN(net87),
    .CK(clknet_leaf_394_clk),
    .Q(\core.keymem.prev_key1_reg[93] ),
    .QN(_19642_));
 DFFR_X1 \core.keymem.prev_key1_reg[94]$_DFFE_PN0P_  (.D(_03006_),
    .RN(net87),
    .CK(clknet_leaf_417_clk),
    .Q(\core.keymem.prev_key1_reg[94] ),
    .QN(_19641_));
 DFFR_X1 \core.keymem.prev_key1_reg[95]$_DFFE_PN0P_  (.D(_03007_),
    .RN(net82),
    .CK(clknet_leaf_418_clk),
    .Q(\core.keymem.prev_key1_reg[95] ),
    .QN(_19640_));
 DFFR_X1 \core.keymem.prev_key1_reg[96]$_DFFE_PN0P_  (.D(_03008_),
    .RN(net88),
    .CK(clknet_leaf_387_clk),
    .Q(\core.keymem.prev_key1_reg[96] ),
    .QN(_00328_));
 DFFR_X1 \core.keymem.prev_key1_reg[97]$_DFFE_PN0P_  (.D(_03009_),
    .RN(net87),
    .CK(clknet_leaf_39_clk),
    .Q(\core.keymem.prev_key1_reg[97] ),
    .QN(_00372_));
 DFFR_X1 \core.keymem.prev_key1_reg[98]$_DFFE_PN0P_  (.D(_03010_),
    .RN(net82),
    .CK(clknet_leaf_6_clk),
    .Q(\core.keymem.prev_key1_reg[98] ),
    .QN(_00124_));
 DFFR_X1 \core.keymem.prev_key1_reg[99]$_DFFE_PN0P_  (.D(_03011_),
    .RN(net82),
    .CK(clknet_leaf_419_clk),
    .Q(\core.keymem.prev_key1_reg[99] ),
    .QN(_00126_));
 DFFR_X2 \core.keymem.prev_key1_reg[9]$_DFFE_PN0P_  (.D(_03012_),
    .RN(net86),
    .CK(clknet_leaf_399_clk),
    .Q(\core.keymem.prev_key1_reg[9] ),
    .QN(_00395_));
 DFFR_X1 \core.keymem.rcon_reg[0]$_DFFE_PN0P_  (.D(_03013_),
    .RN(net87),
    .CK(clknet_leaf_410_clk),
    .Q(\core.keymem.rcon_reg[0] ),
    .QN(_19639_));
 DFFR_X1 \core.keymem.rcon_reg[1]$_DFFE_PN0P_  (.D(_03014_),
    .RN(net87),
    .CK(clknet_leaf_410_clk),
    .Q(\core.keymem.rcon_logic.tmp_rcon[2] ),
    .QN(_19638_));
 DFFR_X1 \core.keymem.rcon_reg[2]$_DFFE_PN0P_  (.D(_03015_),
    .RN(net87),
    .CK(clknet_leaf_410_clk),
    .Q(\core.keymem.rcon_reg[2] ),
    .QN(_19637_));
 DFFR_X1 \core.keymem.rcon_reg[3]$_DFFE_PN0P_  (.D(_03016_),
    .RN(net87),
    .CK(clknet_leaf_410_clk),
    .Q(\core.keymem.rcon_reg[3] ),
    .QN(_19636_));
 DFFR_X1 \core.keymem.rcon_reg[4]$_DFFE_PN0P_  (.D(_03017_),
    .RN(net87),
    .CK(clknet_leaf_410_clk),
    .Q(\core.keymem.rcon_logic.tmp_rcon[5] ),
    .QN(_19635_));
 DFFR_X1 \core.keymem.rcon_reg[5]$_DFFE_PN0P_  (.D(_03018_),
    .RN(net87),
    .CK(clknet_leaf_411_clk),
    .Q(\core.keymem.rcon_logic.tmp_rcon[6] ),
    .QN(_19634_));
 DFFR_X1 \core.keymem.rcon_reg[6]$_DFFE_PN0P_  (.D(_03019_),
    .RN(net87),
    .CK(clknet_leaf_411_clk),
    .Q(\core.keymem.rcon_logic.tmp_rcon[7] ),
    .QN(_19633_));
 DFFR_X1 \core.keymem.rcon_reg[7]$_DFFE_PN0P_  (.D(_03020_),
    .RN(net87),
    .CK(clknet_leaf_410_clk),
    .Q(\core.keymem.rcon_logic.tmp_rcon[0] ),
    .QN(_19632_));
 DFFR_X2 \core.keymem.ready_reg$_DFFE_PN0P_  (.D(_03021_),
    .RN(net88),
    .CK(clknet_leaf_391_clk),
    .Q(\core.key_ready ),
    .QN(_19631_));
 DFFR_X2 \core.keymem.round_ctr_reg[0]$_DFFE_PN0P_  (.D(_03022_),
    .RN(net88),
    .CK(clknet_leaf_41_clk),
    .Q(\core.keymem.round_ctr_reg[0] ),
    .QN(_22104_));
 DFFR_X2 \core.keymem.round_ctr_reg[1]$_DFFE_PN0P_  (.D(_03023_),
    .RN(net88),
    .CK(clknet_leaf_41_clk),
    .Q(\core.keymem.round_ctr_reg[1] ),
    .QN(_22105_));
 DFFR_X1 \core.keymem.round_ctr_reg[2]$_DFFE_PN0P_  (.D(_03024_),
    .RN(net88),
    .CK(clknet_leaf_44_clk),
    .Q(\core.keymem.round_ctr_reg[2] ),
    .QN(_19630_));
 DFFR_X1 \core.keymem.round_ctr_reg[3]$_DFFE_PN0P_  (.D(_03025_),
    .RN(net88),
    .CK(clknet_leaf_42_clk),
    .Q(\core.keymem.round_ctr_reg[3] ),
    .QN(_00319_));
 DFFS_X2 \core.ready_reg$_DFFE_PN1P_  (.D(_03026_),
    .SN(net84),
    .CK(clknet_leaf_357_clk),
    .Q(\core.ready ),
    .QN(_19629_));
 DFFR_X2 \core.result_valid_reg$_DFFE_PN0P_  (.D(_03027_),
    .RN(net84),
    .CK(clknet_leaf_356_clk),
    .Q(\core.result_valid ),
    .QN(_19628_));
 DFFR_X1 \encdec_reg$_DFFE_PN0P_  (.D(_03028_),
    .RN(net96),
    .CK(clknet_leaf_251_clk),
    .Q(\core.encdec ),
    .QN(_21960_));
 DFFR_X1 \init_reg$_DFF_PN0_  (.D(init_new),
    .RN(net90),
    .CK(clknet_leaf_309_clk),
    .Q(\core.init ),
    .QN(_19627_));
 DFFR_X1 \key_reg[0][0]$_DFFE_PN0P_  (.D(_03029_),
    .RN(net85),
    .CK(clknet_leaf_366_clk),
    .Q(\core.key[224] ),
    .QN(_00121_));
 DFFR_X1 \key_reg[0][10]$_DFFE_PN0P_  (.D(_03030_),
    .RN(net85),
    .CK(clknet_leaf_370_clk),
    .Q(\core.key[234] ),
    .QN(_00135_));
 DFFR_X1 \key_reg[0][11]$_DFFE_PN0P_  (.D(_03031_),
    .RN(net85),
    .CK(clknet_leaf_366_clk),
    .Q(\core.key[235] ),
    .QN(_00137_));
 DFFR_X1 \key_reg[0][12]$_DFFE_PN0P_  (.D(_03032_),
    .RN(net84),
    .CK(clknet_leaf_354_clk),
    .Q(\core.key[236] ),
    .QN(_00139_));
 DFFR_X2 \key_reg[0][13]$_DFFE_PN0P_  (.D(_03033_),
    .RN(net85),
    .CK(clknet_leaf_371_clk),
    .Q(\core.key[237] ),
    .QN(_00141_));
 DFFR_X1 \key_reg[0][14]$_DFFE_PN0P_  (.D(_03034_),
    .RN(net84),
    .CK(clknet_leaf_353_clk),
    .Q(\core.key[238] ),
    .QN(_00142_));
 DFFR_X1 \key_reg[0][15]$_DFFE_PN0P_  (.D(_03035_),
    .RN(net85),
    .CK(clknet_leaf_366_clk),
    .Q(\core.key[239] ),
    .QN(_00143_));
 DFFR_X1 \key_reg[0][16]$_DFFE_PN0P_  (.D(_03036_),
    .RN(net84),
    .CK(clknet_leaf_354_clk),
    .Q(\core.key[240] ),
    .QN(_00145_));
 DFFR_X2 \key_reg[0][17]$_DFFE_PN0P_  (.D(_03037_),
    .RN(net85),
    .CK(clknet_leaf_371_clk),
    .Q(\core.key[241] ),
    .QN(_00146_));
 DFFR_X2 \key_reg[0][18]$_DFFE_PN0P_  (.D(_03038_),
    .RN(net85),
    .CK(clknet_leaf_366_clk),
    .Q(\core.key[242] ),
    .QN(_00147_));
 DFFR_X1 \key_reg[0][19]$_DFFE_PN0P_  (.D(_03039_),
    .RN(net84),
    .CK(clknet_leaf_356_clk),
    .Q(\core.key[243] ),
    .QN(_00149_));
 DFFR_X1 \key_reg[0][1]$_DFFE_PN0P_  (.D(_03040_),
    .RN(net87),
    .CK(clknet_leaf_39_clk),
    .Q(\core.key[225] ),
    .QN(_00122_));
 DFFR_X1 \key_reg[0][20]$_DFFE_PN0P_  (.D(_03041_),
    .RN(net84),
    .CK(clknet_leaf_349_clk),
    .Q(\core.key[244] ),
    .QN(_00151_));
 DFFR_X2 \key_reg[0][21]$_DFFE_PN0P_  (.D(_03042_),
    .RN(net85),
    .CK(clknet_leaf_364_clk),
    .Q(\core.key[245] ),
    .QN(_00153_));
 DFFR_X1 \key_reg[0][22]$_DFFE_PN0P_  (.D(_03043_),
    .RN(net85),
    .CK(clknet_leaf_368_clk),
    .Q(\core.key[246] ),
    .QN(_00154_));
 DFFR_X1 \key_reg[0][23]$_DFFE_PN0P_  (.D(_03044_),
    .RN(net84),
    .CK(clknet_leaf_348_clk),
    .Q(\core.key[247] ),
    .QN(_00155_));
 DFFR_X1 \key_reg[0][24]$_DFFE_PN0P_  (.D(_03045_),
    .RN(net86),
    .CK(clknet_leaf_402_clk),
    .Q(\core.key[248] ),
    .QN(_00157_));
 DFFR_X2 \key_reg[0][25]$_DFFE_PN0P_  (.D(_03046_),
    .RN(net86),
    .CK(clknet_leaf_408_clk),
    .Q(\core.key[249] ),
    .QN(_00159_));
 DFFR_X1 \key_reg[0][26]$_DFFE_PN0P_  (.D(_03047_),
    .RN(net87),
    .CK(clknet_leaf_414_clk),
    .Q(\core.key[250] ),
    .QN(_00161_));
 DFFR_X1 \key_reg[0][27]$_DFFE_PN0P_  (.D(_03048_),
    .RN(net87),
    .CK(clknet_leaf_412_clk),
    .Q(\core.key[251] ),
    .QN(_00163_));
 DFFR_X2 \key_reg[0][28]$_DFFE_PN0P_  (.D(_03049_),
    .RN(net87),
    .CK(clknet_leaf_37_clk),
    .Q(\core.key[252] ),
    .QN(_00165_));
 DFFR_X1 \key_reg[0][29]$_DFFE_PN0P_  (.D(_03050_),
    .RN(net87),
    .CK(clknet_leaf_40_clk),
    .Q(\core.key[253] ),
    .QN(_00167_));
 DFFR_X2 \key_reg[0][2]$_DFFE_PN0P_  (.D(_03051_),
    .RN(net82),
    .CK(clknet_leaf_4_clk),
    .Q(\core.key[226] ),
    .QN(_00123_));
 DFFR_X1 \key_reg[0][30]$_DFFE_PN0P_  (.D(_03052_),
    .RN(net82),
    .CK(clknet_leaf_421_clk),
    .Q(\core.key[254] ),
    .QN(_00169_));
 DFFR_X1 \key_reg[0][31]$_DFFE_PN0P_  (.D(_03053_),
    .RN(net82),
    .CK(clknet_leaf_420_clk),
    .Q(\core.key[255] ),
    .QN(_00171_));
 DFFR_X1 \key_reg[0][3]$_DFFE_PN0P_  (.D(_03054_),
    .RN(net82),
    .CK(clknet_leaf_4_clk),
    .Q(\core.key[227] ),
    .QN(_00125_));
 DFFR_X1 \key_reg[0][4]$_DFFE_PN0P_  (.D(_03055_),
    .RN(net82),
    .CK(clknet_leaf_8_clk),
    .Q(\core.key[228] ),
    .QN(_00127_));
 DFFR_X2 \key_reg[0][5]$_DFFE_PN0P_  (.D(_03056_),
    .RN(net82),
    .CK(clknet_leaf_9_clk),
    .Q(\core.key[229] ),
    .QN(_00129_));
 DFFR_X1 \key_reg[0][6]$_DFFE_PN0P_  (.D(_03057_),
    .RN(net82),
    .CK(clknet_leaf_419_clk),
    .Q(\core.key[230] ),
    .QN(_00130_));
 DFFR_X1 \key_reg[0][7]$_DFFE_PN0P_  (.D(_03058_),
    .RN(net82),
    .CK(clknet_leaf_419_clk),
    .Q(\core.key[231] ),
    .QN(_00131_));
 DFFR_X2 \key_reg[0][8]$_DFFE_PN0P_  (.D(_03059_),
    .RN(net85),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[232] ),
    .QN(_00133_));
 DFFR_X2 \key_reg[0][9]$_DFFE_PN0P_  (.D(_03060_),
    .RN(net89),
    .CK(clknet_leaf_370_clk),
    .Q(\core.key[233] ),
    .QN(_00134_));
 DFFR_X1 \key_reg[1][0]$_DFFE_PN0P_  (.D(_03061_),
    .RN(net84),
    .CK(clknet_leaf_384_clk),
    .Q(\core.key[192] ),
    .QN(_00081_));
 DFFR_X2 \key_reg[1][10]$_DFFE_PN0P_  (.D(_03062_),
    .RN(net85),
    .CK(clknet_leaf_382_clk),
    .Q(\core.key[202] ),
    .QN(_00091_));
 DFFR_X1 \key_reg[1][11]$_DFFE_PN0P_  (.D(_03063_),
    .RN(net85),
    .CK(clknet_leaf_382_clk),
    .Q(\core.key[203] ),
    .QN(_00092_));
 DFFR_X2 \key_reg[1][12]$_DFFE_PN0P_  (.D(_03064_),
    .RN(net89),
    .CK(clknet_leaf_370_clk),
    .Q(\core.key[204] ),
    .QN(_00093_));
 DFFR_X1 \key_reg[1][13]$_DFFE_PN0P_  (.D(_03065_),
    .RN(net85),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[205] ),
    .QN(_00094_));
 DFFR_X1 \key_reg[1][14]$_DFFE_PN0P_  (.D(_03066_),
    .RN(net85),
    .CK(clknet_leaf_369_clk),
    .Q(\core.key[206] ),
    .QN(_00095_));
 DFFR_X1 \key_reg[1][15]$_DFFE_PN0P_  (.D(_03067_),
    .RN(net89),
    .CK(clknet_leaf_370_clk),
    .Q(\core.key[207] ),
    .QN(_00096_));
 DFFR_X2 \key_reg[1][16]$_DFFE_PN0P_  (.D(_03068_),
    .RN(net85),
    .CK(clknet_leaf_369_clk),
    .Q(\core.key[208] ),
    .QN(_00097_));
 DFFR_X1 \key_reg[1][17]$_DFFE_PN0P_  (.D(_03069_),
    .RN(net85),
    .CK(clknet_leaf_369_clk),
    .Q(\core.key[209] ),
    .QN(_00098_));
 DFFR_X2 \key_reg[1][18]$_DFFE_PN0P_  (.D(_03070_),
    .RN(net85),
    .CK(clknet_leaf_382_clk),
    .Q(\core.key[210] ),
    .QN(_00099_));
 DFFR_X1 \key_reg[1][19]$_DFFE_PN0P_  (.D(_03071_),
    .RN(net88),
    .CK(clknet_leaf_42_clk),
    .Q(\core.key[211] ),
    .QN(_00100_));
 DFFR_X2 \key_reg[1][1]$_DFFE_PN0P_  (.D(_03072_),
    .RN(net87),
    .CK(clknet_leaf_40_clk),
    .Q(\core.key[193] ),
    .QN(_00082_));
 DFFR_X1 \key_reg[1][20]$_DFFE_PN0P_  (.D(_03073_),
    .RN(net85),
    .CK(clknet_leaf_368_clk),
    .Q(\core.key[212] ),
    .QN(_00101_));
 DFFR_X1 \key_reg[1][21]$_DFFE_PN0P_  (.D(_03074_),
    .RN(net85),
    .CK(clknet_leaf_370_clk),
    .Q(\core.key[213] ),
    .QN(_00102_));
 DFFR_X1 \key_reg[1][22]$_DFFE_PN0P_  (.D(_03075_),
    .RN(net85),
    .CK(clknet_leaf_369_clk),
    .Q(\core.key[214] ),
    .QN(_00103_));
 DFFR_X1 \key_reg[1][23]$_DFFE_PN0P_  (.D(_03076_),
    .RN(net85),
    .CK(clknet_leaf_369_clk),
    .Q(\core.key[215] ),
    .QN(_00104_));
 DFFR_X2 \key_reg[1][24]$_DFFE_PN0P_  (.D(_03077_),
    .RN(net85),
    .CK(clknet_leaf_370_clk),
    .Q(\core.key[216] ),
    .QN(_00105_));
 DFFR_X2 \key_reg[1][25]$_DFFE_PN0P_  (.D(_03078_),
    .RN(net85),
    .CK(clknet_leaf_384_clk),
    .Q(\core.key[217] ),
    .QN(_00107_));
 DFFR_X2 \key_reg[1][26]$_DFFE_PN0P_  (.D(_03079_),
    .RN(net86),
    .CK(clknet_leaf_41_clk),
    .Q(\core.key[218] ),
    .QN(_00109_));
 DFFR_X2 \key_reg[1][27]$_DFFE_PN0P_  (.D(_03080_),
    .RN(net87),
    .CK(clknet_leaf_41_clk),
    .Q(\core.key[219] ),
    .QN(_00111_));
 DFFR_X2 \key_reg[1][28]$_DFFE_PN0P_  (.D(_03081_),
    .RN(net87),
    .CK(clknet_leaf_36_clk),
    .Q(\core.key[220] ),
    .QN(_00113_));
 DFFR_X2 \key_reg[1][29]$_DFFE_PN0P_  (.D(_03082_),
    .RN(net87),
    .CK(clknet_leaf_40_clk),
    .Q(\core.key[221] ),
    .QN(_00115_));
 DFFR_X2 \key_reg[1][2]$_DFFE_PN0P_  (.D(_03083_),
    .RN(net82),
    .CK(clknet_leaf_9_clk),
    .Q(\core.key[194] ),
    .QN(_00083_));
 DFFR_X2 \key_reg[1][30]$_DFFE_PN0P_  (.D(_03084_),
    .RN(net87),
    .CK(clknet_leaf_37_clk),
    .Q(\core.key[222] ),
    .QN(_00117_));
 DFFR_X2 \key_reg[1][31]$_DFFE_PN0P_  (.D(_03085_),
    .RN(net87),
    .CK(clknet_leaf_37_clk),
    .Q(\core.key[223] ),
    .QN(_00119_));
 DFFR_X2 \key_reg[1][3]$_DFFE_PN0P_  (.D(_03086_),
    .RN(net82),
    .CK(clknet_leaf_35_clk),
    .Q(\core.key[195] ),
    .QN(_00084_));
 DFFR_X1 \key_reg[1][4]$_DFFE_PN0P_  (.D(_03087_),
    .RN(net82),
    .CK(clknet_leaf_9_clk),
    .Q(\core.key[196] ),
    .QN(_00085_));
 DFFR_X2 \key_reg[1][5]$_DFFE_PN0P_  (.D(_03088_),
    .RN(net82),
    .CK(clknet_leaf_36_clk),
    .Q(\core.key[197] ),
    .QN(_00086_));
 DFFR_X1 \key_reg[1][6]$_DFFE_PN0P_  (.D(_03089_),
    .RN(net82),
    .CK(clknet_leaf_9_clk),
    .Q(\core.key[198] ),
    .QN(_00087_));
 DFFR_X1 \key_reg[1][7]$_DFFE_PN0P_  (.D(_03090_),
    .RN(net82),
    .CK(clknet_leaf_9_clk),
    .Q(\core.key[199] ),
    .QN(_00088_));
 DFFR_X1 \key_reg[1][8]$_DFFE_PN0P_  (.D(_03091_),
    .RN(net88),
    .CK(clknet_leaf_389_clk),
    .Q(\core.key[200] ),
    .QN(_00089_));
 DFFR_X1 \key_reg[1][9]$_DFFE_PN0P_  (.D(_03092_),
    .RN(net86),
    .CK(clknet_leaf_393_clk),
    .Q(\core.key[201] ),
    .QN(_00090_));
 DFFR_X1 \key_reg[2][0]$_DFFE_PN0P_  (.D(_03093_),
    .RN(net85),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[160] ),
    .QN(_00041_));
 DFFR_X1 \key_reg[2][10]$_DFFE_PN0P_  (.D(_03094_),
    .RN(net85),
    .CK(clknet_leaf_382_clk),
    .Q(\core.key[170] ),
    .QN(_00051_));
 DFFR_X2 \key_reg[2][11]$_DFFE_PN0P_  (.D(_03095_),
    .RN(net85),
    .CK(clknet_leaf_382_clk),
    .Q(\core.key[171] ),
    .QN(_00052_));
 DFFR_X1 \key_reg[2][12]$_DFFE_PN0P_  (.D(_03096_),
    .RN(net84),
    .CK(clknet_leaf_384_clk),
    .Q(\core.key[172] ),
    .QN(_00053_));
 DFFR_X2 \key_reg[2][13]$_DFFE_PN0P_  (.D(_03097_),
    .RN(net85),
    .CK(clknet_leaf_43_clk),
    .Q(\core.key[173] ),
    .QN(_00054_));
 DFFR_X2 \key_reg[2][14]$_DFFE_PN0P_  (.D(_03098_),
    .RN(net89),
    .CK(clknet_leaf_380_clk),
    .Q(\core.key[174] ),
    .QN(_00055_));
 DFFR_X2 \key_reg[2][15]$_DFFE_PN0P_  (.D(_03099_),
    .RN(net85),
    .CK(clknet_leaf_385_clk),
    .Q(\core.key[175] ),
    .QN(_00056_));
 DFFR_X1 \key_reg[2][16]$_DFFE_PN0P_  (.D(_03100_),
    .RN(net85),
    .CK(clknet_leaf_385_clk),
    .Q(\core.key[176] ),
    .QN(_00057_));
 DFFR_X2 \key_reg[2][17]$_DFFE_PN0P_  (.D(_03101_),
    .RN(net85),
    .CK(clknet_leaf_381_clk),
    .Q(\core.key[177] ),
    .QN(_00058_));
 DFFR_X2 \key_reg[2][18]$_DFFE_PN0P_  (.D(_03102_),
    .RN(net88),
    .CK(clknet_leaf_43_clk),
    .Q(\core.key[178] ),
    .QN(_00059_));
 DFFR_X1 \key_reg[2][19]$_DFFE_PN0P_  (.D(_03103_),
    .RN(net87),
    .CK(clknet_leaf_37_clk),
    .Q(\core.key[179] ),
    .QN(_00060_));
 DFFR_X1 \key_reg[2][1]$_DFFE_PN0P_  (.D(_03104_),
    .RN(net87),
    .CK(clknet_leaf_37_clk),
    .Q(\core.key[161] ),
    .QN(_00042_));
 DFFR_X1 \key_reg[2][20]$_DFFE_PN0P_  (.D(_03105_),
    .RN(net84),
    .CK(clknet_leaf_384_clk),
    .Q(\core.key[180] ),
    .QN(_00061_));
 DFFR_X1 \key_reg[2][21]$_DFFE_PN0P_  (.D(_03106_),
    .RN(net85),
    .CK(clknet_leaf_384_clk),
    .Q(\core.key[181] ),
    .QN(_00062_));
 DFFR_X2 \key_reg[2][22]$_DFFE_PN0P_  (.D(_03107_),
    .RN(net85),
    .CK(clknet_leaf_381_clk),
    .Q(\core.key[182] ),
    .QN(_00063_));
 DFFR_X2 \key_reg[2][23]$_DFFE_PN0P_  (.D(_03108_),
    .RN(net85),
    .CK(clknet_leaf_381_clk),
    .Q(\core.key[183] ),
    .QN(_00064_));
 DFFR_X2 \key_reg[2][24]$_DFFE_PN0P_  (.D(_03109_),
    .RN(net88),
    .CK(clknet_leaf_43_clk),
    .Q(\core.key[184] ),
    .QN(_00065_));
 DFFR_X2 \key_reg[2][25]$_DFFE_PN0P_  (.D(_03110_),
    .RN(net88),
    .CK(clknet_leaf_390_clk),
    .Q(\core.key[185] ),
    .QN(_00067_));
 DFFR_X1 \key_reg[2][26]$_DFFE_PN0P_  (.D(_03111_),
    .RN(net87),
    .CK(clknet_leaf_40_clk),
    .Q(\core.key[186] ),
    .QN(_00069_));
 DFFR_X1 \key_reg[2][27]$_DFFE_PN0P_  (.D(_03112_),
    .RN(net87),
    .CK(clknet_leaf_40_clk),
    .Q(\core.key[187] ),
    .QN(_00071_));
 DFFR_X2 \key_reg[2][28]$_DFFE_PN0P_  (.D(_03113_),
    .RN(net82),
    .CK(clknet_leaf_11_clk),
    .Q(\core.key[188] ),
    .QN(_00073_));
 DFFR_X2 \key_reg[2][29]$_DFFE_PN0P_  (.D(_03114_),
    .RN(net82),
    .CK(clknet_leaf_11_clk),
    .Q(\core.key[189] ),
    .QN(_00075_));
 DFFR_X1 \key_reg[2][2]$_DFFE_PN0P_  (.D(_03115_),
    .RN(net82),
    .CK(clknet_leaf_2_clk),
    .Q(\core.key[162] ),
    .QN(_00043_));
 DFFR_X2 \key_reg[2][30]$_DFFE_PN0P_  (.D(_03116_),
    .RN(net82),
    .CK(clknet_leaf_2_clk),
    .Q(\core.key[190] ),
    .QN(_00077_));
 DFFR_X1 \key_reg[2][31]$_DFFE_PN0P_  (.D(_03117_),
    .RN(net82),
    .CK(clknet_leaf_10_clk),
    .Q(\core.key[191] ),
    .QN(_00079_));
 DFFR_X1 \key_reg[2][3]$_DFFE_PN0P_  (.D(_03118_),
    .RN(net82),
    .CK(clknet_leaf_3_clk),
    .Q(\core.key[163] ),
    .QN(_00044_));
 DFFR_X1 \key_reg[2][4]$_DFFE_PN0P_  (.D(_03119_),
    .RN(net82),
    .CK(clknet_leaf_11_clk),
    .Q(\core.key[164] ),
    .QN(_00045_));
 DFFR_X1 \key_reg[2][5]$_DFFE_PN0P_  (.D(_03120_),
    .RN(net82),
    .CK(clknet_leaf_12_clk),
    .Q(\core.key[165] ),
    .QN(_00046_));
 DFFR_X1 \key_reg[2][6]$_DFFE_PN0P_  (.D(_03121_),
    .RN(net82),
    .CK(clknet_leaf_4_clk),
    .Q(\core.key[166] ),
    .QN(_00047_));
 DFFR_X2 \key_reg[2][7]$_DFFE_PN0P_  (.D(_03122_),
    .RN(net82),
    .CK(clknet_leaf_10_clk),
    .Q(\core.key[167] ),
    .QN(_00048_));
 DFFR_X2 \key_reg[2][8]$_DFFE_PN0P_  (.D(_03123_),
    .RN(net87),
    .CK(clknet_leaf_36_clk),
    .Q(\core.key[168] ),
    .QN(_00049_));
 DFFR_X1 \key_reg[2][9]$_DFFE_PN0P_  (.D(_03124_),
    .RN(net87),
    .CK(clknet_leaf_39_clk),
    .Q(\core.key[169] ),
    .QN(_00050_));
 DFFR_X1 \key_reg[3][0]$_DFFE_PN0P_  (.D(_03125_),
    .RN(net85),
    .CK(clknet_leaf_384_clk),
    .Q(\core.key[128] ),
    .QN(_00327_));
 DFFR_X1 \key_reg[3][10]$_DFFE_PN0P_  (.D(_03126_),
    .RN(net85),
    .CK(clknet_leaf_382_clk),
    .Q(\core.key[138] ),
    .QN(_00405_));
 DFFR_X2 \key_reg[3][11]$_DFFE_PN0P_  (.D(_03127_),
    .RN(net85),
    .CK(clknet_leaf_382_clk),
    .Q(\core.key[139] ),
    .QN(_00406_));
 DFFR_X2 \key_reg[3][12]$_DFFE_PN0P_  (.D(_03128_),
    .RN(net89),
    .CK(clknet_leaf_380_clk),
    .Q(\core.key[140] ),
    .QN(_00407_));
 DFFR_X1 \key_reg[3][13]$_DFFE_PN0P_  (.D(_03129_),
    .RN(net88),
    .CK(clknet_leaf_390_clk),
    .Q(\core.key[141] ),
    .QN(_00408_));
 DFFR_X2 \key_reg[3][14]$_DFFE_PN0P_  (.D(_03130_),
    .RN(net89),
    .CK(clknet_leaf_375_clk),
    .Q(\core.key[142] ),
    .QN(_00409_));
 DFFR_X1 \key_reg[3][15]$_DFFE_PN0P_  (.D(_03131_),
    .RN(net85),
    .CK(clknet_leaf_369_clk),
    .Q(\core.key[143] ),
    .QN(_00410_));
 DFFR_X2 \key_reg[3][16]$_DFFE_PN0P_  (.D(_03132_),
    .RN(net89),
    .CK(clknet_leaf_375_clk),
    .Q(\core.key[144] ),
    .QN(_00411_));
 DFFR_X2 \key_reg[3][17]$_DFFE_PN0P_  (.D(_03133_),
    .RN(net89),
    .CK(clknet_leaf_369_clk),
    .Q(\core.key[145] ),
    .QN(_00434_));
 DFFR_X2 \key_reg[3][18]$_DFFE_PN0P_  (.D(_03134_),
    .RN(net88),
    .CK(clknet_leaf_390_clk),
    .Q(\core.key[146] ),
    .QN(_00435_));
 DFFR_X1 \key_reg[3][19]$_DFFE_PN0P_  (.D(_03135_),
    .RN(net86),
    .CK(clknet_leaf_391_clk),
    .Q(\core.key[147] ),
    .QN(_00436_));
 DFFR_X1 \key_reg[3][1]$_DFFE_PN0P_  (.D(_03136_),
    .RN(net87),
    .CK(clknet_leaf_39_clk),
    .Q(\core.key[129] ),
    .QN(_00371_));
 DFFR_X2 \key_reg[3][20]$_DFFE_PN0P_  (.D(_03137_),
    .RN(net85),
    .CK(clknet_leaf_384_clk),
    .Q(\core.key[148] ),
    .QN(_00437_));
 DFFR_X2 \key_reg[3][21]$_DFFE_PN0P_  (.D(_03138_),
    .RN(net85),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[149] ),
    .QN(_00438_));
 DFFR_X1 \key_reg[3][22]$_DFFE_PN0P_  (.D(_03139_),
    .RN(net85),
    .CK(clknet_leaf_380_clk),
    .Q(\core.key[150] ),
    .QN(_00015_));
 DFFR_X1 \key_reg[3][23]$_DFFE_PN0P_  (.D(_03140_),
    .RN(net86),
    .CK(clknet_leaf_403_clk),
    .Q(\core.key[151] ),
    .QN(_00016_));
 DFFR_X2 \key_reg[3][24]$_DFFE_PN0P_  (.D(_03141_),
    .RN(net88),
    .CK(clknet_leaf_43_clk),
    .Q(\core.key[152] ),
    .QN(_00017_));
 DFFR_X2 \key_reg[3][25]$_DFFE_PN0P_  (.D(_03142_),
    .RN(net88),
    .CK(clknet_leaf_390_clk),
    .Q(\core.key[153] ),
    .QN(_00020_));
 DFFR_X1 \key_reg[3][26]$_DFFE_PN0P_  (.D(_03143_),
    .RN(net87),
    .CK(clknet_leaf_413_clk),
    .Q(\core.key[154] ),
    .QN(_00023_));
 DFFR_X2 \key_reg[3][27]$_DFFE_PN0P_  (.D(_03144_),
    .RN(net87),
    .CK(clknet_leaf_39_clk),
    .Q(\core.key[155] ),
    .QN(_00026_));
 DFFR_X1 \key_reg[3][28]$_DFFE_PN0P_  (.D(_03145_),
    .RN(net82),
    .CK(clknet_leaf_36_clk),
    .Q(\core.key[156] ),
    .QN(_00029_));
 DFFR_X2 \key_reg[3][29]$_DFFE_PN0P_  (.D(_03146_),
    .RN(net87),
    .CK(clknet_leaf_37_clk),
    .Q(\core.key[157] ),
    .QN(_00032_));
 DFFR_X2 \key_reg[3][2]$_DFFE_PN0P_  (.D(_03147_),
    .RN(net86),
    .CK(clknet_leaf_41_clk),
    .Q(\core.key[130] ),
    .QN(_00373_));
 DFFR_X2 \key_reg[3][30]$_DFFE_PN0P_  (.D(_03148_),
    .RN(net87),
    .CK(clknet_leaf_40_clk),
    .Q(\core.key[158] ),
    .QN(_00035_));
 DFFR_X2 \key_reg[3][31]$_DFFE_PN0P_  (.D(_03149_),
    .RN(net87),
    .CK(clknet_leaf_37_clk),
    .Q(\core.key[159] ),
    .QN(_00038_));
 DFFR_X2 \key_reg[3][3]$_DFFE_PN0P_  (.D(_03150_),
    .RN(net87),
    .CK(clknet_leaf_38_clk),
    .Q(\core.key[131] ),
    .QN(_00374_));
 DFFR_X2 \key_reg[3][4]$_DFFE_PN0P_  (.D(_03151_),
    .RN(net82),
    .CK(clknet_leaf_35_clk),
    .Q(\core.key[132] ),
    .QN(_00375_));
 DFFR_X1 \key_reg[3][5]$_DFFE_PN0P_  (.D(_03152_),
    .RN(net82),
    .CK(clknet_leaf_9_clk),
    .Q(\core.key[133] ),
    .QN(_00376_));
 DFFR_X2 \key_reg[3][6]$_DFFE_PN0P_  (.D(_03153_),
    .RN(net87),
    .CK(clknet_leaf_36_clk),
    .Q(\core.key[134] ),
    .QN(_00378_));
 DFFR_X2 \key_reg[3][7]$_DFFE_PN0P_  (.D(_03154_),
    .RN(net88),
    .CK(clknet_leaf_391_clk),
    .Q(\core.key[135] ),
    .QN(_00380_));
 DFFR_X1 \key_reg[3][8]$_DFFE_PN0P_  (.D(_03155_),
    .RN(net89),
    .CK(clknet_leaf_380_clk),
    .Q(\core.key[136] ),
    .QN(_00381_));
 DFFR_X2 \key_reg[3][9]$_DFFE_PN0P_  (.D(_03156_),
    .RN(net85),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[137] ),
    .QN(_00404_));
 DFFR_X1 \key_reg[4][0]$_DFFE_PN0P_  (.D(_03157_),
    .RN(net84),
    .CK(clknet_leaf_385_clk),
    .Q(\core.key[96] ),
    .QN(_19626_));
 DFFR_X1 \key_reg[4][10]$_DFFE_PN0P_  (.D(_03158_),
    .RN(net88),
    .CK(clknet_leaf_389_clk),
    .Q(\core.key[106] ),
    .QN(_19625_));
 DFFR_X1 \key_reg[4][11]$_DFFE_PN0P_  (.D(_03159_),
    .RN(net85),
    .CK(clknet_leaf_368_clk),
    .Q(\core.key[107] ),
    .QN(_19624_));
 DFFR_X1 \key_reg[4][12]$_DFFE_PN0P_  (.D(_03160_),
    .RN(net84),
    .CK(clknet_leaf_355_clk),
    .Q(\core.key[108] ),
    .QN(_19623_));
 DFFR_X1 \key_reg[4][13]$_DFFE_PN0P_  (.D(_03161_),
    .RN(net88),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[109] ),
    .QN(_19622_));
 DFFR_X1 \key_reg[4][14]$_DFFE_PN0P_  (.D(_03162_),
    .RN(net84),
    .CK(clknet_leaf_355_clk),
    .Q(\core.key[110] ),
    .QN(_19621_));
 DFFR_X1 \key_reg[4][15]$_DFFE_PN0P_  (.D(_03163_),
    .RN(net85),
    .CK(clknet_leaf_366_clk),
    .Q(\core.key[111] ),
    .QN(_19620_));
 DFFR_X1 \key_reg[4][16]$_DFFE_PN0P_  (.D(_03164_),
    .RN(net84),
    .CK(clknet_leaf_354_clk),
    .Q(\core.key[112] ),
    .QN(_19619_));
 DFFR_X1 \key_reg[4][17]$_DFFE_PN0P_  (.D(_03165_),
    .RN(net85),
    .CK(clknet_leaf_370_clk),
    .Q(\core.key[113] ),
    .QN(_19618_));
 DFFR_X1 \key_reg[4][18]$_DFFE_PN0P_  (.D(_03166_),
    .RN(net88),
    .CK(clknet_leaf_389_clk),
    .Q(\core.key[114] ),
    .QN(_19617_));
 DFFR_X1 \key_reg[4][19]$_DFFE_PN0P_  (.D(_03167_),
    .RN(net84),
    .CK(clknet_leaf_351_clk),
    .Q(\core.key[115] ),
    .QN(_19616_));
 DFFR_X1 \key_reg[4][1]$_DFFE_PN0P_  (.D(_03168_),
    .RN(net87),
    .CK(clknet_leaf_394_clk),
    .Q(\core.key[97] ),
    .QN(_19615_));
 DFFR_X1 \key_reg[4][20]$_DFFE_PN0P_  (.D(_03169_),
    .RN(net86),
    .CK(clknet_leaf_348_clk),
    .Q(\core.key[116] ),
    .QN(_19614_));
 DFFR_X1 \key_reg[4][21]$_DFFE_PN0P_  (.D(_03170_),
    .RN(net86),
    .CK(clknet_leaf_348_clk),
    .Q(\core.key[117] ),
    .QN(_19613_));
 DFFR_X1 \key_reg[4][22]$_DFFE_PN0P_  (.D(_03171_),
    .RN(net86),
    .CK(clknet_leaf_348_clk),
    .Q(\core.key[118] ),
    .QN(_19612_));
 DFFR_X1 \key_reg[4][23]$_DFFE_PN0P_  (.D(_03172_),
    .RN(net86),
    .CK(clknet_leaf_348_clk),
    .Q(\core.key[119] ),
    .QN(_19611_));
 DFFR_X1 \key_reg[4][24]$_DFFE_PN0P_  (.D(_03173_),
    .RN(net86),
    .CK(clknet_leaf_402_clk),
    .Q(\core.key[120] ),
    .QN(_00158_));
 DFFR_X1 \key_reg[4][25]$_DFFE_PN0P_  (.D(_03174_),
    .RN(net86),
    .CK(clknet_leaf_408_clk),
    .Q(\core.key[121] ),
    .QN(_00160_));
 DFFR_X1 \key_reg[4][26]$_DFFE_PN0P_  (.D(_03175_),
    .RN(net87),
    .CK(clknet_leaf_414_clk),
    .Q(\core.key[122] ),
    .QN(_00162_));
 DFFR_X1 \key_reg[4][27]$_DFFE_PN0P_  (.D(_03176_),
    .RN(net87),
    .CK(clknet_leaf_412_clk),
    .Q(\core.key[123] ),
    .QN(_00164_));
 DFFR_X1 \key_reg[4][28]$_DFFE_PN0P_  (.D(_03177_),
    .RN(net82),
    .CK(clknet_leaf_12_clk),
    .Q(\core.key[124] ),
    .QN(_00166_));
 DFFR_X1 \key_reg[4][29]$_DFFE_PN0P_  (.D(_03178_),
    .RN(net82),
    .CK(clknet_leaf_2_clk),
    .Q(\core.key[125] ),
    .QN(_00168_));
 DFFR_X1 \key_reg[4][2]$_DFFE_PN0P_  (.D(_03179_),
    .RN(net82),
    .CK(clknet_leaf_2_clk),
    .Q(\core.key[98] ),
    .QN(_19610_));
 DFFR_X1 \key_reg[4][30]$_DFFE_PN0P_  (.D(_03180_),
    .RN(net82),
    .CK(clknet_leaf_0_clk),
    .Q(\core.key[126] ),
    .QN(_00170_));
 DFFR_X1 \key_reg[4][31]$_DFFE_PN0P_  (.D(_03181_),
    .RN(net82),
    .CK(clknet_leaf_424_clk),
    .Q(\core.key[127] ),
    .QN(_00172_));
 DFFR_X1 \key_reg[4][3]$_DFFE_PN0P_  (.D(_03182_),
    .RN(net82),
    .CK(clknet_leaf_425_clk),
    .Q(\core.key[99] ),
    .QN(_19609_));
 DFFR_X1 \key_reg[4][4]$_DFFE_PN0P_  (.D(_03183_),
    .RN(net82),
    .CK(clknet_leaf_12_clk),
    .Q(\core.key[100] ),
    .QN(_19608_));
 DFFR_X1 \key_reg[4][5]$_DFFE_PN0P_  (.D(_03184_),
    .RN(net82),
    .CK(clknet_leaf_1_clk),
    .Q(\core.key[101] ),
    .QN(_19607_));
 DFFR_X1 \key_reg[4][6]$_DFFE_PN0P_  (.D(_03185_),
    .RN(net82),
    .CK(clknet_leaf_425_clk),
    .Q(\core.key[102] ),
    .QN(_19606_));
 DFFR_X1 \key_reg[4][7]$_DFFE_PN0P_  (.D(_03186_),
    .RN(net82),
    .CK(clknet_leaf_424_clk),
    .Q(\core.key[103] ),
    .QN(_19605_));
 DFFR_X1 \key_reg[4][8]$_DFFE_PN0P_  (.D(_03187_),
    .RN(net86),
    .CK(clknet_leaf_398_clk),
    .Q(\core.key[104] ),
    .QN(_19604_));
 DFFR_X1 \key_reg[4][9]$_DFFE_PN0P_  (.D(_03188_),
    .RN(net84),
    .CK(clknet_leaf_366_clk),
    .Q(\core.key[105] ),
    .QN(_19603_));
 DFFR_X1 \key_reg[5][0]$_DFFE_PN0P_  (.D(_03189_),
    .RN(net84),
    .CK(clknet_leaf_385_clk),
    .Q(\core.key[64] ),
    .QN(_19602_));
 DFFR_X1 \key_reg[5][10]$_DFFE_PN0P_  (.D(_03190_),
    .RN(net88),
    .CK(clknet_leaf_389_clk),
    .Q(\core.key[74] ),
    .QN(_19601_));
 DFFR_X1 \key_reg[5][11]$_DFFE_PN0P_  (.D(_03191_),
    .RN(net88),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[75] ),
    .QN(_19600_));
 DFFR_X1 \key_reg[5][12]$_DFFE_PN0P_  (.D(_03192_),
    .RN(net85),
    .CK(clknet_leaf_367_clk),
    .Q(\core.key[76] ),
    .QN(_19599_));
 DFFR_X1 \key_reg[5][13]$_DFFE_PN0P_  (.D(_03193_),
    .RN(net88),
    .CK(clknet_leaf_390_clk),
    .Q(\core.key[77] ),
    .QN(_19598_));
 DFFR_X1 \key_reg[5][14]$_DFFE_PN0P_  (.D(_03194_),
    .RN(net85),
    .CK(clknet_leaf_368_clk),
    .Q(\core.key[78] ),
    .QN(_19597_));
 DFFR_X1 \key_reg[5][15]$_DFFE_PN0P_  (.D(_03195_),
    .RN(net85),
    .CK(clknet_leaf_368_clk),
    .Q(\core.key[79] ),
    .QN(_19596_));
 DFFR_X1 \key_reg[5][16]$_DFFE_PN0P_  (.D(_03196_),
    .RN(net84),
    .CK(clknet_leaf_367_clk),
    .Q(\core.key[80] ),
    .QN(_19595_));
 DFFR_X1 \key_reg[5][17]$_DFFE_PN0P_  (.D(_03197_),
    .RN(net85),
    .CK(clknet_leaf_368_clk),
    .Q(\core.key[81] ),
    .QN(_19594_));
 DFFR_X1 \key_reg[5][18]$_DFFE_PN0P_  (.D(_03198_),
    .RN(net88),
    .CK(clknet_leaf_389_clk),
    .Q(\core.key[82] ),
    .QN(_19593_));
 DFFR_X1 \key_reg[5][19]$_DFFE_PN0P_  (.D(_03199_),
    .RN(net86),
    .CK(clknet_leaf_395_clk),
    .Q(\core.key[83] ),
    .QN(_19592_));
 DFFR_X1 \key_reg[5][1]$_DFFE_PN0P_  (.D(_03200_),
    .RN(net87),
    .CK(clknet_leaf_417_clk),
    .Q(\core.key[65] ),
    .QN(_19591_));
 DFFR_X1 \key_reg[5][20]$_DFFE_PN0P_  (.D(_03201_),
    .RN(net86),
    .CK(clknet_leaf_348_clk),
    .Q(\core.key[84] ),
    .QN(_19590_));
 DFFR_X1 \key_reg[5][21]$_DFFE_PN0P_  (.D(_03202_),
    .RN(net84),
    .CK(clknet_leaf_353_clk),
    .Q(\core.key[85] ),
    .QN(_19589_));
 DFFR_X1 \key_reg[5][22]$_DFFE_PN0P_  (.D(_03203_),
    .RN(net84),
    .CK(clknet_leaf_350_clk),
    .Q(\core.key[86] ),
    .QN(_19588_));
 DFFR_X1 \key_reg[5][23]$_DFFE_PN0P_  (.D(_03204_),
    .RN(net86),
    .CK(clknet_leaf_347_clk),
    .Q(\core.key[87] ),
    .QN(_19587_));
 DFFR_X1 \key_reg[5][24]$_DFFE_PN0P_  (.D(_03205_),
    .RN(net86),
    .CK(clknet_leaf_408_clk),
    .Q(\core.key[88] ),
    .QN(_00106_));
 DFFR_X1 \key_reg[5][25]$_DFFE_PN0P_  (.D(_03206_),
    .RN(net86),
    .CK(clknet_leaf_408_clk),
    .Q(\core.key[89] ),
    .QN(_00108_));
 DFFR_X1 \key_reg[5][26]$_DFFE_PN0P_  (.D(_03207_),
    .RN(net87),
    .CK(clknet_leaf_413_clk),
    .Q(\core.key[90] ),
    .QN(_00110_));
 DFFR_X1 \key_reg[5][27]$_DFFE_PN0P_  (.D(_03208_),
    .RN(net87),
    .CK(clknet_leaf_416_clk),
    .Q(\core.key[91] ),
    .QN(_00112_));
 DFFR_X1 \key_reg[5][28]$_DFFE_PN0P_  (.D(_03209_),
    .RN(net82),
    .CK(clknet_leaf_11_clk),
    .Q(\core.key[92] ),
    .QN(_00114_));
 DFFR_X1 \key_reg[5][29]$_DFFE_PN0P_  (.D(_03210_),
    .RN(net82),
    .CK(clknet_leaf_1_clk),
    .Q(\core.key[93] ),
    .QN(_00116_));
 DFFR_X1 \key_reg[5][2]$_DFFE_PN0P_  (.D(_03211_),
    .RN(net82),
    .CK(clknet_leaf_2_clk),
    .Q(\core.key[66] ),
    .QN(_19586_));
 DFFR_X1 \key_reg[5][30]$_DFFE_PN0P_  (.D(_03212_),
    .RN(net82),
    .CK(clknet_leaf_1_clk),
    .Q(\core.key[94] ),
    .QN(_00118_));
 DFFR_X1 \key_reg[5][31]$_DFFE_PN0P_  (.D(_03213_),
    .RN(net82),
    .CK(clknet_leaf_3_clk),
    .Q(\core.key[95] ),
    .QN(_00120_));
 DFFR_X1 \key_reg[5][3]$_DFFE_PN0P_  (.D(_03214_),
    .RN(net82),
    .CK(clknet_leaf_3_clk),
    .Q(\core.key[67] ),
    .QN(_19585_));
 DFFR_X1 \key_reg[5][4]$_DFFE_PN0P_  (.D(_03215_),
    .RN(net82),
    .CK(clknet_leaf_8_clk),
    .Q(\core.key[68] ),
    .QN(_19584_));
 DFFR_X1 \key_reg[5][5]$_DFFE_PN0P_  (.D(_03216_),
    .RN(net82),
    .CK(clknet_leaf_12_clk),
    .Q(\core.key[69] ),
    .QN(_19583_));
 DFFR_X1 \key_reg[5][6]$_DFFE_PN0P_  (.D(_03217_),
    .RN(net82),
    .CK(clknet_leaf_3_clk),
    .Q(\core.key[70] ),
    .QN(_19582_));
 DFFR_X1 \key_reg[5][7]$_DFFE_PN0P_  (.D(_03218_),
    .RN(net82),
    .CK(clknet_leaf_4_clk),
    .Q(\core.key[71] ),
    .QN(_19581_));
 DFFR_X1 \key_reg[5][8]$_DFFE_PN0P_  (.D(_03219_),
    .RN(net86),
    .CK(clknet_leaf_397_clk),
    .Q(\core.key[72] ),
    .QN(_19580_));
 DFFR_X1 \key_reg[5][9]$_DFFE_PN0P_  (.D(_03220_),
    .RN(net86),
    .CK(clknet_leaf_391_clk),
    .Q(\core.key[73] ),
    .QN(_19579_));
 DFFR_X1 \key_reg[6][0]$_DFFE_PN0P_  (.D(_03221_),
    .RN(net88),
    .CK(clknet_leaf_384_clk),
    .Q(\core.key[32] ),
    .QN(_19578_));
 DFFR_X1 \key_reg[6][10]$_DFFE_PN0P_  (.D(_03222_),
    .RN(net88),
    .CK(clknet_leaf_390_clk),
    .Q(\core.key[42] ),
    .QN(_19577_));
 DFFR_X1 \key_reg[6][11]$_DFFE_PN0P_  (.D(_03223_),
    .RN(net88),
    .CK(clknet_leaf_389_clk),
    .Q(\core.key[43] ),
    .QN(_19576_));
 DFFR_X1 \key_reg[6][12]$_DFFE_PN0P_  (.D(_03224_),
    .RN(net86),
    .CK(clknet_leaf_400_clk),
    .Q(\core.key[44] ),
    .QN(_19575_));
 DFFR_X1 \key_reg[6][13]$_DFFE_PN0P_  (.D(_03225_),
    .RN(net88),
    .CK(clknet_leaf_391_clk),
    .Q(\core.key[45] ),
    .QN(_19574_));
 DFFR_X1 \key_reg[6][14]$_DFFE_PN0P_  (.D(_03226_),
    .RN(net88),
    .CK(clknet_leaf_400_clk),
    .Q(\core.key[46] ),
    .QN(_19573_));
 DFFR_X1 \key_reg[6][15]$_DFFE_PN0P_  (.D(_03227_),
    .RN(net84),
    .CK(clknet_leaf_385_clk),
    .Q(\core.key[47] ),
    .QN(_19572_));
 DFFR_X1 \key_reg[6][16]$_DFFE_PN0P_  (.D(_03228_),
    .RN(net88),
    .CK(clknet_leaf_399_clk),
    .Q(\core.key[48] ),
    .QN(_19571_));
 DFFR_X1 \key_reg[6][17]$_DFFE_PN0P_  (.D(_03229_),
    .RN(net88),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[49] ),
    .QN(_19570_));
 DFFR_X1 \key_reg[6][18]$_DFFE_PN0P_  (.D(_03230_),
    .RN(net86),
    .CK(clknet_leaf_392_clk),
    .Q(\core.key[50] ),
    .QN(_19569_));
 DFFR_X1 \key_reg[6][19]$_DFFE_PN0P_  (.D(_03231_),
    .RN(net87),
    .CK(clknet_leaf_393_clk),
    .Q(\core.key[51] ),
    .QN(_19568_));
 DFFR_X1 \key_reg[6][1]$_DFFE_PN0P_  (.D(_03232_),
    .RN(net87),
    .CK(clknet_leaf_394_clk),
    .Q(\core.key[33] ),
    .QN(_19567_));
 DFFR_X1 \key_reg[6][20]$_DFFE_PN0P_  (.D(_03233_),
    .RN(net86),
    .CK(clknet_leaf_403_clk),
    .Q(\core.key[52] ),
    .QN(_19566_));
 DFFR_X1 \key_reg[6][21]$_DFFE_PN0P_  (.D(_03234_),
    .RN(net86),
    .CK(clknet_leaf_403_clk),
    .Q(\core.key[53] ),
    .QN(_19565_));
 DFFR_X1 \key_reg[6][22]$_DFFE_PN0P_  (.D(_03235_),
    .RN(net86),
    .CK(clknet_leaf_403_clk),
    .Q(\core.key[54] ),
    .QN(_19564_));
 DFFR_X1 \key_reg[6][23]$_DFFE_PN0P_  (.D(_03236_),
    .RN(net86),
    .CK(clknet_leaf_404_clk),
    .Q(\core.key[55] ),
    .QN(_19563_));
 DFFR_X1 \key_reg[6][24]$_DFFE_PN0P_  (.D(_03237_),
    .RN(net87),
    .CK(clknet_leaf_414_clk),
    .Q(\core.key[56] ),
    .QN(_00066_));
 DFFR_X1 \key_reg[6][25]$_DFFE_PN0P_  (.D(_03238_),
    .RN(net86),
    .CK(clknet_leaf_409_clk),
    .Q(\core.key[57] ),
    .QN(_00068_));
 DFFR_X1 \key_reg[6][26]$_DFFE_PN0P_  (.D(_03239_),
    .RN(net87),
    .CK(clknet_leaf_413_clk),
    .Q(\core.key[58] ),
    .QN(_00070_));
 DFFR_X1 \key_reg[6][27]$_DFFE_PN0P_  (.D(_03240_),
    .RN(net87),
    .CK(clknet_leaf_412_clk),
    .Q(\core.key[59] ),
    .QN(_00072_));
 DFFR_X1 \key_reg[6][28]$_DFFE_PN0P_  (.D(_03241_),
    .RN(net82),
    .CK(clknet_leaf_11_clk),
    .Q(\core.key[60] ),
    .QN(_00074_));
 DFFR_X1 \key_reg[6][29]$_DFFE_PN0P_  (.D(_03242_),
    .RN(net82),
    .CK(clknet_leaf_1_clk),
    .Q(\core.key[61] ),
    .QN(_00076_));
 DFFR_X1 \key_reg[6][2]$_DFFE_PN0P_  (.D(_03243_),
    .RN(net82),
    .CK(clknet_leaf_2_clk),
    .Q(\core.key[34] ),
    .QN(_19562_));
 DFFR_X1 \key_reg[6][30]$_DFFE_PN0P_  (.D(_03244_),
    .RN(net82),
    .CK(clknet_leaf_2_clk),
    .Q(\core.key[62] ),
    .QN(_00078_));
 DFFR_X1 \key_reg[6][31]$_DFFE_PN0P_  (.D(_03245_),
    .RN(net82),
    .CK(clknet_leaf_0_clk),
    .Q(\core.key[63] ),
    .QN(_00080_));
 DFFR_X1 \key_reg[6][3]$_DFFE_PN0P_  (.D(_03246_),
    .RN(net82),
    .CK(clknet_leaf_0_clk),
    .Q(\core.key[35] ),
    .QN(_19561_));
 DFFR_X1 \key_reg[6][4]$_DFFE_PN0P_  (.D(_03247_),
    .RN(net82),
    .CK(clknet_leaf_11_clk),
    .Q(\core.key[36] ),
    .QN(_19560_));
 DFFR_X1 \key_reg[6][5]$_DFFE_PN0P_  (.D(_03248_),
    .RN(net82),
    .CK(clknet_leaf_1_clk),
    .Q(\core.key[37] ),
    .QN(_19559_));
 DFFR_X1 \key_reg[6][6]$_DFFE_PN0P_  (.D(_03249_),
    .RN(net82),
    .CK(clknet_leaf_425_clk),
    .Q(\core.key[38] ),
    .QN(_19558_));
 DFFR_X1 \key_reg[6][7]$_DFFE_PN0P_  (.D(_03250_),
    .RN(net82),
    .CK(clknet_leaf_3_clk),
    .Q(\core.key[39] ),
    .QN(_19557_));
 DFFR_X2 \key_reg[6][8]$_DFFE_PN0P_  (.D(_03251_),
    .RN(net82),
    .CK(clknet_leaf_12_clk),
    .Q(\core.key[40] ),
    .QN(_19556_));
 DFFR_X1 \key_reg[6][9]$_DFFE_PN0P_  (.D(_03252_),
    .RN(net82),
    .CK(clknet_leaf_12_clk),
    .Q(\core.key[41] ),
    .QN(_19555_));
 DFFR_X1 \key_reg[7][0]$_DFFE_PN0P_  (.D(_03253_),
    .RN(net84),
    .CK(clknet_leaf_385_clk),
    .Q(\core.key[0] ),
    .QN(_19554_));
 DFFR_X1 \key_reg[7][10]$_DFFE_PN0P_  (.D(_03254_),
    .RN(net88),
    .CK(clknet_leaf_389_clk),
    .Q(\core.key[10] ),
    .QN(_19553_));
 DFFR_X1 \key_reg[7][11]$_DFFE_PN0P_  (.D(_03255_),
    .RN(net88),
    .CK(clknet_leaf_389_clk),
    .Q(\core.key[11] ),
    .QN(_19552_));
 DFFR_X1 \key_reg[7][12]$_DFFE_PN0P_  (.D(_03256_),
    .RN(net86),
    .CK(clknet_leaf_400_clk),
    .Q(\core.key[12] ),
    .QN(_19551_));
 DFFR_X2 \key_reg[7][13]$_DFFE_PN0P_  (.D(_03257_),
    .RN(net88),
    .CK(clknet_leaf_390_clk),
    .Q(\core.key[13] ),
    .QN(_19550_));
 DFFR_X1 \key_reg[7][14]$_DFFE_PN0P_  (.D(_03258_),
    .RN(net88),
    .CK(clknet_leaf_400_clk),
    .Q(\core.key[14] ),
    .QN(_19549_));
 DFFR_X2 \key_reg[7][15]$_DFFE_PN0P_  (.D(_03259_),
    .RN(net84),
    .CK(clknet_leaf_368_clk),
    .Q(\core.key[15] ),
    .QN(_19548_));
 DFFR_X1 \key_reg[7][16]$_DFFE_PN0P_  (.D(_03260_),
    .RN(net88),
    .CK(clknet_leaf_400_clk),
    .Q(\core.key[16] ),
    .QN(_19547_));
 DFFR_X1 \key_reg[7][17]$_DFFE_PN0P_  (.D(_03261_),
    .RN(net88),
    .CK(clknet_leaf_383_clk),
    .Q(\core.key[17] ),
    .QN(_19546_));
 DFFR_X1 \key_reg[7][18]$_DFFE_PN0P_  (.D(_03262_),
    .RN(net86),
    .CK(clknet_leaf_391_clk),
    .Q(\core.key[18] ),
    .QN(_19545_));
 DFFR_X1 \key_reg[7][19]$_DFFE_PN0P_  (.D(_03263_),
    .RN(net87),
    .CK(clknet_leaf_393_clk),
    .Q(\core.key[19] ),
    .QN(_19544_));
 DFFR_X1 \key_reg[7][1]$_DFFE_PN0P_  (.D(_03264_),
    .RN(net87),
    .CK(clknet_leaf_394_clk),
    .Q(\core.key[1] ),
    .QN(_19543_));
 DFFR_X1 \key_reg[7][20]$_DFFE_PN0P_  (.D(_03265_),
    .RN(net86),
    .CK(clknet_leaf_404_clk),
    .Q(\core.key[20] ),
    .QN(_19542_));
 DFFR_X1 \key_reg[7][21]$_DFFE_PN0P_  (.D(_03266_),
    .RN(net86),
    .CK(clknet_leaf_403_clk),
    .Q(\core.key[21] ),
    .QN(_19541_));
 DFFR_X1 \key_reg[7][22]$_DFFE_PN0P_  (.D(_03267_),
    .RN(net86),
    .CK(clknet_leaf_403_clk),
    .Q(\core.key[22] ),
    .QN(_19540_));
 DFFR_X1 \key_reg[7][23]$_DFFE_PN0P_  (.D(_03268_),
    .RN(net86),
    .CK(clknet_leaf_403_clk),
    .Q(\core.key[23] ),
    .QN(_19539_));
 DFFR_X1 \key_reg[7][24]$_DFFE_PN0P_  (.D(_03269_),
    .RN(net86),
    .CK(clknet_leaf_414_clk),
    .Q(\core.key[24] ),
    .QN(_00019_));
 DFFR_X1 \key_reg[7][25]$_DFFE_PN0P_  (.D(_03270_),
    .RN(net86),
    .CK(clknet_leaf_408_clk),
    .Q(\core.key[25] ),
    .QN(_00022_));
 DFFR_X1 \key_reg[7][26]$_DFFE_PN0P_  (.D(_03271_),
    .RN(net87),
    .CK(clknet_leaf_413_clk),
    .Q(\core.key[26] ),
    .QN(_00025_));
 DFFR_X1 \key_reg[7][27]$_DFFE_PN0P_  (.D(_03272_),
    .RN(net87),
    .CK(clknet_leaf_412_clk),
    .Q(\core.key[27] ),
    .QN(_00028_));
 DFFR_X1 \key_reg[7][28]$_DFFE_PN0P_  (.D(_03273_),
    .RN(net82),
    .CK(clknet_leaf_12_clk),
    .Q(\core.key[28] ),
    .QN(_00031_));
 DFFR_X1 \key_reg[7][29]$_DFFE_PN0P_  (.D(_03274_),
    .RN(net82),
    .CK(clknet_leaf_2_clk),
    .Q(\core.key[29] ),
    .QN(_00034_));
 DFFR_X1 \key_reg[7][2]$_DFFE_PN0P_  (.D(_03275_),
    .RN(net82),
    .CK(clknet_leaf_3_clk),
    .Q(\core.key[2] ),
    .QN(_19538_));
 DFFR_X1 \key_reg[7][30]$_DFFE_PN0P_  (.D(_03276_),
    .RN(net82),
    .CK(clknet_leaf_3_clk),
    .Q(\core.key[30] ),
    .QN(_00037_));
 DFFR_X1 \key_reg[7][31]$_DFFE_PN0P_  (.D(_03277_),
    .RN(net82),
    .CK(clknet_leaf_425_clk),
    .Q(\core.key[31] ),
    .QN(_00040_));
 DFFR_X1 \key_reg[7][3]$_DFFE_PN0P_  (.D(_03278_),
    .RN(net82),
    .CK(clknet_leaf_0_clk),
    .Q(\core.key[3] ),
    .QN(_19537_));
 DFFR_X1 \key_reg[7][4]$_DFFE_PN0P_  (.D(_03279_),
    .RN(net82),
    .CK(clknet_leaf_11_clk),
    .Q(\core.key[4] ),
    .QN(_19536_));
 DFFR_X1 \key_reg[7][5]$_DFFE_PN0P_  (.D(_03280_),
    .RN(net82),
    .CK(clknet_leaf_1_clk),
    .Q(\core.key[5] ),
    .QN(_19535_));
 DFFR_X1 \key_reg[7][6]$_DFFE_PN0P_  (.D(_03281_),
    .RN(net82),
    .CK(clknet_leaf_425_clk),
    .Q(\core.key[6] ),
    .QN(_19534_));
 DFFR_X1 \key_reg[7][7]$_DFFE_PN0P_  (.D(_03282_),
    .RN(net82),
    .CK(clknet_leaf_4_clk),
    .Q(\core.key[7] ),
    .QN(_19533_));
 DFFR_X2 \key_reg[7][8]$_DFFE_PN0P_  (.D(_03283_),
    .RN(net82),
    .CK(clknet_leaf_1_clk),
    .Q(\core.key[8] ),
    .QN(_19532_));
 DFFR_X2 \key_reg[7][9]$_DFFE_PN0P_  (.D(_03284_),
    .RN(net82),
    .CK(clknet_leaf_1_clk),
    .Q(\core.key[9] ),
    .QN(_19531_));
 DFFR_X1 \keylen_reg$_DFFE_PN0P_  (.D(_03285_),
    .RN(net84),
    .CK(clknet_leaf_354_clk),
    .Q(\core.dec_block.keylen ),
    .QN(_22091_));
 DFFR_X1 \next_reg$_DFF_PN0_  (.D(next_new),
    .RN(net90),
    .CK(clknet_leaf_309_clk),
    .Q(\core.next ),
    .QN(_21961_));
 DFFR_X1 \ready_reg$_DFF_PN0_  (.D(\core.ready ),
    .RN(net83),
    .CK(clknet_leaf_315_clk),
    .Q(ready_reg),
    .QN(_21962_));
 DFFR_X1 \result_reg[0]$_DFF_PN0_  (.D(\core.muxed_new_block[0] ),
    .RN(net83),
    .CK(clknet_leaf_326_clk),
    .Q(\result_reg[0] ),
    .QN(_21963_));
 DFFR_X1 \result_reg[100]$_DFF_PN0_  (.D(\core.muxed_new_block[100] ),
    .RN(net83),
    .CK(clknet_leaf_328_clk),
    .Q(\result_reg[100] ),
    .QN(_21964_));
 DFFR_X1 \result_reg[101]$_DFF_PN0_  (.D(\core.muxed_new_block[101] ),
    .RN(net83),
    .CK(clknet_leaf_327_clk),
    .Q(\result_reg[101] ),
    .QN(_21965_));
 DFFR_X1 \result_reg[102]$_DFF_PN0_  (.D(\core.muxed_new_block[102] ),
    .RN(net90),
    .CK(clknet_leaf_307_clk),
    .Q(\result_reg[102] ),
    .QN(_21966_));
 DFFR_X1 \result_reg[103]$_DFF_PN0_  (.D(\core.muxed_new_block[103] ),
    .RN(net83),
    .CK(clknet_leaf_324_clk),
    .Q(\result_reg[103] ),
    .QN(_21967_));
 DFFR_X1 \result_reg[104]$_DFF_PN0_  (.D(\core.muxed_new_block[104] ),
    .RN(net83),
    .CK(clknet_leaf_329_clk),
    .Q(\result_reg[104] ),
    .QN(_21968_));
 DFFR_X1 \result_reg[105]$_DFF_PN0_  (.D(\core.muxed_new_block[105] ),
    .RN(net83),
    .CK(clknet_leaf_329_clk),
    .Q(\result_reg[105] ),
    .QN(_21969_));
 DFFR_X1 \result_reg[106]$_DFF_PN0_  (.D(\core.muxed_new_block[106] ),
    .RN(net83),
    .CK(clknet_leaf_324_clk),
    .Q(\result_reg[106] ),
    .QN(_21970_));
 DFFR_X1 \result_reg[107]$_DFF_PN0_  (.D(\core.muxed_new_block[107] ),
    .RN(net90),
    .CK(clknet_leaf_318_clk),
    .Q(\result_reg[107] ),
    .QN(_21971_));
 DFFR_X1 \result_reg[108]$_DFF_PN0_  (.D(\core.muxed_new_block[108] ),
    .RN(net83),
    .CK(clknet_leaf_327_clk),
    .Q(\result_reg[108] ),
    .QN(_21972_));
 DFFR_X1 \result_reg[109]$_DFF_PN0_  (.D(\core.muxed_new_block[109] ),
    .RN(net83),
    .CK(clknet_leaf_323_clk),
    .Q(\result_reg[109] ),
    .QN(_21973_));
 DFFR_X1 \result_reg[10]$_DFF_PN0_  (.D(\core.muxed_new_block[10] ),
    .RN(net83),
    .CK(clknet_leaf_324_clk),
    .Q(\result_reg[10] ),
    .QN(_21974_));
 DFFR_X1 \result_reg[110]$_DFF_PN0_  (.D(\core.muxed_new_block[110] ),
    .RN(net90),
    .CK(clknet_leaf_321_clk),
    .Q(\result_reg[110] ),
    .QN(_21975_));
 DFFR_X1 \result_reg[111]$_DFF_PN0_  (.D(\core.muxed_new_block[111] ),
    .RN(net90),
    .CK(clknet_leaf_322_clk),
    .Q(\result_reg[111] ),
    .QN(_21976_));
 DFFR_X1 \result_reg[112]$_DFF_PN0_  (.D(\core.muxed_new_block[112] ),
    .RN(net83),
    .CK(clknet_leaf_325_clk),
    .Q(\result_reg[112] ),
    .QN(_21977_));
 DFFR_X1 \result_reg[113]$_DFF_PN0_  (.D(\core.muxed_new_block[113] ),
    .RN(net90),
    .CK(clknet_leaf_321_clk),
    .Q(\result_reg[113] ),
    .QN(_21978_));
 DFFR_X1 \result_reg[114]$_DFF_PN0_  (.D(\core.muxed_new_block[114] ),
    .RN(net83),
    .CK(clknet_leaf_327_clk),
    .Q(\result_reg[114] ),
    .QN(_21979_));
 DFFR_X1 \result_reg[115]$_DFF_PN0_  (.D(\core.muxed_new_block[115] ),
    .RN(net90),
    .CK(clknet_leaf_319_clk),
    .Q(\result_reg[115] ),
    .QN(_21980_));
 DFFR_X1 \result_reg[116]$_DFF_PN0_  (.D(\core.muxed_new_block[116] ),
    .RN(net90),
    .CK(clknet_leaf_319_clk),
    .Q(\result_reg[116] ),
    .QN(_21981_));
 DFFR_X1 \result_reg[117]$_DFF_PN0_  (.D(\core.muxed_new_block[117] ),
    .RN(net90),
    .CK(clknet_leaf_317_clk),
    .Q(\result_reg[117] ),
    .QN(_21982_));
 DFFR_X1 \result_reg[118]$_DFF_PN0_  (.D(\core.muxed_new_block[118] ),
    .RN(net90),
    .CK(clknet_leaf_317_clk),
    .Q(\result_reg[118] ),
    .QN(_21983_));
 DFFR_X1 \result_reg[119]$_DFF_PN0_  (.D(\core.muxed_new_block[119] ),
    .RN(net90),
    .CK(clknet_leaf_320_clk),
    .Q(\result_reg[119] ),
    .QN(_21984_));
 DFFR_X1 \result_reg[11]$_DFF_PN0_  (.D(\core.muxed_new_block[11] ),
    .RN(net90),
    .CK(clknet_leaf_318_clk),
    .Q(\result_reg[11] ),
    .QN(_21985_));
 DFFR_X1 \result_reg[120]$_DFF_PN0_  (.D(\core.muxed_new_block[120] ),
    .RN(net90),
    .CK(clknet_leaf_317_clk),
    .Q(\result_reg[120] ),
    .QN(_21986_));
 DFFR_X1 \result_reg[121]$_DFF_PN0_  (.D(\core.muxed_new_block[121] ),
    .RN(net90),
    .CK(clknet_leaf_320_clk),
    .Q(\result_reg[121] ),
    .QN(_21987_));
 DFFR_X1 \result_reg[122]$_DFF_PN0_  (.D(\core.muxed_new_block[122] ),
    .RN(net90),
    .CK(clknet_leaf_317_clk),
    .Q(\result_reg[122] ),
    .QN(_21988_));
 DFFR_X1 \result_reg[123]$_DFF_PN0_  (.D(\core.muxed_new_block[123] ),
    .RN(net90),
    .CK(clknet_leaf_320_clk),
    .Q(\result_reg[123] ),
    .QN(_21989_));
 DFFR_X1 \result_reg[124]$_DFF_PN0_  (.D(\core.muxed_new_block[124] ),
    .RN(net90),
    .CK(clknet_leaf_313_clk),
    .Q(\result_reg[124] ),
    .QN(_21990_));
 DFFR_X1 \result_reg[125]$_DFF_PN0_  (.D(\core.muxed_new_block[125] ),
    .RN(net83),
    .CK(clknet_leaf_335_clk),
    .Q(\result_reg[125] ),
    .QN(_21991_));
 DFFR_X1 \result_reg[126]$_DFF_PN0_  (.D(\core.muxed_new_block[126] ),
    .RN(net83),
    .CK(clknet_leaf_328_clk),
    .Q(\result_reg[126] ),
    .QN(_21992_));
 DFFR_X1 \result_reg[127]$_DFF_PN0_  (.D(\core.muxed_new_block[127] ),
    .RN(net90),
    .CK(clknet_leaf_322_clk),
    .Q(\result_reg[127] ),
    .QN(_21993_));
 DFFR_X1 \result_reg[12]$_DFF_PN0_  (.D(\core.muxed_new_block[12] ),
    .RN(net83),
    .CK(clknet_leaf_327_clk),
    .Q(\result_reg[12] ),
    .QN(_21994_));
 DFFR_X1 \result_reg[13]$_DFF_PN0_  (.D(\core.muxed_new_block[13] ),
    .RN(net83),
    .CK(clknet_leaf_323_clk),
    .Q(\result_reg[13] ),
    .QN(_21995_));
 DFFR_X1 \result_reg[14]$_DFF_PN0_  (.D(\core.muxed_new_block[14] ),
    .RN(net90),
    .CK(clknet_leaf_322_clk),
    .Q(\result_reg[14] ),
    .QN(_21996_));
 DFFR_X1 \result_reg[15]$_DFF_PN0_  (.D(\core.muxed_new_block[15] ),
    .RN(net90),
    .CK(clknet_leaf_322_clk),
    .Q(\result_reg[15] ),
    .QN(_21997_));
 DFFR_X1 \result_reg[16]$_DFF_PN0_  (.D(\core.muxed_new_block[16] ),
    .RN(net83),
    .CK(clknet_leaf_325_clk),
    .Q(\result_reg[16] ),
    .QN(_21998_));
 DFFR_X1 \result_reg[17]$_DFF_PN0_  (.D(\core.muxed_new_block[17] ),
    .RN(net83),
    .CK(clknet_leaf_325_clk),
    .Q(\result_reg[17] ),
    .QN(_21999_));
 DFFR_X1 \result_reg[18]$_DFF_PN0_  (.D(\core.muxed_new_block[18] ),
    .RN(net83),
    .CK(clknet_leaf_327_clk),
    .Q(\result_reg[18] ),
    .QN(_22000_));
 DFFR_X1 \result_reg[19]$_DFF_PN0_  (.D(\core.muxed_new_block[19] ),
    .RN(net90),
    .CK(clknet_leaf_319_clk),
    .Q(\result_reg[19] ),
    .QN(_22001_));
 DFFR_X1 \result_reg[1]$_DFF_PN0_  (.D(\core.muxed_new_block[1] ),
    .RN(net83),
    .CK(clknet_leaf_315_clk),
    .Q(\result_reg[1] ),
    .QN(_22002_));
 DFFR_X1 \result_reg[20]$_DFF_PN0_  (.D(\core.muxed_new_block[20] ),
    .RN(net90),
    .CK(clknet_leaf_318_clk),
    .Q(\result_reg[20] ),
    .QN(_22003_));
 DFFR_X1 \result_reg[21]$_DFF_PN0_  (.D(\core.muxed_new_block[21] ),
    .RN(net90),
    .CK(clknet_leaf_317_clk),
    .Q(\result_reg[21] ),
    .QN(_22004_));
 DFFR_X1 \result_reg[22]$_DFF_PN0_  (.D(\core.muxed_new_block[22] ),
    .RN(net90),
    .CK(clknet_leaf_316_clk),
    .Q(\result_reg[22] ),
    .QN(_22005_));
 DFFR_X1 \result_reg[23]$_DFF_PN0_  (.D(\core.muxed_new_block[23] ),
    .RN(net90),
    .CK(clknet_leaf_322_clk),
    .Q(\result_reg[23] ),
    .QN(_22006_));
 DFFR_X1 \result_reg[24]$_DFF_PN0_  (.D(\core.muxed_new_block[24] ),
    .RN(net83),
    .CK(clknet_leaf_323_clk),
    .Q(\result_reg[24] ),
    .QN(_22007_));
 DFFR_X1 \result_reg[25]$_DFF_PN0_  (.D(\core.muxed_new_block[25] ),
    .RN(net90),
    .CK(clknet_leaf_321_clk),
    .Q(\result_reg[25] ),
    .QN(_22008_));
 DFFR_X1 \result_reg[26]$_DFF_PN0_  (.D(\core.muxed_new_block[26] ),
    .RN(net90),
    .CK(clknet_leaf_317_clk),
    .Q(\result_reg[26] ),
    .QN(_22009_));
 DFFR_X1 \result_reg[27]$_DFF_PN0_  (.D(\core.muxed_new_block[27] ),
    .RN(net90),
    .CK(clknet_leaf_320_clk),
    .Q(\result_reg[27] ),
    .QN(_22010_));
 DFFR_X1 \result_reg[28]$_DFF_PN0_  (.D(\core.muxed_new_block[28] ),
    .RN(net90),
    .CK(clknet_leaf_313_clk),
    .Q(\result_reg[28] ),
    .QN(_22011_));
 DFFR_X1 \result_reg[29]$_DFF_PN0_  (.D(\core.muxed_new_block[29] ),
    .RN(net83),
    .CK(clknet_leaf_315_clk),
    .Q(\result_reg[29] ),
    .QN(_22012_));
 DFFR_X1 \result_reg[2]$_DFF_PN0_  (.D(\core.muxed_new_block[2] ),
    .RN(net83),
    .CK(clknet_leaf_314_clk),
    .Q(\result_reg[2] ),
    .QN(_22013_));
 DFFR_X1 \result_reg[30]$_DFF_PN0_  (.D(\core.muxed_new_block[30] ),
    .RN(net83),
    .CK(clknet_leaf_328_clk),
    .Q(\result_reg[30] ),
    .QN(_22014_));
 DFFR_X1 \result_reg[31]$_DFF_PN0_  (.D(\core.muxed_new_block[31] ),
    .RN(net90),
    .CK(clknet_leaf_321_clk),
    .Q(\result_reg[31] ),
    .QN(_22015_));
 DFFR_X1 \result_reg[32]$_DFF_PN0_  (.D(\core.muxed_new_block[32] ),
    .RN(net83),
    .CK(clknet_leaf_326_clk),
    .Q(\result_reg[32] ),
    .QN(_22016_));
 DFFR_X1 \result_reg[33]$_DFF_PN0_  (.D(\core.muxed_new_block[33] ),
    .RN(net83),
    .CK(clknet_leaf_315_clk),
    .Q(\result_reg[33] ),
    .QN(_22017_));
 DFFR_X1 \result_reg[34]$_DFF_PN0_  (.D(\core.muxed_new_block[34] ),
    .RN(net83),
    .CK(clknet_leaf_314_clk),
    .Q(\result_reg[34] ),
    .QN(_22018_));
 DFFR_X1 \result_reg[35]$_DFF_PN0_  (.D(\core.muxed_new_block[35] ),
    .RN(net83),
    .CK(clknet_leaf_314_clk),
    .Q(\result_reg[35] ),
    .QN(_22019_));
 DFFR_X1 \result_reg[36]$_DFF_PN0_  (.D(\core.muxed_new_block[36] ),
    .RN(net83),
    .CK(clknet_leaf_323_clk),
    .Q(\result_reg[36] ),
    .QN(_22020_));
 DFFR_X1 \result_reg[37]$_DFF_PN0_  (.D(\core.muxed_new_block[37] ),
    .RN(net90),
    .CK(clknet_leaf_313_clk),
    .Q(\result_reg[37] ),
    .QN(_22021_));
 DFFR_X1 \result_reg[38]$_DFF_PN0_  (.D(\core.muxed_new_block[38] ),
    .RN(net90),
    .CK(clknet_leaf_320_clk),
    .Q(\result_reg[38] ),
    .QN(_22022_));
 DFFR_X1 \result_reg[39]$_DFF_PN0_  (.D(\core.muxed_new_block[39] ),
    .RN(net90),
    .CK(clknet_leaf_316_clk),
    .Q(\result_reg[39] ),
    .QN(_22023_));
 DFFR_X1 \result_reg[3]$_DFF_PN0_  (.D(\core.muxed_new_block[3] ),
    .RN(net83),
    .CK(clknet_leaf_314_clk),
    .Q(\result_reg[3] ),
    .QN(_22024_));
 DFFR_X1 \result_reg[40]$_DFF_PN0_  (.D(\core.muxed_new_block[40] ),
    .RN(net90),
    .CK(clknet_leaf_309_clk),
    .Q(\result_reg[40] ),
    .QN(_22025_));
 DFFR_X1 \result_reg[41]$_DFF_PN0_  (.D(\core.muxed_new_block[41] ),
    .RN(net83),
    .CK(clknet_leaf_329_clk),
    .Q(\result_reg[41] ),
    .QN(_22026_));
 DFFR_X1 \result_reg[42]$_DFF_PN0_  (.D(\core.muxed_new_block[42] ),
    .RN(net83),
    .CK(clknet_leaf_324_clk),
    .Q(\result_reg[42] ),
    .QN(_22027_));
 DFFR_X1 \result_reg[43]$_DFF_PN0_  (.D(\core.muxed_new_block[43] ),
    .RN(net90),
    .CK(clknet_leaf_318_clk),
    .Q(\result_reg[43] ),
    .QN(_22028_));
 DFFR_X1 \result_reg[44]$_DFF_PN0_  (.D(\core.muxed_new_block[44] ),
    .RN(net83),
    .CK(clknet_leaf_327_clk),
    .Q(\result_reg[44] ),
    .QN(_22029_));
 DFFR_X1 \result_reg[45]$_DFF_PN0_  (.D(\core.muxed_new_block[45] ),
    .RN(net90),
    .CK(clknet_leaf_308_clk),
    .Q(\result_reg[45] ),
    .QN(_22030_));
 DFFR_X1 \result_reg[46]$_DFF_PN0_  (.D(\core.muxed_new_block[46] ),
    .RN(net90),
    .CK(clknet_leaf_307_clk),
    .Q(\result_reg[46] ),
    .QN(_22031_));
 DFFR_X1 \result_reg[47]$_DFF_PN0_  (.D(\core.muxed_new_block[47] ),
    .RN(net90),
    .CK(clknet_leaf_322_clk),
    .Q(\result_reg[47] ),
    .QN(_22032_));
 DFFR_X1 \result_reg[48]$_DFF_PN0_  (.D(\core.muxed_new_block[48] ),
    .RN(net83),
    .CK(clknet_leaf_325_clk),
    .Q(\result_reg[48] ),
    .QN(_22033_));
 DFFR_X1 \result_reg[49]$_DFF_PN0_  (.D(\core.muxed_new_block[49] ),
    .RN(net90),
    .CK(clknet_leaf_325_clk),
    .Q(\result_reg[49] ),
    .QN(_22034_));
 DFFR_X1 \result_reg[4]$_DFF_PN0_  (.D(\core.muxed_new_block[4] ),
    .RN(net83),
    .CK(clknet_leaf_323_clk),
    .Q(\result_reg[4] ),
    .QN(_22035_));
 DFFR_X1 \result_reg[50]$_DFF_PN0_  (.D(\core.muxed_new_block[50] ),
    .RN(net83),
    .CK(clknet_leaf_326_clk),
    .Q(\result_reg[50] ),
    .QN(_22036_));
 DFFR_X1 \result_reg[51]$_DFF_PN0_  (.D(\core.muxed_new_block[51] ),
    .RN(net90),
    .CK(clknet_leaf_307_clk),
    .Q(\result_reg[51] ),
    .QN(_22037_));
 DFFR_X1 \result_reg[52]$_DFF_PN0_  (.D(\core.muxed_new_block[52] ),
    .RN(net90),
    .CK(clknet_leaf_319_clk),
    .Q(\result_reg[52] ),
    .QN(_22038_));
 DFFR_X1 \result_reg[53]$_DFF_PN0_  (.D(\core.muxed_new_block[53] ),
    .RN(net90),
    .CK(clknet_leaf_308_clk),
    .Q(\result_reg[53] ),
    .QN(_22039_));
 DFFR_X1 \result_reg[54]$_DFF_PN0_  (.D(\core.muxed_new_block[54] ),
    .RN(net90),
    .CK(clknet_leaf_316_clk),
    .Q(\result_reg[54] ),
    .QN(_22040_));
 DFFR_X1 \result_reg[55]$_DFF_PN0_  (.D(\core.muxed_new_block[55] ),
    .RN(net90),
    .CK(clknet_leaf_322_clk),
    .Q(\result_reg[55] ),
    .QN(_22041_));
 DFFR_X1 \result_reg[56]$_DFF_PN0_  (.D(\core.muxed_new_block[56] ),
    .RN(net83),
    .CK(clknet_leaf_323_clk),
    .Q(\result_reg[56] ),
    .QN(_22042_));
 DFFR_X1 \result_reg[57]$_DFF_PN0_  (.D(\core.muxed_new_block[57] ),
    .RN(net90),
    .CK(clknet_leaf_321_clk),
    .Q(\result_reg[57] ),
    .QN(_22043_));
 DFFR_X1 \result_reg[58]$_DFF_PN0_  (.D(\core.muxed_new_block[58] ),
    .RN(net90),
    .CK(clknet_leaf_317_clk),
    .Q(\result_reg[58] ),
    .QN(_22044_));
 DFFR_X1 \result_reg[59]$_DFF_PN0_  (.D(\core.muxed_new_block[59] ),
    .RN(net90),
    .CK(clknet_leaf_318_clk),
    .Q(\result_reg[59] ),
    .QN(_22045_));
 DFFR_X1 \result_reg[5]$_DFF_PN0_  (.D(\core.muxed_new_block[5] ),
    .RN(net90),
    .CK(clknet_leaf_313_clk),
    .Q(\result_reg[5] ),
    .QN(_22046_));
 DFFR_X1 \result_reg[60]$_DFF_PN0_  (.D(\core.muxed_new_block[60] ),
    .RN(net83),
    .CK(clknet_leaf_314_clk),
    .Q(\result_reg[60] ),
    .QN(_22047_));
 DFFR_X1 \result_reg[61]$_DFF_PN0_  (.D(\core.muxed_new_block[61] ),
    .RN(net83),
    .CK(clknet_leaf_335_clk),
    .Q(\result_reg[61] ),
    .QN(_22048_));
 DFFR_X1 \result_reg[62]$_DFF_PN0_  (.D(\core.muxed_new_block[62] ),
    .RN(net83),
    .CK(clknet_leaf_328_clk),
    .Q(\result_reg[62] ),
    .QN(_22049_));
 DFFR_X1 \result_reg[63]$_DFF_PN0_  (.D(\core.muxed_new_block[63] ),
    .RN(net90),
    .CK(clknet_leaf_318_clk),
    .Q(\result_reg[63] ),
    .QN(_22050_));
 DFFR_X1 \result_reg[64]$_DFF_PN0_  (.D(\core.muxed_new_block[64] ),
    .RN(net83),
    .CK(clknet_leaf_326_clk),
    .Q(\result_reg[64] ),
    .QN(_22051_));
 DFFR_X1 \result_reg[65]$_DFF_PN0_  (.D(\core.muxed_new_block[65] ),
    .RN(net83),
    .CK(clknet_leaf_330_clk),
    .Q(\result_reg[65] ),
    .QN(_22052_));
 DFFR_X1 \result_reg[66]$_DFF_PN0_  (.D(\core.muxed_new_block[66] ),
    .RN(net83),
    .CK(clknet_leaf_330_clk),
    .Q(\result_reg[66] ),
    .QN(_22053_));
 DFFR_X1 \result_reg[67]$_DFF_PN0_  (.D(\core.muxed_new_block[67] ),
    .RN(net83),
    .CK(clknet_leaf_329_clk),
    .Q(\result_reg[67] ),
    .QN(_22054_));
 DFFR_X1 \result_reg[68]$_DFF_PN0_  (.D(\core.muxed_new_block[68] ),
    .RN(net83),
    .CK(clknet_leaf_328_clk),
    .Q(\result_reg[68] ),
    .QN(_22055_));
 DFFR_X1 \result_reg[69]$_DFF_PN0_  (.D(\core.muxed_new_block[69] ),
    .RN(net83),
    .CK(clknet_leaf_328_clk),
    .Q(\result_reg[69] ),
    .QN(_22056_));
 DFFR_X1 \result_reg[6]$_DFF_PN0_  (.D(\core.muxed_new_block[6] ),
    .RN(net90),
    .CK(clknet_leaf_319_clk),
    .Q(\result_reg[6] ),
    .QN(_22057_));
 DFFR_X1 \result_reg[70]$_DFF_PN0_  (.D(\core.muxed_new_block[70] ),
    .RN(net90),
    .CK(clknet_leaf_319_clk),
    .Q(\result_reg[70] ),
    .QN(_22058_));
 DFFR_X1 \result_reg[71]$_DFF_PN0_  (.D(\core.muxed_new_block[71] ),
    .RN(net83),
    .CK(clknet_leaf_324_clk),
    .Q(\result_reg[71] ),
    .QN(_22059_));
 DFFR_X1 \result_reg[72]$_DFF_PN0_  (.D(\core.muxed_new_block[72] ),
    .RN(net83),
    .CK(clknet_leaf_326_clk),
    .Q(\result_reg[72] ),
    .QN(_22060_));
 DFFR_X1 \result_reg[73]$_DFF_PN0_  (.D(\core.muxed_new_block[73] ),
    .RN(net83),
    .CK(clknet_leaf_326_clk),
    .Q(\result_reg[73] ),
    .QN(_22061_));
 DFFR_X1 \result_reg[74]$_DFF_PN0_  (.D(\core.muxed_new_block[74] ),
    .RN(net83),
    .CK(clknet_leaf_324_clk),
    .Q(\result_reg[74] ),
    .QN(_22062_));
 DFFR_X1 \result_reg[75]$_DFF_PN0_  (.D(\core.muxed_new_block[75] ),
    .RN(net90),
    .CK(clknet_leaf_318_clk),
    .Q(\result_reg[75] ),
    .QN(_22063_));
 DFFR_X1 \result_reg[76]$_DFF_PN0_  (.D(\core.muxed_new_block[76] ),
    .RN(net83),
    .CK(clknet_leaf_327_clk),
    .Q(\result_reg[76] ),
    .QN(_22064_));
 DFFR_X1 \result_reg[77]$_DFF_PN0_  (.D(\core.muxed_new_block[77] ),
    .RN(net83),
    .CK(clknet_leaf_323_clk),
    .Q(\result_reg[77] ),
    .QN(_22065_));
 DFFR_X1 \result_reg[78]$_DFF_PN0_  (.D(\core.muxed_new_block[78] ),
    .RN(net90),
    .CK(clknet_leaf_321_clk),
    .Q(\result_reg[78] ),
    .QN(_22066_));
 DFFR_X1 \result_reg[79]$_DFF_PN0_  (.D(\core.muxed_new_block[79] ),
    .RN(net90),
    .CK(clknet_leaf_318_clk),
    .Q(\result_reg[79] ),
    .QN(_22067_));
 DFFR_X1 \result_reg[7]$_DFF_PN0_  (.D(\core.muxed_new_block[7] ),
    .RN(net90),
    .CK(clknet_leaf_316_clk),
    .Q(\result_reg[7] ),
    .QN(_22068_));
 DFFR_X1 \result_reg[80]$_DFF_PN0_  (.D(\core.muxed_new_block[80] ),
    .RN(net83),
    .CK(clknet_leaf_325_clk),
    .Q(\result_reg[80] ),
    .QN(_22069_));
 DFFR_X1 \result_reg[81]$_DFF_PN0_  (.D(\core.muxed_new_block[81] ),
    .RN(net90),
    .CK(clknet_leaf_321_clk),
    .Q(\result_reg[81] ),
    .QN(_22070_));
 DFFR_X1 \result_reg[82]$_DFF_PN0_  (.D(\core.muxed_new_block[82] ),
    .RN(net83),
    .CK(clknet_leaf_324_clk),
    .Q(\result_reg[82] ),
    .QN(_22071_));
 DFFR_X1 \result_reg[83]$_DFF_PN0_  (.D(\core.muxed_new_block[83] ),
    .RN(net90),
    .CK(clknet_leaf_307_clk),
    .Q(\result_reg[83] ),
    .QN(_22072_));
 DFFR_X1 \result_reg[84]$_DFF_PN0_  (.D(\core.muxed_new_block[84] ),
    .RN(net90),
    .CK(clknet_leaf_319_clk),
    .Q(\result_reg[84] ),
    .QN(_22073_));
 DFFR_X1 \result_reg[85]$_DFF_PN0_  (.D(\core.muxed_new_block[85] ),
    .RN(net90),
    .CK(clknet_leaf_308_clk),
    .Q(\result_reg[85] ),
    .QN(_22074_));
 DFFR_X1 \result_reg[86]$_DFF_PN0_  (.D(\core.muxed_new_block[86] ),
    .RN(net90),
    .CK(clknet_leaf_308_clk),
    .Q(\result_reg[86] ),
    .QN(_22075_));
 DFFR_X1 \result_reg[87]$_DFF_PN0_  (.D(\core.muxed_new_block[87] ),
    .RN(net90),
    .CK(clknet_leaf_307_clk),
    .Q(\result_reg[87] ),
    .QN(_22076_));
 DFFR_X1 \result_reg[88]$_DFF_PN0_  (.D(\core.muxed_new_block[88] ),
    .RN(net83),
    .CK(clknet_leaf_323_clk),
    .Q(\result_reg[88] ),
    .QN(_22077_));
 DFFR_X1 \result_reg[89]$_DFF_PN0_  (.D(\core.muxed_new_block[89] ),
    .RN(net90),
    .CK(clknet_leaf_320_clk),
    .Q(\result_reg[89] ),
    .QN(_22078_));
 DFFR_X1 \result_reg[8]$_DFF_PN0_  (.D(\core.muxed_new_block[8] ),
    .RN(net83),
    .CK(clknet_leaf_328_clk),
    .Q(\result_reg[8] ),
    .QN(_22079_));
 DFFR_X1 \result_reg[90]$_DFF_PN0_  (.D(\core.muxed_new_block[90] ),
    .RN(net90),
    .CK(clknet_leaf_317_clk),
    .Q(\result_reg[90] ),
    .QN(_22080_));
 DFFR_X1 \result_reg[91]$_DFF_PN0_  (.D(\core.muxed_new_block[91] ),
    .RN(net90),
    .CK(clknet_leaf_320_clk),
    .Q(\result_reg[91] ),
    .QN(_22081_));
 DFFR_X1 \result_reg[92]$_DFF_PN0_  (.D(\core.muxed_new_block[92] ),
    .RN(net83),
    .CK(clknet_leaf_315_clk),
    .Q(\result_reg[92] ),
    .QN(_22082_));
 DFFR_X1 \result_reg[93]$_DFF_PN0_  (.D(\core.muxed_new_block[93] ),
    .RN(net83),
    .CK(clknet_leaf_315_clk),
    .Q(\result_reg[93] ),
    .QN(_22083_));
 DFFR_X1 \result_reg[94]$_DFF_PN0_  (.D(\core.muxed_new_block[94] ),
    .RN(net83),
    .CK(clknet_leaf_328_clk),
    .Q(\result_reg[94] ),
    .QN(_22084_));
 DFFR_X1 \result_reg[95]$_DFF_PN0_  (.D(\core.muxed_new_block[95] ),
    .RN(net90),
    .CK(clknet_leaf_322_clk),
    .Q(\result_reg[95] ),
    .QN(_22085_));
 DFFR_X1 \result_reg[96]$_DFF_PN0_  (.D(\core.muxed_new_block[96] ),
    .RN(net83),
    .CK(clknet_leaf_326_clk),
    .Q(\result_reg[96] ),
    .QN(_22086_));
 DFFR_X1 \result_reg[97]$_DFF_PN0_  (.D(\core.muxed_new_block[97] ),
    .RN(net83),
    .CK(clknet_leaf_331_clk),
    .Q(\result_reg[97] ),
    .QN(_22087_));
 DFFR_X1 \result_reg[98]$_DFF_PN0_  (.D(\core.muxed_new_block[98] ),
    .RN(net83),
    .CK(clknet_leaf_330_clk),
    .Q(\result_reg[98] ),
    .QN(_22088_));
 DFFR_X1 \result_reg[99]$_DFF_PN0_  (.D(\core.muxed_new_block[99] ),
    .RN(net83),
    .CK(clknet_leaf_329_clk),
    .Q(\result_reg[99] ),
    .QN(_22089_));
 DFFR_X1 \result_reg[9]$_DFF_PN0_  (.D(\core.muxed_new_block[9] ),
    .RN(net83),
    .CK(clknet_leaf_330_clk),
    .Q(\result_reg[9] ),
    .QN(_22090_));
 DFFR_X1 \valid_reg$_DFF_PN0_  (.D(\core.result_valid ),
    .RN(net83),
    .CK(clknet_leaf_315_clk),
    .Q(valid_reg),
    .QN(_19530_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_447 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_448 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_449 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_450 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_451 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_452 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_673 ();
 BUF_X2 wire9 (.A(_12677_),
    .Z(net9));
 BUF_X2 wire10 (.A(_12427_),
    .Z(net10));
 BUF_X2 wire11 (.A(_11995_),
    .Z(net11));
 BUF_X2 wire12 (.A(_11834_),
    .Z(net12));
 CLKBUF_X2 wire13 (.A(_12020_),
    .Z(net13));
 BUF_X1 max_cap14 (.A(_08660_),
    .Z(net14));
 BUF_X1 max_cap15 (.A(_18152_),
    .Z(net15));
 BUF_X4 input1 (.A(address[1]),
    .Z(net1));
 CLKBUF_X3 input2 (.A(address[2]),
    .Z(net2));
 BUF_X2 input3 (.A(address[3]),
    .Z(net3));
 CLKBUF_X3 input4 (.A(address[4]),
    .Z(net4));
 CLKBUF_X2 input5 (.A(address[5]),
    .Z(net5));
 BUF_X2 input6 (.A(address[6]),
    .Z(net6));
 BUF_X2 input7 (.A(address[7]),
    .Z(net7));
 CLKBUF_X3 input8 (.A(cs),
    .Z(net8));
 BUF_X32 input9 (.A(reset_n),
    .Z(net16));
 BUF_X2 input10 (.A(we),
    .Z(net17));
 CLKBUF_X3 input11 (.A(write_data[0]),
    .Z(net18));
 BUF_X2 input12 (.A(write_data[10]),
    .Z(net19));
 BUF_X2 input13 (.A(write_data[11]),
    .Z(net20));
 BUF_X2 input14 (.A(write_data[12]),
    .Z(net21));
 BUF_X2 input15 (.A(write_data[13]),
    .Z(net22));
 BUF_X2 input16 (.A(write_data[14]),
    .Z(net23));
 BUF_X2 input17 (.A(write_data[15]),
    .Z(net24));
 BUF_X2 input18 (.A(write_data[16]),
    .Z(net25));
 BUF_X2 input19 (.A(write_data[17]),
    .Z(net26));
 BUF_X2 input20 (.A(write_data[18]),
    .Z(net27));
 BUF_X2 input21 (.A(write_data[19]),
    .Z(net28));
 BUF_X2 input22 (.A(write_data[1]),
    .Z(net29));
 CLKBUF_X2 input23 (.A(write_data[20]),
    .Z(net30));
 BUF_X2 input24 (.A(write_data[21]),
    .Z(net31));
 CLKBUF_X2 input25 (.A(write_data[22]),
    .Z(net32));
 CLKBUF_X2 input26 (.A(write_data[23]),
    .Z(net33));
 BUF_X2 input27 (.A(write_data[24]),
    .Z(net34));
 BUF_X2 input28 (.A(write_data[25]),
    .Z(net35));
 BUF_X2 input29 (.A(write_data[26]),
    .Z(net36));
 BUF_X2 input30 (.A(write_data[27]),
    .Z(net37));
 CLKBUF_X2 input31 (.A(write_data[28]),
    .Z(net38));
 BUF_X1 input32 (.A(write_data[29]),
    .Z(net39));
 BUF_X1 input33 (.A(write_data[2]),
    .Z(net40));
 BUF_X1 input34 (.A(write_data[30]),
    .Z(net41));
 BUF_X2 input35 (.A(write_data[31]),
    .Z(net42));
 BUF_X1 input36 (.A(write_data[3]),
    .Z(net43));
 BUF_X1 input37 (.A(write_data[4]),
    .Z(net44));
 BUF_X1 input38 (.A(write_data[5]),
    .Z(net45));
 BUF_X1 input39 (.A(write_data[6]),
    .Z(net46));
 CLKBUF_X2 input40 (.A(write_data[7]),
    .Z(net47));
 BUF_X1 input41 (.A(write_data[8]),
    .Z(net48));
 BUF_X1 input42 (.A(write_data[9]),
    .Z(net49));
 BUF_X1 output43 (.A(net50),
    .Z(read_data[0]));
 BUF_X1 output44 (.A(net51),
    .Z(read_data[10]));
 BUF_X1 output45 (.A(net52),
    .Z(read_data[11]));
 BUF_X1 output46 (.A(net53),
    .Z(read_data[12]));
 BUF_X1 output47 (.A(net54),
    .Z(read_data[13]));
 BUF_X1 output48 (.A(net55),
    .Z(read_data[14]));
 BUF_X1 output49 (.A(net56),
    .Z(read_data[15]));
 BUF_X1 output50 (.A(net57),
    .Z(read_data[16]));
 BUF_X1 output51 (.A(net58),
    .Z(read_data[17]));
 BUF_X1 output52 (.A(net59),
    .Z(read_data[18]));
 BUF_X1 output53 (.A(net60),
    .Z(read_data[19]));
 BUF_X1 output54 (.A(net61),
    .Z(read_data[1]));
 BUF_X1 output55 (.A(net62),
    .Z(read_data[20]));
 BUF_X1 output56 (.A(net63),
    .Z(read_data[21]));
 BUF_X1 output57 (.A(net64),
    .Z(read_data[22]));
 BUF_X1 output58 (.A(net65),
    .Z(read_data[23]));
 BUF_X1 output59 (.A(net66),
    .Z(read_data[24]));
 BUF_X1 output60 (.A(net67),
    .Z(read_data[25]));
 BUF_X1 output61 (.A(net68),
    .Z(read_data[26]));
 BUF_X1 output62 (.A(net69),
    .Z(read_data[27]));
 BUF_X1 output63 (.A(net70),
    .Z(read_data[28]));
 BUF_X1 output64 (.A(net71),
    .Z(read_data[29]));
 BUF_X1 output65 (.A(net72),
    .Z(read_data[2]));
 BUF_X1 output66 (.A(net73),
    .Z(read_data[30]));
 BUF_X1 output67 (.A(net74),
    .Z(read_data[31]));
 BUF_X1 output68 (.A(net75),
    .Z(read_data[3]));
 BUF_X1 output69 (.A(net76),
    .Z(read_data[4]));
 BUF_X1 output70 (.A(net77),
    .Z(read_data[5]));
 BUF_X1 output71 (.A(net78),
    .Z(read_data[6]));
 BUF_X1 output72 (.A(net79),
    .Z(read_data[7]));
 BUF_X1 output73 (.A(net80),
    .Z(read_data[8]));
 BUF_X1 output74 (.A(net81),
    .Z(read_data[9]));
 BUF_X32 max_length75 (.A(net100),
    .Z(net82));
 BUF_X32 max_length76 (.A(net84),
    .Z(net83));
 BUF_X32 max_length77 (.A(net85),
    .Z(net84));
 BUF_X32 max_length78 (.A(net89),
    .Z(net85));
 BUF_X32 max_length79 (.A(net88),
    .Z(net86));
 BUF_X32 max_length80 (.A(net88),
    .Z(net87));
 BUF_X32 max_length81 (.A(net89),
    .Z(net88));
 BUF_X32 max_length82 (.A(net100),
    .Z(net89));
 BUF_X32 max_length83 (.A(net91),
    .Z(net90));
 BUF_X32 max_length84 (.A(net92),
    .Z(net91));
 BUF_X32 max_length85 (.A(net93),
    .Z(net92));
 BUF_X32 max_length86 (.A(net95),
    .Z(net93));
 BUF_X32 max_length87 (.A(net95),
    .Z(net94));
 BUF_X32 max_length88 (.A(net99),
    .Z(net95));
 BUF_X32 max_length89 (.A(net98),
    .Z(net96));
 BUF_X32 max_length90 (.A(net98),
    .Z(net97));
 BUF_X32 max_length91 (.A(net16),
    .Z(net98));
 BUF_X32 max_length92 (.A(net16),
    .Z(net99));
 BUF_X32 max_length93 (.A(net16),
    .Z(net100));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_leaf_80_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_80_clk));
 CLKBUF_X3 clkbuf_leaf_81_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_81_clk));
 CLKBUF_X3 clkbuf_leaf_82_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_82_clk));
 CLKBUF_X3 clkbuf_leaf_83_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_83_clk));
 CLKBUF_X3 clkbuf_leaf_84_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_84_clk));
 CLKBUF_X3 clkbuf_leaf_85_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_85_clk));
 CLKBUF_X3 clkbuf_leaf_86_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_86_clk));
 CLKBUF_X3 clkbuf_leaf_87_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_87_clk));
 CLKBUF_X3 clkbuf_leaf_88_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_88_clk));
 CLKBUF_X3 clkbuf_leaf_89_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_89_clk));
 CLKBUF_X3 clkbuf_leaf_90_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_90_clk));
 CLKBUF_X3 clkbuf_leaf_91_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_91_clk));
 CLKBUF_X3 clkbuf_leaf_92_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_92_clk));
 CLKBUF_X3 clkbuf_leaf_93_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_93_clk));
 CLKBUF_X3 clkbuf_leaf_94_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_94_clk));
 CLKBUF_X3 clkbuf_leaf_95_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_95_clk));
 CLKBUF_X3 clkbuf_leaf_96_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_96_clk));
 CLKBUF_X3 clkbuf_leaf_97_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_97_clk));
 CLKBUF_X3 clkbuf_leaf_98_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_98_clk));
 CLKBUF_X3 clkbuf_leaf_99_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_99_clk));
 CLKBUF_X3 clkbuf_leaf_100_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_100_clk));
 CLKBUF_X3 clkbuf_leaf_101_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_101_clk));
 CLKBUF_X3 clkbuf_leaf_102_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_102_clk));
 CLKBUF_X3 clkbuf_leaf_103_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_103_clk));
 CLKBUF_X3 clkbuf_leaf_104_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_104_clk));
 CLKBUF_X3 clkbuf_leaf_105_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_105_clk));
 CLKBUF_X3 clkbuf_leaf_106_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_106_clk));
 CLKBUF_X3 clkbuf_leaf_107_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_107_clk));
 CLKBUF_X3 clkbuf_leaf_108_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_108_clk));
 CLKBUF_X3 clkbuf_leaf_109_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_109_clk));
 CLKBUF_X3 clkbuf_leaf_110_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_110_clk));
 CLKBUF_X3 clkbuf_leaf_111_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_111_clk));
 CLKBUF_X3 clkbuf_leaf_112_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_112_clk));
 CLKBUF_X3 clkbuf_leaf_113_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_113_clk));
 CLKBUF_X3 clkbuf_leaf_114_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_114_clk));
 CLKBUF_X3 clkbuf_leaf_115_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_115_clk));
 CLKBUF_X3 clkbuf_leaf_116_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_116_clk));
 CLKBUF_X3 clkbuf_leaf_117_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_117_clk));
 CLKBUF_X3 clkbuf_leaf_118_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_118_clk));
 CLKBUF_X3 clkbuf_leaf_119_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_119_clk));
 CLKBUF_X3 clkbuf_leaf_120_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_120_clk));
 CLKBUF_X3 clkbuf_leaf_121_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_121_clk));
 CLKBUF_X3 clkbuf_leaf_122_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_122_clk));
 CLKBUF_X3 clkbuf_leaf_123_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_123_clk));
 CLKBUF_X3 clkbuf_leaf_124_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_124_clk));
 CLKBUF_X3 clkbuf_leaf_125_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_125_clk));
 CLKBUF_X3 clkbuf_leaf_126_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_126_clk));
 CLKBUF_X3 clkbuf_leaf_127_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_127_clk));
 CLKBUF_X3 clkbuf_leaf_128_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_128_clk));
 CLKBUF_X3 clkbuf_leaf_129_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_129_clk));
 CLKBUF_X3 clkbuf_leaf_130_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_130_clk));
 CLKBUF_X3 clkbuf_leaf_131_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_131_clk));
 CLKBUF_X3 clkbuf_leaf_132_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_132_clk));
 CLKBUF_X3 clkbuf_leaf_133_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_133_clk));
 CLKBUF_X3 clkbuf_leaf_134_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_134_clk));
 CLKBUF_X3 clkbuf_leaf_135_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_135_clk));
 CLKBUF_X3 clkbuf_leaf_136_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_136_clk));
 CLKBUF_X3 clkbuf_leaf_137_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_137_clk));
 CLKBUF_X3 clkbuf_leaf_138_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_138_clk));
 CLKBUF_X3 clkbuf_leaf_139_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_139_clk));
 CLKBUF_X3 clkbuf_leaf_140_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_140_clk));
 CLKBUF_X3 clkbuf_leaf_141_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_141_clk));
 CLKBUF_X3 clkbuf_leaf_142_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_142_clk));
 CLKBUF_X3 clkbuf_leaf_143_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_143_clk));
 CLKBUF_X3 clkbuf_leaf_144_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_144_clk));
 CLKBUF_X3 clkbuf_leaf_145_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_145_clk));
 CLKBUF_X3 clkbuf_leaf_146_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_146_clk));
 CLKBUF_X3 clkbuf_leaf_147_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_147_clk));
 CLKBUF_X3 clkbuf_leaf_148_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_148_clk));
 CLKBUF_X3 clkbuf_leaf_149_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_149_clk));
 CLKBUF_X3 clkbuf_leaf_150_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_150_clk));
 CLKBUF_X3 clkbuf_leaf_151_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_151_clk));
 CLKBUF_X3 clkbuf_leaf_152_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_152_clk));
 CLKBUF_X3 clkbuf_leaf_153_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_153_clk));
 CLKBUF_X3 clkbuf_leaf_154_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_154_clk));
 CLKBUF_X3 clkbuf_leaf_155_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_155_clk));
 CLKBUF_X3 clkbuf_leaf_156_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_156_clk));
 CLKBUF_X3 clkbuf_leaf_157_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_157_clk));
 CLKBUF_X3 clkbuf_leaf_158_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_158_clk));
 CLKBUF_X3 clkbuf_leaf_159_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_159_clk));
 CLKBUF_X3 clkbuf_leaf_160_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_160_clk));
 CLKBUF_X3 clkbuf_leaf_161_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_161_clk));
 CLKBUF_X3 clkbuf_leaf_162_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_162_clk));
 CLKBUF_X3 clkbuf_leaf_163_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_163_clk));
 CLKBUF_X3 clkbuf_leaf_164_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_164_clk));
 CLKBUF_X3 clkbuf_leaf_165_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_165_clk));
 CLKBUF_X3 clkbuf_leaf_166_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_166_clk));
 CLKBUF_X3 clkbuf_leaf_167_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_167_clk));
 CLKBUF_X3 clkbuf_leaf_168_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_168_clk));
 CLKBUF_X3 clkbuf_leaf_169_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_169_clk));
 CLKBUF_X3 clkbuf_leaf_170_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_170_clk));
 CLKBUF_X3 clkbuf_leaf_171_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_171_clk));
 CLKBUF_X3 clkbuf_leaf_172_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_172_clk));
 CLKBUF_X3 clkbuf_leaf_173_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_173_clk));
 CLKBUF_X3 clkbuf_leaf_174_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_174_clk));
 CLKBUF_X3 clkbuf_leaf_175_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_175_clk));
 CLKBUF_X3 clkbuf_leaf_176_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_176_clk));
 CLKBUF_X3 clkbuf_leaf_177_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_177_clk));
 CLKBUF_X3 clkbuf_leaf_178_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_178_clk));
 CLKBUF_X3 clkbuf_leaf_179_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_179_clk));
 CLKBUF_X3 clkbuf_leaf_180_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_180_clk));
 CLKBUF_X3 clkbuf_leaf_181_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_181_clk));
 CLKBUF_X3 clkbuf_leaf_182_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_182_clk));
 CLKBUF_X3 clkbuf_leaf_183_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_183_clk));
 CLKBUF_X3 clkbuf_leaf_184_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_184_clk));
 CLKBUF_X3 clkbuf_leaf_185_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_185_clk));
 CLKBUF_X3 clkbuf_leaf_186_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_186_clk));
 CLKBUF_X3 clkbuf_leaf_187_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_187_clk));
 CLKBUF_X3 clkbuf_leaf_188_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_188_clk));
 CLKBUF_X3 clkbuf_leaf_189_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_189_clk));
 CLKBUF_X3 clkbuf_leaf_190_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_190_clk));
 CLKBUF_X3 clkbuf_leaf_191_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_191_clk));
 CLKBUF_X3 clkbuf_leaf_192_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_192_clk));
 CLKBUF_X3 clkbuf_leaf_193_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_193_clk));
 CLKBUF_X3 clkbuf_leaf_194_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_194_clk));
 CLKBUF_X3 clkbuf_leaf_195_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_195_clk));
 CLKBUF_X3 clkbuf_leaf_196_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_196_clk));
 CLKBUF_X3 clkbuf_leaf_197_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_197_clk));
 CLKBUF_X3 clkbuf_leaf_198_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_198_clk));
 CLKBUF_X3 clkbuf_leaf_199_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_199_clk));
 CLKBUF_X3 clkbuf_leaf_200_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_200_clk));
 CLKBUF_X3 clkbuf_leaf_201_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_201_clk));
 CLKBUF_X3 clkbuf_leaf_202_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_202_clk));
 CLKBUF_X3 clkbuf_leaf_203_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_203_clk));
 CLKBUF_X3 clkbuf_leaf_204_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_204_clk));
 CLKBUF_X3 clkbuf_leaf_205_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_205_clk));
 CLKBUF_X3 clkbuf_leaf_206_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_206_clk));
 CLKBUF_X3 clkbuf_leaf_207_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_207_clk));
 CLKBUF_X3 clkbuf_leaf_208_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_208_clk));
 CLKBUF_X3 clkbuf_leaf_209_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_209_clk));
 CLKBUF_X3 clkbuf_leaf_210_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_210_clk));
 CLKBUF_X3 clkbuf_leaf_211_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_211_clk));
 CLKBUF_X3 clkbuf_leaf_212_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_212_clk));
 CLKBUF_X3 clkbuf_leaf_213_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_213_clk));
 CLKBUF_X3 clkbuf_leaf_214_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_214_clk));
 CLKBUF_X3 clkbuf_leaf_215_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_215_clk));
 CLKBUF_X3 clkbuf_leaf_216_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_216_clk));
 CLKBUF_X3 clkbuf_leaf_217_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_217_clk));
 CLKBUF_X3 clkbuf_leaf_218_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_218_clk));
 CLKBUF_X3 clkbuf_leaf_219_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_219_clk));
 CLKBUF_X3 clkbuf_leaf_220_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_220_clk));
 CLKBUF_X3 clkbuf_leaf_221_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_221_clk));
 CLKBUF_X3 clkbuf_leaf_222_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_222_clk));
 CLKBUF_X3 clkbuf_leaf_223_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_223_clk));
 CLKBUF_X3 clkbuf_leaf_224_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_224_clk));
 CLKBUF_X3 clkbuf_leaf_225_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_225_clk));
 CLKBUF_X3 clkbuf_leaf_226_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_226_clk));
 CLKBUF_X3 clkbuf_leaf_227_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_227_clk));
 CLKBUF_X3 clkbuf_leaf_228_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_228_clk));
 CLKBUF_X3 clkbuf_leaf_229_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_229_clk));
 CLKBUF_X3 clkbuf_leaf_230_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_230_clk));
 CLKBUF_X3 clkbuf_leaf_231_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_231_clk));
 CLKBUF_X3 clkbuf_leaf_232_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_232_clk));
 CLKBUF_X3 clkbuf_leaf_233_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_233_clk));
 CLKBUF_X3 clkbuf_leaf_234_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_234_clk));
 CLKBUF_X3 clkbuf_leaf_235_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_235_clk));
 CLKBUF_X3 clkbuf_leaf_236_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_236_clk));
 CLKBUF_X3 clkbuf_leaf_237_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_237_clk));
 CLKBUF_X3 clkbuf_leaf_238_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_238_clk));
 CLKBUF_X3 clkbuf_leaf_239_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_239_clk));
 CLKBUF_X3 clkbuf_leaf_240_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_240_clk));
 CLKBUF_X3 clkbuf_leaf_241_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_241_clk));
 CLKBUF_X3 clkbuf_leaf_242_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_242_clk));
 CLKBUF_X3 clkbuf_leaf_243_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_243_clk));
 CLKBUF_X3 clkbuf_leaf_244_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_244_clk));
 CLKBUF_X3 clkbuf_leaf_245_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_245_clk));
 CLKBUF_X3 clkbuf_leaf_246_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_246_clk));
 CLKBUF_X3 clkbuf_leaf_247_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_247_clk));
 CLKBUF_X3 clkbuf_leaf_248_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_248_clk));
 CLKBUF_X3 clkbuf_leaf_249_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_249_clk));
 CLKBUF_X3 clkbuf_leaf_250_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_250_clk));
 CLKBUF_X3 clkbuf_leaf_251_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_251_clk));
 CLKBUF_X3 clkbuf_leaf_252_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_252_clk));
 CLKBUF_X3 clkbuf_leaf_253_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_253_clk));
 CLKBUF_X3 clkbuf_leaf_254_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_254_clk));
 CLKBUF_X3 clkbuf_leaf_255_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_255_clk));
 CLKBUF_X3 clkbuf_leaf_256_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_256_clk));
 CLKBUF_X3 clkbuf_leaf_257_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_257_clk));
 CLKBUF_X3 clkbuf_leaf_258_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_258_clk));
 CLKBUF_X3 clkbuf_leaf_259_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_259_clk));
 CLKBUF_X3 clkbuf_leaf_260_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_260_clk));
 CLKBUF_X3 clkbuf_leaf_261_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_261_clk));
 CLKBUF_X3 clkbuf_leaf_262_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_262_clk));
 CLKBUF_X3 clkbuf_leaf_263_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_263_clk));
 CLKBUF_X3 clkbuf_leaf_264_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_264_clk));
 CLKBUF_X3 clkbuf_leaf_265_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_265_clk));
 CLKBUF_X3 clkbuf_leaf_266_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_266_clk));
 CLKBUF_X3 clkbuf_leaf_267_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_267_clk));
 CLKBUF_X3 clkbuf_leaf_268_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_268_clk));
 CLKBUF_X3 clkbuf_leaf_269_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_269_clk));
 CLKBUF_X3 clkbuf_leaf_270_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_270_clk));
 CLKBUF_X3 clkbuf_leaf_271_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_271_clk));
 CLKBUF_X3 clkbuf_leaf_272_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_272_clk));
 CLKBUF_X3 clkbuf_leaf_273_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_273_clk));
 CLKBUF_X3 clkbuf_leaf_274_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_274_clk));
 CLKBUF_X3 clkbuf_leaf_275_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_275_clk));
 CLKBUF_X3 clkbuf_leaf_276_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_276_clk));
 CLKBUF_X3 clkbuf_leaf_277_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_277_clk));
 CLKBUF_X3 clkbuf_leaf_278_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_278_clk));
 CLKBUF_X3 clkbuf_leaf_279_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_279_clk));
 CLKBUF_X3 clkbuf_leaf_280_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_280_clk));
 CLKBUF_X3 clkbuf_leaf_281_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_281_clk));
 CLKBUF_X3 clkbuf_leaf_282_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_282_clk));
 CLKBUF_X3 clkbuf_leaf_283_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_283_clk));
 CLKBUF_X3 clkbuf_leaf_284_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_284_clk));
 CLKBUF_X3 clkbuf_leaf_285_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_285_clk));
 CLKBUF_X3 clkbuf_leaf_286_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_286_clk));
 CLKBUF_X3 clkbuf_leaf_287_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_287_clk));
 CLKBUF_X3 clkbuf_leaf_288_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_288_clk));
 CLKBUF_X3 clkbuf_leaf_289_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_289_clk));
 CLKBUF_X3 clkbuf_leaf_290_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_290_clk));
 CLKBUF_X3 clkbuf_leaf_291_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_291_clk));
 CLKBUF_X3 clkbuf_leaf_292_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_292_clk));
 CLKBUF_X3 clkbuf_leaf_293_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_293_clk));
 CLKBUF_X3 clkbuf_leaf_294_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_294_clk));
 CLKBUF_X3 clkbuf_leaf_295_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_295_clk));
 CLKBUF_X3 clkbuf_leaf_296_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_296_clk));
 CLKBUF_X3 clkbuf_leaf_297_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_297_clk));
 CLKBUF_X3 clkbuf_leaf_298_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_298_clk));
 CLKBUF_X3 clkbuf_leaf_299_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_299_clk));
 CLKBUF_X3 clkbuf_leaf_300_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_300_clk));
 CLKBUF_X3 clkbuf_leaf_301_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_301_clk));
 CLKBUF_X3 clkbuf_leaf_302_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_302_clk));
 CLKBUF_X3 clkbuf_leaf_303_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_303_clk));
 CLKBUF_X3 clkbuf_leaf_304_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_304_clk));
 CLKBUF_X3 clkbuf_leaf_305_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_305_clk));
 CLKBUF_X3 clkbuf_leaf_306_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_306_clk));
 CLKBUF_X3 clkbuf_leaf_307_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_307_clk));
 CLKBUF_X3 clkbuf_leaf_308_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_308_clk));
 CLKBUF_X3 clkbuf_leaf_309_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_309_clk));
 CLKBUF_X3 clkbuf_leaf_310_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_310_clk));
 CLKBUF_X3 clkbuf_leaf_311_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_311_clk));
 CLKBUF_X3 clkbuf_leaf_312_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_312_clk));
 CLKBUF_X3 clkbuf_leaf_313_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_313_clk));
 CLKBUF_X3 clkbuf_leaf_314_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_314_clk));
 CLKBUF_X3 clkbuf_leaf_315_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_315_clk));
 CLKBUF_X3 clkbuf_leaf_316_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_316_clk));
 CLKBUF_X3 clkbuf_leaf_317_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_317_clk));
 CLKBUF_X3 clkbuf_leaf_318_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_318_clk));
 CLKBUF_X3 clkbuf_leaf_319_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_319_clk));
 CLKBUF_X3 clkbuf_leaf_320_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_320_clk));
 CLKBUF_X3 clkbuf_leaf_321_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_321_clk));
 CLKBUF_X3 clkbuf_leaf_322_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_322_clk));
 CLKBUF_X3 clkbuf_leaf_323_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_323_clk));
 CLKBUF_X3 clkbuf_leaf_324_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_324_clk));
 CLKBUF_X3 clkbuf_leaf_325_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_325_clk));
 CLKBUF_X3 clkbuf_leaf_326_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_326_clk));
 CLKBUF_X3 clkbuf_leaf_327_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_327_clk));
 CLKBUF_X3 clkbuf_leaf_328_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_328_clk));
 CLKBUF_X3 clkbuf_leaf_329_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_329_clk));
 CLKBUF_X3 clkbuf_leaf_330_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_330_clk));
 CLKBUF_X3 clkbuf_leaf_331_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_331_clk));
 CLKBUF_X3 clkbuf_leaf_332_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_332_clk));
 CLKBUF_X3 clkbuf_leaf_333_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_333_clk));
 CLKBUF_X3 clkbuf_leaf_334_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_334_clk));
 CLKBUF_X3 clkbuf_leaf_335_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_335_clk));
 CLKBUF_X3 clkbuf_leaf_336_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_336_clk));
 CLKBUF_X3 clkbuf_leaf_337_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_337_clk));
 CLKBUF_X3 clkbuf_leaf_338_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_338_clk));
 CLKBUF_X3 clkbuf_leaf_339_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_339_clk));
 CLKBUF_X3 clkbuf_leaf_340_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_340_clk));
 CLKBUF_X3 clkbuf_leaf_341_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_341_clk));
 CLKBUF_X3 clkbuf_leaf_342_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_342_clk));
 CLKBUF_X3 clkbuf_leaf_343_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_343_clk));
 CLKBUF_X3 clkbuf_leaf_344_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_344_clk));
 CLKBUF_X3 clkbuf_leaf_345_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_345_clk));
 CLKBUF_X3 clkbuf_leaf_346_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_346_clk));
 CLKBUF_X3 clkbuf_leaf_347_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_347_clk));
 CLKBUF_X3 clkbuf_leaf_348_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_348_clk));
 CLKBUF_X3 clkbuf_leaf_349_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_349_clk));
 CLKBUF_X3 clkbuf_leaf_350_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_350_clk));
 CLKBUF_X3 clkbuf_leaf_351_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_351_clk));
 CLKBUF_X3 clkbuf_leaf_352_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_352_clk));
 CLKBUF_X3 clkbuf_leaf_353_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_353_clk));
 CLKBUF_X3 clkbuf_leaf_354_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_354_clk));
 CLKBUF_X3 clkbuf_leaf_355_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_355_clk));
 CLKBUF_X3 clkbuf_leaf_356_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_356_clk));
 CLKBUF_X3 clkbuf_leaf_357_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_357_clk));
 CLKBUF_X3 clkbuf_leaf_358_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_358_clk));
 CLKBUF_X3 clkbuf_leaf_359_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_359_clk));
 CLKBUF_X3 clkbuf_leaf_360_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_360_clk));
 CLKBUF_X3 clkbuf_leaf_361_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_361_clk));
 CLKBUF_X3 clkbuf_leaf_362_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_362_clk));
 CLKBUF_X3 clkbuf_leaf_363_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_363_clk));
 CLKBUF_X3 clkbuf_leaf_364_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_364_clk));
 CLKBUF_X3 clkbuf_leaf_365_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_365_clk));
 CLKBUF_X3 clkbuf_leaf_366_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_366_clk));
 CLKBUF_X3 clkbuf_leaf_367_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_367_clk));
 CLKBUF_X3 clkbuf_leaf_368_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_368_clk));
 CLKBUF_X3 clkbuf_leaf_369_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_369_clk));
 CLKBUF_X3 clkbuf_leaf_370_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_370_clk));
 CLKBUF_X3 clkbuf_leaf_371_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_371_clk));
 CLKBUF_X3 clkbuf_leaf_372_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_372_clk));
 CLKBUF_X3 clkbuf_leaf_373_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_373_clk));
 CLKBUF_X3 clkbuf_leaf_374_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_374_clk));
 CLKBUF_X3 clkbuf_leaf_375_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_375_clk));
 CLKBUF_X3 clkbuf_leaf_376_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_376_clk));
 CLKBUF_X3 clkbuf_leaf_377_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_377_clk));
 CLKBUF_X3 clkbuf_leaf_378_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_378_clk));
 CLKBUF_X3 clkbuf_leaf_379_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_379_clk));
 CLKBUF_X3 clkbuf_leaf_380_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_380_clk));
 CLKBUF_X3 clkbuf_leaf_381_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_381_clk));
 CLKBUF_X3 clkbuf_leaf_382_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_382_clk));
 CLKBUF_X3 clkbuf_leaf_383_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_383_clk));
 CLKBUF_X3 clkbuf_leaf_384_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_384_clk));
 CLKBUF_X3 clkbuf_leaf_385_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_385_clk));
 CLKBUF_X3 clkbuf_leaf_386_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_386_clk));
 CLKBUF_X3 clkbuf_leaf_387_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_387_clk));
 CLKBUF_X3 clkbuf_leaf_388_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_388_clk));
 CLKBUF_X3 clkbuf_leaf_389_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_389_clk));
 CLKBUF_X3 clkbuf_leaf_390_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_390_clk));
 CLKBUF_X3 clkbuf_leaf_391_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_391_clk));
 CLKBUF_X3 clkbuf_leaf_392_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_392_clk));
 CLKBUF_X3 clkbuf_leaf_393_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_393_clk));
 CLKBUF_X3 clkbuf_leaf_394_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_394_clk));
 CLKBUF_X3 clkbuf_leaf_395_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_395_clk));
 CLKBUF_X3 clkbuf_leaf_396_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_396_clk));
 CLKBUF_X3 clkbuf_leaf_397_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_397_clk));
 CLKBUF_X3 clkbuf_leaf_398_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_398_clk));
 CLKBUF_X3 clkbuf_leaf_399_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_399_clk));
 CLKBUF_X3 clkbuf_leaf_400_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_400_clk));
 CLKBUF_X3 clkbuf_leaf_401_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_401_clk));
 CLKBUF_X3 clkbuf_leaf_402_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_402_clk));
 CLKBUF_X3 clkbuf_leaf_403_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_403_clk));
 CLKBUF_X3 clkbuf_leaf_404_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_404_clk));
 CLKBUF_X3 clkbuf_leaf_405_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_405_clk));
 CLKBUF_X3 clkbuf_leaf_406_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_406_clk));
 CLKBUF_X3 clkbuf_leaf_407_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_407_clk));
 CLKBUF_X3 clkbuf_leaf_408_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_408_clk));
 CLKBUF_X3 clkbuf_leaf_409_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_409_clk));
 CLKBUF_X3 clkbuf_leaf_410_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_410_clk));
 CLKBUF_X3 clkbuf_leaf_411_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_411_clk));
 CLKBUF_X3 clkbuf_leaf_412_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_412_clk));
 CLKBUF_X3 clkbuf_leaf_413_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_413_clk));
 CLKBUF_X3 clkbuf_leaf_414_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_414_clk));
 CLKBUF_X3 clkbuf_leaf_415_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_415_clk));
 CLKBUF_X3 clkbuf_leaf_416_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_416_clk));
 CLKBUF_X3 clkbuf_leaf_417_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_417_clk));
 CLKBUF_X3 clkbuf_leaf_418_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_418_clk));
 CLKBUF_X3 clkbuf_leaf_419_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_419_clk));
 CLKBUF_X3 clkbuf_leaf_420_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_420_clk));
 CLKBUF_X3 clkbuf_leaf_421_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_421_clk));
 CLKBUF_X3 clkbuf_leaf_422_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_422_clk));
 CLKBUF_X3 clkbuf_leaf_423_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_423_clk));
 CLKBUF_X3 clkbuf_leaf_424_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_424_clk));
 CLKBUF_X3 clkbuf_leaf_425_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_425_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_3_0_0_clk));
 CLKBUF_X3 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_3_1_0_clk));
 CLKBUF_X3 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_3_2_0_clk));
 CLKBUF_X3 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_3_3_0_clk));
 CLKBUF_X3 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_3_4_0_clk));
 CLKBUF_X3 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_3_5_0_clk));
 CLKBUF_X3 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_3_6_0_clk));
 CLKBUF_X3 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_3_7_0_clk));
 CLKBUF_X3 clkbuf_5_0__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_5_0__leaf_clk));
 CLKBUF_X3 clkbuf_5_1__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_5_1__leaf_clk));
 CLKBUF_X3 clkbuf_5_2__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_5_2__leaf_clk));
 CLKBUF_X3 clkbuf_5_3__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_5_3__leaf_clk));
 CLKBUF_X3 clkbuf_5_4__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_5_4__leaf_clk));
 CLKBUF_X3 clkbuf_5_5__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_5_5__leaf_clk));
 CLKBUF_X3 clkbuf_5_6__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_5_6__leaf_clk));
 CLKBUF_X3 clkbuf_5_7__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_5_7__leaf_clk));
 CLKBUF_X3 clkbuf_5_8__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_5_8__leaf_clk));
 CLKBUF_X3 clkbuf_5_9__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_5_9__leaf_clk));
 CLKBUF_X3 clkbuf_5_10__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_5_10__leaf_clk));
 CLKBUF_X3 clkbuf_5_11__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_5_11__leaf_clk));
 CLKBUF_X3 clkbuf_5_12__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_5_12__leaf_clk));
 CLKBUF_X3 clkbuf_5_13__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_5_13__leaf_clk));
 CLKBUF_X3 clkbuf_5_14__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_5_14__leaf_clk));
 CLKBUF_X3 clkbuf_5_15__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_5_15__leaf_clk));
 CLKBUF_X3 clkbuf_5_16__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_5_16__leaf_clk));
 CLKBUF_X3 clkbuf_5_17__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_5_17__leaf_clk));
 CLKBUF_X3 clkbuf_5_18__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_5_18__leaf_clk));
 CLKBUF_X3 clkbuf_5_19__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_5_19__leaf_clk));
 CLKBUF_X3 clkbuf_5_20__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_5_20__leaf_clk));
 CLKBUF_X3 clkbuf_5_21__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_5_21__leaf_clk));
 CLKBUF_X3 clkbuf_5_22__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_5_22__leaf_clk));
 CLKBUF_X3 clkbuf_5_23__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_5_23__leaf_clk));
 CLKBUF_X3 clkbuf_5_24__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_5_24__leaf_clk));
 CLKBUF_X3 clkbuf_5_25__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_5_25__leaf_clk));
 CLKBUF_X3 clkbuf_5_26__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_5_26__leaf_clk));
 CLKBUF_X3 clkbuf_5_27__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_5_27__leaf_clk));
 CLKBUF_X3 clkbuf_5_28__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_5_28__leaf_clk));
 CLKBUF_X3 clkbuf_5_29__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_5_29__leaf_clk));
 CLKBUF_X3 clkbuf_5_30__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_5_30__leaf_clk));
 CLKBUF_X3 clkbuf_5_31__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_5_31__leaf_clk));
 INV_X4 clkload0 (.A(clknet_5_0__leaf_clk));
 INV_X8 clkload1 (.A(clknet_5_1__leaf_clk));
 INV_X2 clkload2 (.A(clknet_5_4__leaf_clk));
 INV_X4 clkload3 (.A(clknet_5_5__leaf_clk));
 INV_X4 clkload4 (.A(clknet_5_6__leaf_clk));
 CLKBUF_X3 clkload5 (.A(clknet_5_9__leaf_clk));
 INV_X8 clkload6 (.A(clknet_5_10__leaf_clk));
 INV_X4 clkload7 (.A(clknet_5_11__leaf_clk));
 CLKBUF_X3 clkload8 (.A(clknet_5_12__leaf_clk));
 INV_X4 clkload9 (.A(clknet_5_14__leaf_clk));
 INV_X4 clkload10 (.A(clknet_5_15__leaf_clk));
 CLKBUF_X3 clkload11 (.A(clknet_5_16__leaf_clk));
 INV_X2 clkload12 (.A(clknet_5_17__leaf_clk));
 INV_X2 clkload13 (.A(clknet_5_19__leaf_clk));
 INV_X2 clkload14 (.A(clknet_5_20__leaf_clk));
 INV_X4 clkload15 (.A(clknet_5_22__leaf_clk));
 CLKBUF_X3 clkload16 (.A(clknet_5_23__leaf_clk));
 INV_X2 clkload17 (.A(clknet_5_24__leaf_clk));
 INV_X4 clkload18 (.A(clknet_5_25__leaf_clk));
 INV_X2 clkload19 (.A(clknet_5_27__leaf_clk));
 INV_X2 clkload20 (.A(clknet_5_29__leaf_clk));
 INV_X4 clkload21 (.A(clknet_5_30__leaf_clk));
 INV_X4 clkload22 (.A(clknet_5_31__leaf_clk));
 INV_X2 clkload23 (.A(clknet_leaf_0_clk));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_1_clk));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_2_clk));
 CLKBUF_X1 clkload26 (.A(clknet_leaf_10_clk));
 CLKBUF_X1 clkload27 (.A(clknet_leaf_11_clk));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_12_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_13_clk));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_14_clk));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_16_clk));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_24_clk));
 INV_X2 clkload33 (.A(clknet_leaf_425_clk));
 INV_X1 clkload34 (.A(clknet_leaf_4_clk));
 INV_X1 clkload35 (.A(clknet_leaf_5_clk));
 INV_X1 clkload36 (.A(clknet_leaf_8_clk));
 INV_X1 clkload37 (.A(clknet_leaf_9_clk));
 CLKBUF_X1 clkload38 (.A(clknet_leaf_32_clk));
 CLKBUF_X1 clkload39 (.A(clknet_leaf_34_clk));
 INV_X1 clkload40 (.A(clknet_leaf_35_clk));
 INV_X2 clkload41 (.A(clknet_leaf_419_clk));
 INV_X1 clkload42 (.A(clknet_leaf_423_clk));
 INV_X1 clkload43 (.A(clknet_leaf_424_clk));
 CLKBUF_X1 clkload44 (.A(clknet_leaf_17_clk));
 CLKBUF_X1 clkload45 (.A(clknet_leaf_18_clk));
 INV_X1 clkload46 (.A(clknet_leaf_22_clk));
 CLKBUF_X1 clkload47 (.A(clknet_leaf_23_clk));
 CLKBUF_X1 clkload48 (.A(clknet_leaf_94_clk));
 INV_X1 clkload49 (.A(clknet_leaf_95_clk));
 INV_X1 clkload50 (.A(clknet_leaf_97_clk));
 CLKBUF_X1 clkload51 (.A(clknet_leaf_98_clk));
 CLKBUF_X1 clkload52 (.A(clknet_leaf_100_clk));
 CLKBUF_X1 clkload53 (.A(clknet_leaf_101_clk));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_104_clk));
 INV_X1 clkload55 (.A(clknet_leaf_25_clk));
 INV_X2 clkload56 (.A(clknet_leaf_26_clk));
 CLKBUF_X1 clkload57 (.A(clknet_leaf_27_clk));
 CLKBUF_X1 clkload58 (.A(clknet_leaf_28_clk));
 INV_X1 clkload59 (.A(clknet_leaf_30_clk));
 CLKBUF_X1 clkload60 (.A(clknet_leaf_31_clk));
 INV_X1 clkload61 (.A(clknet_leaf_83_clk));
 INV_X1 clkload62 (.A(clknet_leaf_84_clk));
 CLKBUF_X1 clkload63 (.A(clknet_leaf_85_clk));
 INV_X2 clkload64 (.A(clknet_leaf_86_clk));
 CLKBUF_X1 clkload65 (.A(clknet_leaf_88_clk));
 INV_X1 clkload66 (.A(clknet_leaf_89_clk));
 CLKBUF_X1 clkload67 (.A(clknet_leaf_90_clk));
 INV_X1 clkload68 (.A(clknet_leaf_91_clk));
 INV_X1 clkload69 (.A(clknet_leaf_92_clk));
 CLKBUF_X1 clkload70 (.A(clknet_leaf_93_clk));
 INV_X2 clkload71 (.A(clknet_leaf_6_clk));
 INV_X1 clkload72 (.A(clknet_leaf_7_clk));
 CLKBUF_X1 clkload73 (.A(clknet_leaf_37_clk));
 INV_X1 clkload74 (.A(clknet_leaf_38_clk));
 INV_X2 clkload75 (.A(clknet_leaf_394_clk));
 CLKBUF_X1 clkload76 (.A(clknet_leaf_411_clk));
 CLKBUF_X1 clkload77 (.A(clknet_leaf_412_clk));
 INV_X1 clkload78 (.A(clknet_leaf_413_clk));
 CLKBUF_X1 clkload79 (.A(clknet_leaf_416_clk));
 CLKBUF_X1 clkload80 (.A(clknet_leaf_417_clk));
 INV_X1 clkload81 (.A(clknet_leaf_418_clk));
 INV_X1 clkload82 (.A(clknet_leaf_420_clk));
 CLKBUF_X1 clkload83 (.A(clknet_leaf_421_clk));
 INV_X1 clkload84 (.A(clknet_leaf_422_clk));
 INV_X2 clkload85 (.A(clknet_leaf_388_clk));
 INV_X1 clkload86 (.A(clknet_leaf_392_clk));
 CLKBUF_X1 clkload87 (.A(clknet_leaf_393_clk));
 INV_X1 clkload88 (.A(clknet_leaf_395_clk));
 INV_X1 clkload89 (.A(clknet_leaf_396_clk));
 INV_X1 clkload90 (.A(clknet_leaf_397_clk));
 INV_X1 clkload91 (.A(clknet_leaf_398_clk));
 INV_X2 clkload92 (.A(clknet_leaf_402_clk));
 CLKBUF_X1 clkload93 (.A(clknet_leaf_407_clk));
 INV_X1 clkload94 (.A(clknet_leaf_409_clk));
 CLKBUF_X1 clkload95 (.A(clknet_leaf_410_clk));
 CLKBUF_X1 clkload96 (.A(clknet_leaf_414_clk));
 INV_X2 clkload97 (.A(clknet_leaf_415_clk));
 CLKBUF_X1 clkload98 (.A(clknet_leaf_36_clk));
 CLKBUF_X1 clkload99 (.A(clknet_leaf_40_clk));
 INV_X1 clkload100 (.A(clknet_leaf_41_clk));
 INV_X1 clkload101 (.A(clknet_leaf_42_clk));
 CLKBUF_X1 clkload102 (.A(clknet_leaf_44_clk));
 CLKBUF_X1 clkload103 (.A(clknet_leaf_45_clk));
 CLKBUF_X1 clkload104 (.A(clknet_leaf_46_clk));
 CLKBUF_X1 clkload105 (.A(clknet_leaf_47_clk));
 CLKBUF_X1 clkload106 (.A(clknet_leaf_67_clk));
 CLKBUF_X1 clkload107 (.A(clknet_leaf_68_clk));
 INV_X1 clkload108 (.A(clknet_leaf_43_clk));
 INV_X1 clkload109 (.A(clknet_leaf_49_clk));
 CLKBUF_X1 clkload110 (.A(clknet_leaf_50_clk));
 INV_X1 clkload111 (.A(clknet_leaf_52_clk));
 INV_X1 clkload112 (.A(clknet_leaf_53_clk));
 CLKBUF_X1 clkload113 (.A(clknet_leaf_54_clk));
 INV_X2 clkload114 (.A(clknet_leaf_55_clk));
 CLKBUF_X1 clkload115 (.A(clknet_leaf_56_clk));
 CLKBUF_X1 clkload116 (.A(clknet_leaf_57_clk));
 INV_X1 clkload117 (.A(clknet_leaf_59_clk));
 INV_X1 clkload118 (.A(clknet_leaf_64_clk));
 CLKBUF_X1 clkload119 (.A(clknet_leaf_65_clk));
 CLKBUF_X1 clkload120 (.A(clknet_leaf_199_clk));
 CLKBUF_X1 clkload121 (.A(clknet_leaf_382_clk));
 CLKBUF_X1 clkload122 (.A(clknet_leaf_389_clk));
 INV_X1 clkload123 (.A(clknet_leaf_390_clk));
 CLKBUF_X1 clkload124 (.A(clknet_leaf_391_clk));
 CLKBUF_X1 clkload125 (.A(clknet_leaf_106_clk));
 CLKBUF_X1 clkload126 (.A(clknet_leaf_107_clk));
 CLKBUF_X1 clkload127 (.A(clknet_leaf_109_clk));
 CLKBUF_X1 clkload128 (.A(clknet_leaf_111_clk));
 INV_X1 clkload129 (.A(clknet_leaf_112_clk));
 INV_X1 clkload130 (.A(clknet_leaf_114_clk));
 CLKBUF_X1 clkload131 (.A(clknet_leaf_115_clk));
 CLKBUF_X1 clkload132 (.A(clknet_leaf_116_clk));
 CLKBUF_X1 clkload133 (.A(clknet_leaf_129_clk));
 INV_X2 clkload134 (.A(clknet_leaf_130_clk));
 CLKBUF_X1 clkload135 (.A(clknet_leaf_69_clk));
 INV_X1 clkload136 (.A(clknet_leaf_70_clk));
 INV_X2 clkload137 (.A(clknet_leaf_71_clk));
 CLKBUF_X1 clkload138 (.A(clknet_leaf_73_clk));
 CLKBUF_X1 clkload139 (.A(clknet_leaf_74_clk));
 CLKBUF_X1 clkload140 (.A(clknet_leaf_75_clk));
 CLKBUF_X1 clkload141 (.A(clknet_leaf_77_clk));
 CLKBUF_X1 clkload142 (.A(clknet_leaf_78_clk));
 CLKBUF_X1 clkload143 (.A(clknet_leaf_79_clk));
 CLKBUF_X1 clkload144 (.A(clknet_leaf_80_clk));
 CLKBUF_X1 clkload145 (.A(clknet_leaf_81_clk));
 CLKBUF_X1 clkload146 (.A(clknet_leaf_117_clk));
 CLKBUF_X1 clkload147 (.A(clknet_leaf_118_clk));
 CLKBUF_X1 clkload148 (.A(clknet_leaf_121_clk));
 INV_X1 clkload149 (.A(clknet_leaf_120_clk));
 INV_X1 clkload150 (.A(clknet_leaf_124_clk));
 INV_X1 clkload151 (.A(clknet_leaf_125_clk));
 INV_X2 clkload152 (.A(clknet_leaf_131_clk));
 INV_X1 clkload153 (.A(clknet_leaf_135_clk));
 INV_X1 clkload154 (.A(clknet_leaf_136_clk));
 CLKBUF_X1 clkload155 (.A(clknet_leaf_137_clk));
 CLKBUF_X1 clkload156 (.A(clknet_leaf_138_clk));
 CLKBUF_X1 clkload157 (.A(clknet_leaf_140_clk));
 INV_X1 clkload158 (.A(clknet_leaf_132_clk));
 INV_X1 clkload159 (.A(clknet_leaf_139_clk));
 INV_X1 clkload160 (.A(clknet_leaf_141_clk));
 INV_X1 clkload161 (.A(clknet_leaf_142_clk));
 INV_X1 clkload162 (.A(clknet_leaf_143_clk));
 CLKBUF_X1 clkload163 (.A(clknet_leaf_144_clk));
 INV_X2 clkload164 (.A(clknet_leaf_145_clk));
 INV_X2 clkload165 (.A(clknet_leaf_148_clk));
 CLKBUF_X1 clkload166 (.A(clknet_leaf_149_clk));
 INV_X2 clkload167 (.A(clknet_leaf_151_clk));
 INV_X1 clkload168 (.A(clknet_leaf_176_clk));
 INV_X1 clkload169 (.A(clknet_leaf_177_clk));
 CLKBUF_X1 clkload170 (.A(clknet_leaf_60_clk));
 INV_X1 clkload171 (.A(clknet_leaf_61_clk));
 CLKBUF_X1 clkload172 (.A(clknet_leaf_62_clk));
 CLKBUF_X1 clkload173 (.A(clknet_leaf_63_clk));
 INV_X2 clkload174 (.A(clknet_leaf_72_clk));
 INV_X1 clkload175 (.A(clknet_leaf_179_clk));
 INV_X1 clkload176 (.A(clknet_leaf_180_clk));
 CLKBUF_X1 clkload177 (.A(clknet_leaf_181_clk));
 INV_X1 clkload178 (.A(clknet_leaf_182_clk));
 INV_X1 clkload179 (.A(clknet_leaf_183_clk));
 INV_X1 clkload180 (.A(clknet_leaf_184_clk));
 INV_X1 clkload181 (.A(clknet_leaf_185_clk));
 INV_X1 clkload182 (.A(clknet_leaf_186_clk));
 INV_X1 clkload183 (.A(clknet_leaf_187_clk));
 CLKBUF_X1 clkload184 (.A(clknet_leaf_193_clk));
 INV_X1 clkload185 (.A(clknet_leaf_194_clk));
 INV_X1 clkload186 (.A(clknet_leaf_195_clk));
 CLKBUF_X1 clkload187 (.A(clknet_leaf_188_clk));
 CLKBUF_X1 clkload188 (.A(clknet_leaf_189_clk));
 CLKBUF_X1 clkload189 (.A(clknet_leaf_191_clk));
 INV_X1 clkload190 (.A(clknet_leaf_196_clk));
 CLKBUF_X1 clkload191 (.A(clknet_leaf_200_clk));
 CLKBUF_X1 clkload192 (.A(clknet_leaf_201_clk));
 INV_X1 clkload193 (.A(clknet_leaf_202_clk));
 CLKBUF_X1 clkload194 (.A(clknet_leaf_206_clk));
 INV_X1 clkload195 (.A(clknet_leaf_207_clk));
 INV_X1 clkload196 (.A(clknet_leaf_208_clk));
 CLKBUF_X1 clkload197 (.A(clknet_leaf_209_clk));
 CLKBUF_X1 clkload198 (.A(clknet_leaf_210_clk));
 INV_X1 clkload199 (.A(clknet_leaf_146_clk));
 INV_X1 clkload200 (.A(clknet_leaf_147_clk));
 INV_X1 clkload201 (.A(clknet_leaf_152_clk));
 INV_X1 clkload202 (.A(clknet_leaf_153_clk));
 INV_X1 clkload203 (.A(clknet_leaf_154_clk));
 CLKBUF_X1 clkload204 (.A(clknet_leaf_155_clk));
 INV_X1 clkload205 (.A(clknet_leaf_156_clk));
 CLKBUF_X1 clkload206 (.A(clknet_leaf_157_clk));
 INV_X1 clkload207 (.A(clknet_leaf_164_clk));
 INV_X1 clkload208 (.A(clknet_leaf_170_clk));
 INV_X1 clkload209 (.A(clknet_leaf_171_clk));
 CLKBUF_X1 clkload210 (.A(clknet_leaf_172_clk));
 INV_X1 clkload211 (.A(clknet_leaf_174_clk));
 CLKBUF_X1 clkload212 (.A(clknet_leaf_175_clk));
 INV_X2 clkload213 (.A(clknet_leaf_158_clk));
 CLKBUF_X1 clkload214 (.A(clknet_leaf_159_clk));
 CLKBUF_X1 clkload215 (.A(clknet_leaf_160_clk));
 INV_X1 clkload216 (.A(clknet_leaf_161_clk));
 INV_X1 clkload217 (.A(clknet_leaf_162_clk));
 INV_X1 clkload218 (.A(clknet_leaf_163_clk));
 INV_X2 clkload219 (.A(clknet_leaf_165_clk));
 INV_X1 clkload220 (.A(clknet_leaf_168_clk));
 CLKBUF_X1 clkload221 (.A(clknet_leaf_229_clk));
 INV_X1 clkload222 (.A(clknet_leaf_230_clk));
 INV_X1 clkload223 (.A(clknet_leaf_231_clk));
 INV_X2 clkload224 (.A(clknet_leaf_236_clk));
 INV_X1 clkload225 (.A(clknet_leaf_237_clk));
 CLKBUF_X1 clkload226 (.A(clknet_leaf_346_clk));
 CLKBUF_X1 clkload227 (.A(clknet_leaf_347_clk));
 INV_X1 clkload228 (.A(clknet_leaf_350_clk));
 INV_X1 clkload229 (.A(clknet_leaf_351_clk));
 CLKBUF_X1 clkload230 (.A(clknet_leaf_353_clk));
 CLKBUF_X1 clkload231 (.A(clknet_leaf_399_clk));
 INV_X1 clkload232 (.A(clknet_leaf_400_clk));
 INV_X2 clkload233 (.A(clknet_leaf_401_clk));
 CLKBUF_X1 clkload234 (.A(clknet_leaf_403_clk));
 CLKBUF_X1 clkload235 (.A(clknet_leaf_404_clk));
 CLKBUF_X1 clkload236 (.A(clknet_leaf_405_clk));
 INV_X1 clkload237 (.A(clknet_leaf_406_clk));
 CLKBUF_X1 clkload238 (.A(clknet_leaf_339_clk));
 CLKBUF_X1 clkload239 (.A(clknet_leaf_340_clk));
 CLKBUF_X1 clkload240 (.A(clknet_leaf_343_clk));
 CLKBUF_X1 clkload241 (.A(clknet_leaf_344_clk));
 CLKBUF_X1 clkload242 (.A(clknet_leaf_345_clk));
 CLKBUF_X1 clkload243 (.A(clknet_leaf_349_clk));
 CLKBUF_X1 clkload244 (.A(clknet_leaf_356_clk));
 CLKBUF_X1 clkload245 (.A(clknet_leaf_357_clk));
 CLKBUF_X1 clkload246 (.A(clknet_leaf_358_clk));
 INV_X1 clkload247 (.A(clknet_leaf_359_clk));
 INV_X2 clkload248 (.A(clknet_leaf_352_clk));
 CLKBUF_X1 clkload249 (.A(clknet_leaf_367_clk));
 INV_X1 clkload250 (.A(clknet_leaf_368_clk));
 INV_X1 clkload251 (.A(clknet_leaf_369_clk));
 INV_X1 clkload252 (.A(clknet_leaf_370_clk));
 INV_X1 clkload253 (.A(clknet_leaf_374_clk));
 INV_X1 clkload254 (.A(clknet_leaf_375_clk));
 INV_X2 clkload255 (.A(clknet_leaf_380_clk));
 INV_X1 clkload256 (.A(clknet_leaf_381_clk));
 CLKBUF_X1 clkload257 (.A(clknet_leaf_384_clk));
 INV_X2 clkload258 (.A(clknet_leaf_385_clk));
 INV_X2 clkload259 (.A(clknet_leaf_386_clk));
 INV_X2 clkload260 (.A(clknet_leaf_387_clk));
 CLKBUF_X1 clkload261 (.A(clknet_leaf_286_clk));
 INV_X1 clkload262 (.A(clknet_leaf_292_clk));
 INV_X2 clkload263 (.A(clknet_leaf_360_clk));
 CLKBUF_X1 clkload264 (.A(clknet_leaf_361_clk));
 CLKBUF_X1 clkload265 (.A(clknet_leaf_362_clk));
 CLKBUF_X1 clkload266 (.A(clknet_leaf_365_clk));
 CLKBUF_X1 clkload267 (.A(clknet_leaf_366_clk));
 CLKBUF_X1 clkload268 (.A(clknet_leaf_372_clk));
 CLKBUF_X1 clkload269 (.A(clknet_leaf_373_clk));
 CLKBUF_X1 clkload270 (.A(clknet_leaf_332_clk));
 INV_X2 clkload271 (.A(clknet_leaf_333_clk));
 INV_X1 clkload272 (.A(clknet_leaf_334_clk));
 CLKBUF_X1 clkload273 (.A(clknet_leaf_335_clk));
 INV_X2 clkload274 (.A(clknet_leaf_336_clk));
 CLKBUF_X1 clkload275 (.A(clknet_leaf_337_clk));
 INV_X1 clkload276 (.A(clknet_leaf_338_clk));
 INV_X1 clkload277 (.A(clknet_leaf_341_clk));
 CLKBUF_X1 clkload278 (.A(clknet_leaf_342_clk));
 INV_X1 clkload279 (.A(clknet_leaf_314_clk));
 CLKBUF_X1 clkload280 (.A(clknet_leaf_315_clk));
 INV_X2 clkload281 (.A(clknet_leaf_316_clk));
 CLKBUF_X1 clkload282 (.A(clknet_leaf_321_clk));
 CLKBUF_X1 clkload283 (.A(clknet_leaf_324_clk));
 INV_X1 clkload284 (.A(clknet_leaf_325_clk));
 CLKBUF_X1 clkload285 (.A(clknet_leaf_326_clk));
 CLKBUF_X1 clkload286 (.A(clknet_leaf_327_clk));
 INV_X1 clkload287 (.A(clknet_leaf_329_clk));
 INV_X2 clkload288 (.A(clknet_leaf_293_clk));
 CLKBUF_X1 clkload289 (.A(clknet_leaf_294_clk));
 INV_X1 clkload290 (.A(clknet_leaf_295_clk));
 INV_X2 clkload291 (.A(clknet_leaf_296_clk));
 INV_X1 clkload292 (.A(clknet_leaf_300_clk));
 INV_X1 clkload293 (.A(clknet_leaf_312_clk));
 INV_X1 clkload294 (.A(clknet_leaf_313_clk));
 CLKBUF_X1 clkload295 (.A(clknet_leaf_301_clk));
 INV_X1 clkload296 (.A(clknet_leaf_304_clk));
 CLKBUF_X1 clkload297 (.A(clknet_leaf_305_clk));
 CLKBUF_X1 clkload298 (.A(clknet_leaf_306_clk));
 INV_X1 clkload299 (.A(clknet_leaf_307_clk));
 INV_X1 clkload300 (.A(clknet_leaf_308_clk));
 INV_X1 clkload301 (.A(clknet_leaf_309_clk));
 INV_X1 clkload302 (.A(clknet_leaf_310_clk));
 CLKBUF_X1 clkload303 (.A(clknet_leaf_319_clk));
 CLKBUF_X1 clkload304 (.A(clknet_leaf_320_clk));
 CLKBUF_X1 clkload305 (.A(clknet_leaf_205_clk));
 CLKBUF_X1 clkload306 (.A(clknet_leaf_281_clk));
 CLKBUF_X1 clkload307 (.A(clknet_leaf_283_clk));
 CLKBUF_X1 clkload308 (.A(clknet_leaf_376_clk));
 CLKBUF_X1 clkload309 (.A(clknet_leaf_377_clk));
 CLKBUF_X1 clkload310 (.A(clknet_leaf_378_clk));
 CLKBUF_X1 clkload311 (.A(clknet_leaf_379_clk));
 CLKBUF_X1 clkload312 (.A(clknet_leaf_215_clk));
 CLKBUF_X1 clkload313 (.A(clknet_leaf_216_clk));
 CLKBUF_X1 clkload314 (.A(clknet_leaf_284_clk));
 CLKBUF_X1 clkload315 (.A(clknet_leaf_285_clk));
 CLKBUF_X1 clkload316 (.A(clknet_leaf_213_clk));
 CLKBUF_X1 clkload317 (.A(clknet_leaf_224_clk));
 INV_X1 clkload318 (.A(clknet_leaf_225_clk));
 CLKBUF_X1 clkload319 (.A(clknet_leaf_226_clk));
 CLKBUF_X1 clkload320 (.A(clknet_leaf_227_clk));
 CLKBUF_X1 clkload321 (.A(clknet_leaf_228_clk));
 CLKBUF_X1 clkload322 (.A(clknet_leaf_232_clk));
 INV_X1 clkload323 (.A(clknet_leaf_233_clk));
 CLKBUF_X1 clkload324 (.A(clknet_leaf_234_clk));
 INV_X1 clkload325 (.A(clknet_leaf_235_clk));
 CLKBUF_X1 clkload326 (.A(clknet_leaf_240_clk));
 INV_X1 clkload327 (.A(clknet_leaf_241_clk));
 INV_X1 clkload328 (.A(clknet_leaf_243_clk));
 INV_X1 clkload329 (.A(clknet_leaf_218_clk));
 INV_X1 clkload330 (.A(clknet_leaf_219_clk));
 CLKBUF_X1 clkload331 (.A(clknet_leaf_220_clk));
 INV_X1 clkload332 (.A(clknet_leaf_221_clk));
 CLKBUF_X1 clkload333 (.A(clknet_leaf_222_clk));
 INV_X2 clkload334 (.A(clknet_leaf_223_clk));
 INV_X2 clkload335 (.A(clknet_leaf_244_clk));
 CLKBUF_X1 clkload336 (.A(clknet_leaf_245_clk));
 INV_X1 clkload337 (.A(clknet_leaf_246_clk));
 CLKBUF_X1 clkload338 (.A(clknet_leaf_247_clk));
 CLKBUF_X1 clkload339 (.A(clknet_leaf_262_clk));
 CLKBUF_X1 clkload340 (.A(clknet_leaf_269_clk));
 INV_X1 clkload341 (.A(clknet_leaf_270_clk));
 INV_X1 clkload342 (.A(clknet_leaf_271_clk));
 CLKBUF_X1 clkload343 (.A(clknet_leaf_272_clk));
 CLKBUF_X1 clkload344 (.A(clknet_leaf_273_clk));
 INV_X1 clkload345 (.A(clknet_leaf_274_clk));
 CLKBUF_X1 clkload346 (.A(clknet_leaf_275_clk));
 INV_X1 clkload347 (.A(clknet_leaf_276_clk));
 CLKBUF_X1 clkload348 (.A(clknet_leaf_288_clk));
 INV_X1 clkload349 (.A(clknet_leaf_289_clk));
 INV_X1 clkload350 (.A(clknet_leaf_290_clk));
 INV_X2 clkload351 (.A(clknet_leaf_291_clk));
 CLKBUF_X1 clkload352 (.A(clknet_leaf_253_clk));
 CLKBUF_X1 clkload353 (.A(clknet_leaf_254_clk));
 INV_X1 clkload354 (.A(clknet_leaf_256_clk));
 CLKBUF_X1 clkload355 (.A(clknet_leaf_257_clk));
 CLKBUF_X1 clkload356 (.A(clknet_leaf_297_clk));
 CLKBUF_X1 clkload357 (.A(clknet_leaf_298_clk));
 CLKBUF_X1 clkload358 (.A(clknet_leaf_299_clk));
 CLKBUF_X1 clkload359 (.A(clknet_leaf_302_clk));
 CLKBUF_X1 clkload360 (.A(clknet_leaf_303_clk));
 INV_X4 clkload361 (.A(clknet_leaf_251_clk));
 INV_X1 clkload362 (.A(clknet_leaf_252_clk));
 INV_X2 clkload363 (.A(clknet_leaf_258_clk));
 CLKBUF_X1 clkload364 (.A(clknet_leaf_259_clk));
 INV_X1 clkload365 (.A(clknet_leaf_261_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X4 FILLER_0_225 ();
 FILLCELL_X16 FILLER_0_233 ();
 FILLCELL_X8 FILLER_0_249 ();
 FILLCELL_X4 FILLER_0_257 ();
 FILLCELL_X2 FILLER_0_261 ();
 FILLCELL_X16 FILLER_0_287 ();
 FILLCELL_X8 FILLER_0_303 ();
 FILLCELL_X2 FILLER_0_311 ();
 FILLCELL_X16 FILLER_0_322 ();
 FILLCELL_X8 FILLER_0_338 ();
 FILLCELL_X4 FILLER_0_346 ();
 FILLCELL_X1 FILLER_0_350 ();
 FILLCELL_X32 FILLER_0_360 ();
 FILLCELL_X16 FILLER_0_392 ();
 FILLCELL_X4 FILLER_0_408 ();
 FILLCELL_X1 FILLER_0_412 ();
 FILLCELL_X8 FILLER_0_417 ();
 FILLCELL_X2 FILLER_0_425 ();
 FILLCELL_X32 FILLER_0_431 ();
 FILLCELL_X2 FILLER_0_463 ();
 FILLCELL_X32 FILLER_0_469 ();
 FILLCELL_X16 FILLER_0_501 ();
 FILLCELL_X2 FILLER_0_517 ();
 FILLCELL_X1 FILLER_0_519 ();
 FILLCELL_X8 FILLER_0_523 ();
 FILLCELL_X4 FILLER_0_531 ();
 FILLCELL_X32 FILLER_0_538 ();
 FILLCELL_X32 FILLER_0_570 ();
 FILLCELL_X16 FILLER_0_602 ();
 FILLCELL_X8 FILLER_0_618 ();
 FILLCELL_X4 FILLER_0_626 ();
 FILLCELL_X1 FILLER_0_630 ();
 FILLCELL_X1 FILLER_0_632 ();
 FILLCELL_X4 FILLER_0_637 ();
 FILLCELL_X4 FILLER_0_649 ();
 FILLCELL_X1 FILLER_0_653 ();
 FILLCELL_X8 FILLER_0_658 ();
 FILLCELL_X2 FILLER_0_666 ();
 FILLCELL_X1 FILLER_0_668 ();
 FILLCELL_X8 FILLER_0_673 ();
 FILLCELL_X2 FILLER_0_681 ();
 FILLCELL_X1 FILLER_0_683 ();
 FILLCELL_X2 FILLER_0_688 ();
 FILLCELL_X8 FILLER_0_694 ();
 FILLCELL_X2 FILLER_0_702 ();
 FILLCELL_X32 FILLER_0_708 ();
 FILLCELL_X32 FILLER_0_740 ();
 FILLCELL_X16 FILLER_0_772 ();
 FILLCELL_X4 FILLER_0_788 ();
 FILLCELL_X2 FILLER_0_792 ();
 FILLCELL_X1 FILLER_0_794 ();
 FILLCELL_X32 FILLER_0_800 ();
 FILLCELL_X32 FILLER_0_832 ();
 FILLCELL_X32 FILLER_0_864 ();
 FILLCELL_X16 FILLER_0_896 ();
 FILLCELL_X8 FILLER_0_912 ();
 FILLCELL_X2 FILLER_0_920 ();
 FILLCELL_X32 FILLER_0_929 ();
 FILLCELL_X32 FILLER_0_961 ();
 FILLCELL_X32 FILLER_0_993 ();
 FILLCELL_X32 FILLER_0_1025 ();
 FILLCELL_X32 FILLER_0_1057 ();
 FILLCELL_X32 FILLER_0_1089 ();
 FILLCELL_X32 FILLER_0_1121 ();
 FILLCELL_X32 FILLER_0_1153 ();
 FILLCELL_X32 FILLER_0_1185 ();
 FILLCELL_X32 FILLER_0_1217 ();
 FILLCELL_X8 FILLER_0_1249 ();
 FILLCELL_X4 FILLER_0_1257 ();
 FILLCELL_X1 FILLER_0_1261 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X32 FILLER_0_1295 ();
 FILLCELL_X32 FILLER_0_1327 ();
 FILLCELL_X32 FILLER_0_1359 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X32 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1487 ();
 FILLCELL_X32 FILLER_0_1519 ();
 FILLCELL_X32 FILLER_0_1551 ();
 FILLCELL_X32 FILLER_0_1583 ();
 FILLCELL_X32 FILLER_0_1615 ();
 FILLCELL_X4 FILLER_0_1647 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X1 FILLER_1_257 ();
 FILLCELL_X16 FILLER_1_278 ();
 FILLCELL_X1 FILLER_1_294 ();
 FILLCELL_X1 FILLER_1_298 ();
 FILLCELL_X2 FILLER_1_316 ();
 FILLCELL_X8 FILLER_1_330 ();
 FILLCELL_X4 FILLER_1_338 ();
 FILLCELL_X1 FILLER_1_342 ();
 FILLCELL_X4 FILLER_1_352 ();
 FILLCELL_X2 FILLER_1_356 ();
 FILLCELL_X1 FILLER_1_358 ();
 FILLCELL_X32 FILLER_1_368 ();
 FILLCELL_X32 FILLER_1_400 ();
 FILLCELL_X16 FILLER_1_432 ();
 FILLCELL_X8 FILLER_1_448 ();
 FILLCELL_X2 FILLER_1_456 ();
 FILLCELL_X1 FILLER_1_458 ();
 FILLCELL_X2 FILLER_1_466 ();
 FILLCELL_X2 FILLER_1_475 ();
 FILLCELL_X1 FILLER_1_477 ();
 FILLCELL_X1 FILLER_1_485 ();
 FILLCELL_X2 FILLER_1_489 ();
 FILLCELL_X1 FILLER_1_491 ();
 FILLCELL_X4 FILLER_1_509 ();
 FILLCELL_X2 FILLER_1_513 ();
 FILLCELL_X1 FILLER_1_519 ();
 FILLCELL_X1 FILLER_1_527 ();
 FILLCELL_X1 FILLER_1_531 ();
 FILLCELL_X2 FILLER_1_556 ();
 FILLCELL_X2 FILLER_1_563 ();
 FILLCELL_X1 FILLER_1_565 ();
 FILLCELL_X4 FILLER_1_573 ();
 FILLCELL_X1 FILLER_1_577 ();
 FILLCELL_X1 FILLER_1_587 ();
 FILLCELL_X1 FILLER_1_602 ();
 FILLCELL_X1 FILLER_1_610 ();
 FILLCELL_X8 FILLER_1_618 ();
 FILLCELL_X4 FILLER_1_626 ();
 FILLCELL_X2 FILLER_1_630 ();
 FILLCELL_X16 FILLER_1_639 ();
 FILLCELL_X2 FILLER_1_655 ();
 FILLCELL_X32 FILLER_1_664 ();
 FILLCELL_X32 FILLER_1_696 ();
 FILLCELL_X16 FILLER_1_728 ();
 FILLCELL_X2 FILLER_1_744 ();
 FILLCELL_X1 FILLER_1_746 ();
 FILLCELL_X8 FILLER_1_754 ();
 FILLCELL_X1 FILLER_1_762 ();
 FILLCELL_X2 FILLER_1_767 ();
 FILLCELL_X4 FILLER_1_778 ();
 FILLCELL_X4 FILLER_1_789 ();
 FILLCELL_X4 FILLER_1_800 ();
 FILLCELL_X16 FILLER_1_815 ();
 FILLCELL_X8 FILLER_1_831 ();
 FILLCELL_X8 FILLER_1_843 ();
 FILLCELL_X2 FILLER_1_851 ();
 FILLCELL_X1 FILLER_1_853 ();
 FILLCELL_X4 FILLER_1_858 ();
 FILLCELL_X2 FILLER_1_862 ();
 FILLCELL_X1 FILLER_1_864 ();
 FILLCELL_X4 FILLER_1_872 ();
 FILLCELL_X16 FILLER_1_883 ();
 FILLCELL_X4 FILLER_1_899 ();
 FILLCELL_X2 FILLER_1_903 ();
 FILLCELL_X1 FILLER_1_905 ();
 FILLCELL_X8 FILLER_1_913 ();
 FILLCELL_X4 FILLER_1_921 ();
 FILLCELL_X2 FILLER_1_925 ();
 FILLCELL_X1 FILLER_1_927 ();
 FILLCELL_X32 FILLER_1_935 ();
 FILLCELL_X32 FILLER_1_967 ();
 FILLCELL_X32 FILLER_1_999 ();
 FILLCELL_X32 FILLER_1_1031 ();
 FILLCELL_X16 FILLER_1_1063 ();
 FILLCELL_X4 FILLER_1_1079 ();
 FILLCELL_X1 FILLER_1_1083 ();
 FILLCELL_X4 FILLER_1_1091 ();
 FILLCELL_X2 FILLER_1_1095 ();
 FILLCELL_X1 FILLER_1_1097 ();
 FILLCELL_X4 FILLER_1_1105 ();
 FILLCELL_X2 FILLER_1_1109 ();
 FILLCELL_X16 FILLER_1_1114 ();
 FILLCELL_X8 FILLER_1_1137 ();
 FILLCELL_X2 FILLER_1_1145 ();
 FILLCELL_X1 FILLER_1_1147 ();
 FILLCELL_X4 FILLER_1_1159 ();
 FILLCELL_X2 FILLER_1_1163 ();
 FILLCELL_X8 FILLER_1_1175 ();
 FILLCELL_X4 FILLER_1_1183 ();
 FILLCELL_X1 FILLER_1_1187 ();
 FILLCELL_X32 FILLER_1_1229 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X32 FILLER_1_1424 ();
 FILLCELL_X32 FILLER_1_1456 ();
 FILLCELL_X32 FILLER_1_1488 ();
 FILLCELL_X32 FILLER_1_1520 ();
 FILLCELL_X32 FILLER_1_1552 ();
 FILLCELL_X32 FILLER_1_1584 ();
 FILLCELL_X32 FILLER_1_1616 ();
 FILLCELL_X2 FILLER_1_1648 ();
 FILLCELL_X1 FILLER_1_1650 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X8 FILLER_2_225 ();
 FILLCELL_X4 FILLER_2_233 ();
 FILLCELL_X4 FILLER_2_241 ();
 FILLCELL_X2 FILLER_2_245 ();
 FILLCELL_X4 FILLER_2_268 ();
 FILLCELL_X4 FILLER_2_279 ();
 FILLCELL_X2 FILLER_2_283 ();
 FILLCELL_X1 FILLER_2_305 ();
 FILLCELL_X4 FILLER_2_313 ();
 FILLCELL_X2 FILLER_2_317 ();
 FILLCELL_X8 FILLER_2_360 ();
 FILLCELL_X2 FILLER_2_368 ();
 FILLCELL_X1 FILLER_2_370 ();
 FILLCELL_X8 FILLER_2_378 ();
 FILLCELL_X4 FILLER_2_386 ();
 FILLCELL_X32 FILLER_2_397 ();
 FILLCELL_X16 FILLER_2_429 ();
 FILLCELL_X8 FILLER_2_445 ();
 FILLCELL_X4 FILLER_2_453 ();
 FILLCELL_X2 FILLER_2_457 ();
 FILLCELL_X2 FILLER_2_479 ();
 FILLCELL_X4 FILLER_2_512 ();
 FILLCELL_X1 FILLER_2_516 ();
 FILLCELL_X2 FILLER_2_525 ();
 FILLCELL_X1 FILLER_2_527 ();
 FILLCELL_X4 FILLER_2_535 ();
 FILLCELL_X2 FILLER_2_539 ();
 FILLCELL_X1 FILLER_2_541 ();
 FILLCELL_X1 FILLER_2_551 ();
 FILLCELL_X2 FILLER_2_559 ();
 FILLCELL_X1 FILLER_2_561 ();
 FILLCELL_X2 FILLER_2_576 ();
 FILLCELL_X4 FILLER_2_599 ();
 FILLCELL_X1 FILLER_2_603 ();
 FILLCELL_X2 FILLER_2_610 ();
 FILLCELL_X1 FILLER_2_612 ();
 FILLCELL_X4 FILLER_2_632 ();
 FILLCELL_X4 FILLER_2_643 ();
 FILLCELL_X2 FILLER_2_647 ();
 FILLCELL_X1 FILLER_2_649 ();
 FILLCELL_X32 FILLER_2_671 ();
 FILLCELL_X32 FILLER_2_703 ();
 FILLCELL_X8 FILLER_2_735 ();
 FILLCELL_X4 FILLER_2_743 ();
 FILLCELL_X8 FILLER_2_758 ();
 FILLCELL_X2 FILLER_2_766 ();
 FILLCELL_X1 FILLER_2_768 ();
 FILLCELL_X1 FILLER_2_784 ();
 FILLCELL_X1 FILLER_2_791 ();
 FILLCELL_X2 FILLER_2_795 ();
 FILLCELL_X2 FILLER_2_810 ();
 FILLCELL_X1 FILLER_2_812 ();
 FILLCELL_X1 FILLER_2_822 ();
 FILLCELL_X2 FILLER_2_827 ();
 FILLCELL_X1 FILLER_2_829 ();
 FILLCELL_X8 FILLER_2_833 ();
 FILLCELL_X2 FILLER_2_841 ();
 FILLCELL_X1 FILLER_2_846 ();
 FILLCELL_X8 FILLER_2_855 ();
 FILLCELL_X2 FILLER_2_863 ();
 FILLCELL_X1 FILLER_2_870 ();
 FILLCELL_X2 FILLER_2_889 ();
 FILLCELL_X1 FILLER_2_891 ();
 FILLCELL_X4 FILLER_2_896 ();
 FILLCELL_X4 FILLER_2_907 ();
 FILLCELL_X1 FILLER_2_915 ();
 FILLCELL_X4 FILLER_2_923 ();
 FILLCELL_X8 FILLER_2_934 ();
 FILLCELL_X32 FILLER_2_953 ();
 FILLCELL_X32 FILLER_2_985 ();
 FILLCELL_X32 FILLER_2_1017 ();
 FILLCELL_X16 FILLER_2_1049 ();
 FILLCELL_X4 FILLER_2_1065 ();
 FILLCELL_X2 FILLER_2_1094 ();
 FILLCELL_X2 FILLER_2_1115 ();
 FILLCELL_X1 FILLER_2_1117 ();
 FILLCELL_X4 FILLER_2_1130 ();
 FILLCELL_X2 FILLER_2_1134 ();
 FILLCELL_X4 FILLER_2_1145 ();
 FILLCELL_X1 FILLER_2_1149 ();
 FILLCELL_X8 FILLER_2_1191 ();
 FILLCELL_X2 FILLER_2_1199 ();
 FILLCELL_X32 FILLER_2_1228 ();
 FILLCELL_X32 FILLER_2_1260 ();
 FILLCELL_X32 FILLER_2_1292 ();
 FILLCELL_X32 FILLER_2_1324 ();
 FILLCELL_X32 FILLER_2_1356 ();
 FILLCELL_X32 FILLER_2_1388 ();
 FILLCELL_X32 FILLER_2_1420 ();
 FILLCELL_X32 FILLER_2_1452 ();
 FILLCELL_X32 FILLER_2_1484 ();
 FILLCELL_X32 FILLER_2_1516 ();
 FILLCELL_X32 FILLER_2_1548 ();
 FILLCELL_X32 FILLER_2_1580 ();
 FILLCELL_X32 FILLER_2_1612 ();
 FILLCELL_X4 FILLER_2_1644 ();
 FILLCELL_X2 FILLER_2_1648 ();
 FILLCELL_X1 FILLER_2_1650 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X16 FILLER_3_193 ();
 FILLCELL_X8 FILLER_3_209 ();
 FILLCELL_X4 FILLER_3_217 ();
 FILLCELL_X1 FILLER_3_221 ();
 FILLCELL_X4 FILLER_3_226 ();
 FILLCELL_X2 FILLER_3_237 ();
 FILLCELL_X1 FILLER_3_239 ();
 FILLCELL_X2 FILLER_3_247 ();
 FILLCELL_X4 FILLER_3_267 ();
 FILLCELL_X2 FILLER_3_288 ();
 FILLCELL_X4 FILLER_3_297 ();
 FILLCELL_X4 FILLER_3_321 ();
 FILLCELL_X1 FILLER_3_325 ();
 FILLCELL_X1 FILLER_3_335 ();
 FILLCELL_X8 FILLER_3_379 ();
 FILLCELL_X4 FILLER_3_387 ();
 FILLCELL_X1 FILLER_3_391 ();
 FILLCELL_X1 FILLER_3_399 ();
 FILLCELL_X32 FILLER_3_413 ();
 FILLCELL_X8 FILLER_3_445 ();
 FILLCELL_X4 FILLER_3_460 ();
 FILLCELL_X2 FILLER_3_484 ();
 FILLCELL_X8 FILLER_3_495 ();
 FILLCELL_X2 FILLER_3_503 ();
 FILLCELL_X2 FILLER_3_518 ();
 FILLCELL_X4 FILLER_3_524 ();
 FILLCELL_X1 FILLER_3_528 ();
 FILLCELL_X4 FILLER_3_550 ();
 FILLCELL_X1 FILLER_3_554 ();
 FILLCELL_X4 FILLER_3_558 ();
 FILLCELL_X2 FILLER_3_562 ();
 FILLCELL_X4 FILLER_3_573 ();
 FILLCELL_X4 FILLER_3_602 ();
 FILLCELL_X2 FILLER_3_606 ();
 FILLCELL_X2 FILLER_3_616 ();
 FILLCELL_X1 FILLER_3_618 ();
 FILLCELL_X4 FILLER_3_632 ();
 FILLCELL_X2 FILLER_3_636 ();
 FILLCELL_X1 FILLER_3_645 ();
 FILLCELL_X1 FILLER_3_662 ();
 FILLCELL_X4 FILLER_3_670 ();
 FILLCELL_X2 FILLER_3_674 ();
 FILLCELL_X1 FILLER_3_676 ();
 FILLCELL_X32 FILLER_3_684 ();
 FILLCELL_X32 FILLER_3_716 ();
 FILLCELL_X16 FILLER_3_748 ();
 FILLCELL_X2 FILLER_3_778 ();
 FILLCELL_X4 FILLER_3_788 ();
 FILLCELL_X1 FILLER_3_792 ();
 FILLCELL_X8 FILLER_3_797 ();
 FILLCELL_X4 FILLER_3_805 ();
 FILLCELL_X2 FILLER_3_809 ();
 FILLCELL_X1 FILLER_3_811 ();
 FILLCELL_X8 FILLER_3_819 ();
 FILLCELL_X1 FILLER_3_834 ();
 FILLCELL_X4 FILLER_3_847 ();
 FILLCELL_X4 FILLER_3_856 ();
 FILLCELL_X2 FILLER_3_864 ();
 FILLCELL_X1 FILLER_3_866 ();
 FILLCELL_X8 FILLER_3_884 ();
 FILLCELL_X1 FILLER_3_892 ();
 FILLCELL_X4 FILLER_3_902 ();
 FILLCELL_X1 FILLER_3_906 ();
 FILLCELL_X1 FILLER_3_914 ();
 FILLCELL_X2 FILLER_3_922 ();
 FILLCELL_X1 FILLER_3_924 ();
 FILLCELL_X2 FILLER_3_937 ();
 FILLCELL_X1 FILLER_3_939 ();
 FILLCELL_X32 FILLER_3_947 ();
 FILLCELL_X32 FILLER_3_979 ();
 FILLCELL_X32 FILLER_3_1011 ();
 FILLCELL_X8 FILLER_3_1043 ();
 FILLCELL_X4 FILLER_3_1051 ();
 FILLCELL_X2 FILLER_3_1055 ();
 FILLCELL_X1 FILLER_3_1057 ();
 FILLCELL_X2 FILLER_3_1100 ();
 FILLCELL_X1 FILLER_3_1102 ();
 FILLCELL_X4 FILLER_3_1113 ();
 FILLCELL_X1 FILLER_3_1117 ();
 FILLCELL_X1 FILLER_3_1127 ();
 FILLCELL_X2 FILLER_3_1132 ();
 FILLCELL_X1 FILLER_3_1134 ();
 FILLCELL_X4 FILLER_3_1139 ();
 FILLCELL_X1 FILLER_3_1143 ();
 FILLCELL_X8 FILLER_3_1172 ();
 FILLCELL_X2 FILLER_3_1180 ();
 FILLCELL_X1 FILLER_3_1182 ();
 FILLCELL_X4 FILLER_3_1213 ();
 FILLCELL_X2 FILLER_3_1217 ();
 FILLCELL_X1 FILLER_3_1219 ();
 FILLCELL_X32 FILLER_3_1227 ();
 FILLCELL_X4 FILLER_3_1259 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1296 ();
 FILLCELL_X32 FILLER_3_1328 ();
 FILLCELL_X32 FILLER_3_1360 ();
 FILLCELL_X32 FILLER_3_1392 ();
 FILLCELL_X32 FILLER_3_1424 ();
 FILLCELL_X32 FILLER_3_1456 ();
 FILLCELL_X32 FILLER_3_1488 ();
 FILLCELL_X32 FILLER_3_1520 ();
 FILLCELL_X32 FILLER_3_1552 ();
 FILLCELL_X32 FILLER_3_1584 ();
 FILLCELL_X32 FILLER_3_1616 ();
 FILLCELL_X2 FILLER_3_1648 ();
 FILLCELL_X1 FILLER_3_1650 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X16 FILLER_4_193 ();
 FILLCELL_X1 FILLER_4_209 ();
 FILLCELL_X1 FILLER_4_227 ();
 FILLCELL_X4 FILLER_4_247 ();
 FILLCELL_X8 FILLER_4_266 ();
 FILLCELL_X4 FILLER_4_274 ();
 FILLCELL_X8 FILLER_4_285 ();
 FILLCELL_X4 FILLER_4_293 ();
 FILLCELL_X4 FILLER_4_311 ();
 FILLCELL_X2 FILLER_4_315 ();
 FILLCELL_X1 FILLER_4_317 ();
 FILLCELL_X4 FILLER_4_327 ();
 FILLCELL_X2 FILLER_4_331 ();
 FILLCELL_X2 FILLER_4_340 ();
 FILLCELL_X1 FILLER_4_342 ();
 FILLCELL_X8 FILLER_4_361 ();
 FILLCELL_X1 FILLER_4_369 ();
 FILLCELL_X32 FILLER_4_388 ();
 FILLCELL_X32 FILLER_4_420 ();
 FILLCELL_X8 FILLER_4_452 ();
 FILLCELL_X2 FILLER_4_460 ();
 FILLCELL_X4 FILLER_4_497 ();
 FILLCELL_X2 FILLER_4_501 ();
 FILLCELL_X1 FILLER_4_503 ();
 FILLCELL_X4 FILLER_4_518 ();
 FILLCELL_X1 FILLER_4_522 ();
 FILLCELL_X2 FILLER_4_546 ();
 FILLCELL_X1 FILLER_4_557 ();
 FILLCELL_X1 FILLER_4_576 ();
 FILLCELL_X16 FILLER_4_586 ();
 FILLCELL_X2 FILLER_4_602 ();
 FILLCELL_X2 FILLER_4_607 ();
 FILLCELL_X1 FILLER_4_609 ();
 FILLCELL_X1 FILLER_4_623 ();
 FILLCELL_X8 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_666 ();
 FILLCELL_X32 FILLER_4_698 ();
 FILLCELL_X8 FILLER_4_730 ();
 FILLCELL_X1 FILLER_4_738 ();
 FILLCELL_X4 FILLER_4_793 ();
 FILLCELL_X2 FILLER_4_797 ();
 FILLCELL_X8 FILLER_4_804 ();
 FILLCELL_X4 FILLER_4_812 ();
 FILLCELL_X2 FILLER_4_816 ();
 FILLCELL_X1 FILLER_4_818 ();
 FILLCELL_X2 FILLER_4_831 ();
 FILLCELL_X1 FILLER_4_833 ();
 FILLCELL_X2 FILLER_4_842 ();
 FILLCELL_X1 FILLER_4_848 ();
 FILLCELL_X8 FILLER_4_864 ();
 FILLCELL_X2 FILLER_4_872 ();
 FILLCELL_X1 FILLER_4_874 ();
 FILLCELL_X2 FILLER_4_894 ();
 FILLCELL_X1 FILLER_4_896 ();
 FILLCELL_X16 FILLER_4_921 ();
 FILLCELL_X1 FILLER_4_937 ();
 FILLCELL_X32 FILLER_4_967 ();
 FILLCELL_X32 FILLER_4_999 ();
 FILLCELL_X8 FILLER_4_1031 ();
 FILLCELL_X1 FILLER_4_1039 ();
 FILLCELL_X8 FILLER_4_1047 ();
 FILLCELL_X2 FILLER_4_1055 ();
 FILLCELL_X4 FILLER_4_1068 ();
 FILLCELL_X2 FILLER_4_1072 ();
 FILLCELL_X1 FILLER_4_1092 ();
 FILLCELL_X2 FILLER_4_1097 ();
 FILLCELL_X2 FILLER_4_1106 ();
 FILLCELL_X1 FILLER_4_1122 ();
 FILLCELL_X8 FILLER_4_1131 ();
 FILLCELL_X4 FILLER_4_1139 ();
 FILLCELL_X2 FILLER_4_1143 ();
 FILLCELL_X4 FILLER_4_1194 ();
 FILLCELL_X4 FILLER_4_1219 ();
 FILLCELL_X1 FILLER_4_1223 ();
 FILLCELL_X4 FILLER_4_1231 ();
 FILLCELL_X2 FILLER_4_1235 ();
 FILLCELL_X32 FILLER_4_1250 ();
 FILLCELL_X32 FILLER_4_1282 ();
 FILLCELL_X32 FILLER_4_1314 ();
 FILLCELL_X32 FILLER_4_1346 ();
 FILLCELL_X32 FILLER_4_1378 ();
 FILLCELL_X32 FILLER_4_1410 ();
 FILLCELL_X32 FILLER_4_1442 ();
 FILLCELL_X32 FILLER_4_1474 ();
 FILLCELL_X32 FILLER_4_1506 ();
 FILLCELL_X32 FILLER_4_1538 ();
 FILLCELL_X32 FILLER_4_1570 ();
 FILLCELL_X32 FILLER_4_1602 ();
 FILLCELL_X16 FILLER_4_1634 ();
 FILLCELL_X1 FILLER_4_1650 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X16 FILLER_5_161 ();
 FILLCELL_X8 FILLER_5_177 ();
 FILLCELL_X4 FILLER_5_196 ();
 FILLCELL_X2 FILLER_5_200 ();
 FILLCELL_X8 FILLER_5_215 ();
 FILLCELL_X1 FILLER_5_223 ();
 FILLCELL_X8 FILLER_5_249 ();
 FILLCELL_X2 FILLER_5_257 ();
 FILLCELL_X1 FILLER_5_259 ();
 FILLCELL_X2 FILLER_5_265 ();
 FILLCELL_X1 FILLER_5_290 ();
 FILLCELL_X4 FILLER_5_316 ();
 FILLCELL_X4 FILLER_5_331 ();
 FILLCELL_X1 FILLER_5_335 ();
 FILLCELL_X32 FILLER_5_391 ();
 FILLCELL_X32 FILLER_5_423 ();
 FILLCELL_X1 FILLER_5_455 ();
 FILLCELL_X4 FILLER_5_514 ();
 FILLCELL_X1 FILLER_5_518 ();
 FILLCELL_X2 FILLER_5_530 ();
 FILLCELL_X1 FILLER_5_532 ();
 FILLCELL_X16 FILLER_5_577 ();
 FILLCELL_X8 FILLER_5_593 ();
 FILLCELL_X2 FILLER_5_601 ();
 FILLCELL_X1 FILLER_5_603 ();
 FILLCELL_X8 FILLER_5_626 ();
 FILLCELL_X2 FILLER_5_648 ();
 FILLCELL_X2 FILLER_5_657 ();
 FILLCELL_X32 FILLER_5_663 ();
 FILLCELL_X32 FILLER_5_695 ();
 FILLCELL_X16 FILLER_5_727 ();
 FILLCELL_X8 FILLER_5_752 ();
 FILLCELL_X4 FILLER_5_760 ();
 FILLCELL_X4 FILLER_5_769 ();
 FILLCELL_X2 FILLER_5_788 ();
 FILLCELL_X1 FILLER_5_790 ();
 FILLCELL_X2 FILLER_5_797 ();
 FILLCELL_X1 FILLER_5_799 ();
 FILLCELL_X4 FILLER_5_808 ();
 FILLCELL_X2 FILLER_5_819 ();
 FILLCELL_X1 FILLER_5_830 ();
 FILLCELL_X16 FILLER_5_836 ();
 FILLCELL_X2 FILLER_5_861 ();
 FILLCELL_X2 FILLER_5_877 ();
 FILLCELL_X2 FILLER_5_888 ();
 FILLCELL_X1 FILLER_5_890 ();
 FILLCELL_X8 FILLER_5_895 ();
 FILLCELL_X2 FILLER_5_903 ();
 FILLCELL_X4 FILLER_5_944 ();
 FILLCELL_X32 FILLER_5_952 ();
 FILLCELL_X32 FILLER_5_984 ();
 FILLCELL_X8 FILLER_5_1016 ();
 FILLCELL_X4 FILLER_5_1024 ();
 FILLCELL_X1 FILLER_5_1028 ();
 FILLCELL_X1 FILLER_5_1040 ();
 FILLCELL_X2 FILLER_5_1053 ();
 FILLCELL_X2 FILLER_5_1076 ();
 FILLCELL_X2 FILLER_5_1097 ();
 FILLCELL_X2 FILLER_5_1103 ();
 FILLCELL_X2 FILLER_5_1112 ();
 FILLCELL_X1 FILLER_5_1114 ();
 FILLCELL_X2 FILLER_5_1119 ();
 FILLCELL_X1 FILLER_5_1121 ();
 FILLCELL_X8 FILLER_5_1127 ();
 FILLCELL_X4 FILLER_5_1135 ();
 FILLCELL_X1 FILLER_5_1139 ();
 FILLCELL_X2 FILLER_5_1143 ();
 FILLCELL_X1 FILLER_5_1145 ();
 FILLCELL_X4 FILLER_5_1153 ();
 FILLCELL_X2 FILLER_5_1157 ();
 FILLCELL_X2 FILLER_5_1177 ();
 FILLCELL_X1 FILLER_5_1179 ();
 FILLCELL_X4 FILLER_5_1190 ();
 FILLCELL_X1 FILLER_5_1194 ();
 FILLCELL_X4 FILLER_5_1215 ();
 FILLCELL_X1 FILLER_5_1219 ();
 FILLCELL_X4 FILLER_5_1232 ();
 FILLCELL_X2 FILLER_5_1236 ();
 FILLCELL_X8 FILLER_5_1248 ();
 FILLCELL_X4 FILLER_5_1256 ();
 FILLCELL_X2 FILLER_5_1260 ();
 FILLCELL_X1 FILLER_5_1262 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X32 FILLER_5_1296 ();
 FILLCELL_X32 FILLER_5_1328 ();
 FILLCELL_X32 FILLER_5_1360 ();
 FILLCELL_X32 FILLER_5_1392 ();
 FILLCELL_X32 FILLER_5_1424 ();
 FILLCELL_X32 FILLER_5_1456 ();
 FILLCELL_X32 FILLER_5_1488 ();
 FILLCELL_X32 FILLER_5_1520 ();
 FILLCELL_X32 FILLER_5_1552 ();
 FILLCELL_X32 FILLER_5_1584 ();
 FILLCELL_X32 FILLER_5_1616 ();
 FILLCELL_X2 FILLER_5_1648 ();
 FILLCELL_X1 FILLER_5_1650 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X16 FILLER_6_161 ();
 FILLCELL_X4 FILLER_6_177 ();
 FILLCELL_X1 FILLER_6_181 ();
 FILLCELL_X4 FILLER_6_199 ();
 FILLCELL_X2 FILLER_6_203 ();
 FILLCELL_X2 FILLER_6_227 ();
 FILLCELL_X1 FILLER_6_229 ();
 FILLCELL_X1 FILLER_6_234 ();
 FILLCELL_X8 FILLER_6_249 ();
 FILLCELL_X4 FILLER_6_257 ();
 FILLCELL_X2 FILLER_6_261 ();
 FILLCELL_X2 FILLER_6_275 ();
 FILLCELL_X4 FILLER_6_280 ();
 FILLCELL_X2 FILLER_6_284 ();
 FILLCELL_X1 FILLER_6_286 ();
 FILLCELL_X4 FILLER_6_296 ();
 FILLCELL_X4 FILLER_6_321 ();
 FILLCELL_X2 FILLER_6_325 ();
 FILLCELL_X4 FILLER_6_336 ();
 FILLCELL_X2 FILLER_6_354 ();
 FILLCELL_X1 FILLER_6_356 ();
 FILLCELL_X1 FILLER_6_361 ();
 FILLCELL_X1 FILLER_6_369 ();
 FILLCELL_X1 FILLER_6_379 ();
 FILLCELL_X4 FILLER_6_399 ();
 FILLCELL_X1 FILLER_6_403 ();
 FILLCELL_X32 FILLER_6_411 ();
 FILLCELL_X8 FILLER_6_443 ();
 FILLCELL_X2 FILLER_6_451 ();
 FILLCELL_X1 FILLER_6_453 ();
 FILLCELL_X1 FILLER_6_471 ();
 FILLCELL_X4 FILLER_6_496 ();
 FILLCELL_X16 FILLER_6_507 ();
 FILLCELL_X4 FILLER_6_523 ();
 FILLCELL_X2 FILLER_6_527 ();
 FILLCELL_X8 FILLER_6_545 ();
 FILLCELL_X4 FILLER_6_557 ();
 FILLCELL_X2 FILLER_6_561 ();
 FILLCELL_X1 FILLER_6_563 ();
 FILLCELL_X8 FILLER_6_571 ();
 FILLCELL_X2 FILLER_6_579 ();
 FILLCELL_X8 FILLER_6_595 ();
 FILLCELL_X4 FILLER_6_603 ();
 FILLCELL_X2 FILLER_6_607 ();
 FILLCELL_X2 FILLER_6_614 ();
 FILLCELL_X1 FILLER_6_616 ();
 FILLCELL_X2 FILLER_6_621 ();
 FILLCELL_X1 FILLER_6_623 ();
 FILLCELL_X2 FILLER_6_632 ();
 FILLCELL_X1 FILLER_6_655 ();
 FILLCELL_X2 FILLER_6_663 ();
 FILLCELL_X4 FILLER_6_676 ();
 FILLCELL_X1 FILLER_6_680 ();
 FILLCELL_X32 FILLER_6_688 ();
 FILLCELL_X16 FILLER_6_720 ();
 FILLCELL_X4 FILLER_6_736 ();
 FILLCELL_X2 FILLER_6_740 ();
 FILLCELL_X1 FILLER_6_742 ();
 FILLCELL_X4 FILLER_6_746 ();
 FILLCELL_X1 FILLER_6_750 ();
 FILLCELL_X8 FILLER_6_765 ();
 FILLCELL_X2 FILLER_6_787 ();
 FILLCELL_X2 FILLER_6_792 ();
 FILLCELL_X2 FILLER_6_821 ();
 FILLCELL_X2 FILLER_6_826 ();
 FILLCELL_X1 FILLER_6_828 ();
 FILLCELL_X4 FILLER_6_834 ();
 FILLCELL_X1 FILLER_6_838 ();
 FILLCELL_X2 FILLER_6_848 ();
 FILLCELL_X4 FILLER_6_880 ();
 FILLCELL_X1 FILLER_6_884 ();
 FILLCELL_X1 FILLER_6_895 ();
 FILLCELL_X1 FILLER_6_901 ();
 FILLCELL_X2 FILLER_6_917 ();
 FILLCELL_X1 FILLER_6_919 ();
 FILLCELL_X2 FILLER_6_939 ();
 FILLCELL_X4 FILLER_6_955 ();
 FILLCELL_X2 FILLER_6_959 ();
 FILLCELL_X1 FILLER_6_961 ();
 FILLCELL_X1 FILLER_6_967 ();
 FILLCELL_X32 FILLER_6_974 ();
 FILLCELL_X16 FILLER_6_1006 ();
 FILLCELL_X4 FILLER_6_1022 ();
 FILLCELL_X1 FILLER_6_1026 ();
 FILLCELL_X2 FILLER_6_1036 ();
 FILLCELL_X1 FILLER_6_1038 ();
 FILLCELL_X1 FILLER_6_1043 ();
 FILLCELL_X1 FILLER_6_1049 ();
 FILLCELL_X1 FILLER_6_1059 ();
 FILLCELL_X2 FILLER_6_1076 ();
 FILLCELL_X1 FILLER_6_1078 ();
 FILLCELL_X4 FILLER_6_1163 ();
 FILLCELL_X2 FILLER_6_1167 ();
 FILLCELL_X1 FILLER_6_1173 ();
 FILLCELL_X2 FILLER_6_1177 ();
 FILLCELL_X2 FILLER_6_1190 ();
 FILLCELL_X1 FILLER_6_1201 ();
 FILLCELL_X1 FILLER_6_1210 ();
 FILLCELL_X2 FILLER_6_1227 ();
 FILLCELL_X1 FILLER_6_1238 ();
 FILLCELL_X16 FILLER_6_1246 ();
 FILLCELL_X32 FILLER_6_1280 ();
 FILLCELL_X32 FILLER_6_1312 ();
 FILLCELL_X32 FILLER_6_1344 ();
 FILLCELL_X32 FILLER_6_1376 ();
 FILLCELL_X32 FILLER_6_1408 ();
 FILLCELL_X32 FILLER_6_1440 ();
 FILLCELL_X32 FILLER_6_1472 ();
 FILLCELL_X32 FILLER_6_1504 ();
 FILLCELL_X32 FILLER_6_1536 ();
 FILLCELL_X32 FILLER_6_1568 ();
 FILLCELL_X32 FILLER_6_1600 ();
 FILLCELL_X16 FILLER_6_1632 ();
 FILLCELL_X2 FILLER_6_1648 ();
 FILLCELL_X1 FILLER_6_1650 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X1 FILLER_7_193 ();
 FILLCELL_X2 FILLER_7_201 ();
 FILLCELL_X8 FILLER_7_208 ();
 FILLCELL_X4 FILLER_7_216 ();
 FILLCELL_X2 FILLER_7_229 ();
 FILLCELL_X1 FILLER_7_231 ();
 FILLCELL_X2 FILLER_7_241 ();
 FILLCELL_X1 FILLER_7_243 ();
 FILLCELL_X4 FILLER_7_258 ();
 FILLCELL_X1 FILLER_7_262 ();
 FILLCELL_X4 FILLER_7_268 ();
 FILLCELL_X1 FILLER_7_288 ();
 FILLCELL_X2 FILLER_7_320 ();
 FILLCELL_X4 FILLER_7_329 ();
 FILLCELL_X8 FILLER_7_374 ();
 FILLCELL_X1 FILLER_7_382 ();
 FILLCELL_X2 FILLER_7_390 ();
 FILLCELL_X1 FILLER_7_392 ();
 FILLCELL_X16 FILLER_7_411 ();
 FILLCELL_X8 FILLER_7_427 ();
 FILLCELL_X1 FILLER_7_435 ();
 FILLCELL_X4 FILLER_7_453 ();
 FILLCELL_X1 FILLER_7_457 ();
 FILLCELL_X1 FILLER_7_465 ();
 FILLCELL_X2 FILLER_7_473 ();
 FILLCELL_X2 FILLER_7_486 ();
 FILLCELL_X2 FILLER_7_498 ();
 FILLCELL_X1 FILLER_7_500 ();
 FILLCELL_X1 FILLER_7_505 ();
 FILLCELL_X2 FILLER_7_511 ();
 FILLCELL_X1 FILLER_7_513 ();
 FILLCELL_X4 FILLER_7_527 ();
 FILLCELL_X2 FILLER_7_531 ();
 FILLCELL_X2 FILLER_7_559 ();
 FILLCELL_X1 FILLER_7_561 ();
 FILLCELL_X4 FILLER_7_570 ();
 FILLCELL_X16 FILLER_7_592 ();
 FILLCELL_X8 FILLER_7_608 ();
 FILLCELL_X4 FILLER_7_616 ();
 FILLCELL_X8 FILLER_7_624 ();
 FILLCELL_X2 FILLER_7_632 ();
 FILLCELL_X8 FILLER_7_645 ();
 FILLCELL_X2 FILLER_7_653 ();
 FILLCELL_X4 FILLER_7_659 ();
 FILLCELL_X2 FILLER_7_663 ();
 FILLCELL_X32 FILLER_7_669 ();
 FILLCELL_X32 FILLER_7_701 ();
 FILLCELL_X16 FILLER_7_733 ();
 FILLCELL_X4 FILLER_7_749 ();
 FILLCELL_X1 FILLER_7_753 ();
 FILLCELL_X1 FILLER_7_794 ();
 FILLCELL_X2 FILLER_7_800 ();
 FILLCELL_X4 FILLER_7_815 ();
 FILLCELL_X2 FILLER_7_819 ();
 FILLCELL_X1 FILLER_7_838 ();
 FILLCELL_X4 FILLER_7_864 ();
 FILLCELL_X1 FILLER_7_868 ();
 FILLCELL_X2 FILLER_7_873 ();
 FILLCELL_X2 FILLER_7_879 ();
 FILLCELL_X1 FILLER_7_881 ();
 FILLCELL_X8 FILLER_7_886 ();
 FILLCELL_X2 FILLER_7_894 ();
 FILLCELL_X8 FILLER_7_903 ();
 FILLCELL_X4 FILLER_7_911 ();
 FILLCELL_X4 FILLER_7_925 ();
 FILLCELL_X2 FILLER_7_929 ();
 FILLCELL_X1 FILLER_7_952 ();
 FILLCELL_X32 FILLER_7_957 ();
 FILLCELL_X32 FILLER_7_989 ();
 FILLCELL_X4 FILLER_7_1021 ();
 FILLCELL_X2 FILLER_7_1025 ();
 FILLCELL_X2 FILLER_7_1044 ();
 FILLCELL_X1 FILLER_7_1063 ();
 FILLCELL_X1 FILLER_7_1081 ();
 FILLCELL_X1 FILLER_7_1092 ();
 FILLCELL_X2 FILLER_7_1097 ();
 FILLCELL_X2 FILLER_7_1113 ();
 FILLCELL_X1 FILLER_7_1115 ();
 FILLCELL_X4 FILLER_7_1123 ();
 FILLCELL_X4 FILLER_7_1134 ();
 FILLCELL_X1 FILLER_7_1138 ();
 FILLCELL_X2 FILLER_7_1143 ();
 FILLCELL_X1 FILLER_7_1149 ();
 FILLCELL_X1 FILLER_7_1167 ();
 FILLCELL_X1 FILLER_7_1172 ();
 FILLCELL_X2 FILLER_7_1178 ();
 FILLCELL_X8 FILLER_7_1188 ();
 FILLCELL_X4 FILLER_7_1196 ();
 FILLCELL_X2 FILLER_7_1200 ();
 FILLCELL_X4 FILLER_7_1209 ();
 FILLCELL_X2 FILLER_7_1213 ();
 FILLCELL_X1 FILLER_7_1215 ();
 FILLCELL_X4 FILLER_7_1259 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X32 FILLER_7_1296 ();
 FILLCELL_X32 FILLER_7_1328 ();
 FILLCELL_X32 FILLER_7_1360 ();
 FILLCELL_X32 FILLER_7_1392 ();
 FILLCELL_X32 FILLER_7_1424 ();
 FILLCELL_X32 FILLER_7_1456 ();
 FILLCELL_X32 FILLER_7_1488 ();
 FILLCELL_X32 FILLER_7_1520 ();
 FILLCELL_X32 FILLER_7_1552 ();
 FILLCELL_X32 FILLER_7_1584 ();
 FILLCELL_X32 FILLER_7_1616 ();
 FILLCELL_X2 FILLER_7_1648 ();
 FILLCELL_X1 FILLER_7_1650 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X16 FILLER_8_161 ();
 FILLCELL_X8 FILLER_8_177 ();
 FILLCELL_X4 FILLER_8_185 ();
 FILLCELL_X2 FILLER_8_189 ();
 FILLCELL_X8 FILLER_8_200 ();
 FILLCELL_X1 FILLER_8_208 ();
 FILLCELL_X2 FILLER_8_219 ();
 FILLCELL_X16 FILLER_8_225 ();
 FILLCELL_X1 FILLER_8_241 ();
 FILLCELL_X8 FILLER_8_258 ();
 FILLCELL_X4 FILLER_8_266 ();
 FILLCELL_X1 FILLER_8_270 ();
 FILLCELL_X2 FILLER_8_284 ();
 FILLCELL_X1 FILLER_8_286 ();
 FILLCELL_X2 FILLER_8_297 ();
 FILLCELL_X8 FILLER_8_366 ();
 FILLCELL_X2 FILLER_8_374 ();
 FILLCELL_X1 FILLER_8_376 ();
 FILLCELL_X16 FILLER_8_420 ();
 FILLCELL_X1 FILLER_8_436 ();
 FILLCELL_X1 FILLER_8_454 ();
 FILLCELL_X1 FILLER_8_462 ();
 FILLCELL_X4 FILLER_8_467 ();
 FILLCELL_X1 FILLER_8_471 ();
 FILLCELL_X2 FILLER_8_480 ();
 FILLCELL_X1 FILLER_8_485 ();
 FILLCELL_X1 FILLER_8_491 ();
 FILLCELL_X1 FILLER_8_496 ();
 FILLCELL_X2 FILLER_8_511 ();
 FILLCELL_X8 FILLER_8_533 ();
 FILLCELL_X2 FILLER_8_541 ();
 FILLCELL_X1 FILLER_8_543 ();
 FILLCELL_X4 FILLER_8_548 ();
 FILLCELL_X1 FILLER_8_567 ();
 FILLCELL_X4 FILLER_8_572 ();
 FILLCELL_X4 FILLER_8_594 ();
 FILLCELL_X1 FILLER_8_598 ();
 FILLCELL_X2 FILLER_8_603 ();
 FILLCELL_X2 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_632 ();
 FILLCELL_X1 FILLER_8_641 ();
 FILLCELL_X4 FILLER_8_659 ();
 FILLCELL_X2 FILLER_8_663 ();
 FILLCELL_X1 FILLER_8_665 ();
 FILLCELL_X2 FILLER_8_674 ();
 FILLCELL_X32 FILLER_8_680 ();
 FILLCELL_X16 FILLER_8_712 ();
 FILLCELL_X8 FILLER_8_728 ();
 FILLCELL_X2 FILLER_8_736 ();
 FILLCELL_X1 FILLER_8_738 ();
 FILLCELL_X8 FILLER_8_749 ();
 FILLCELL_X1 FILLER_8_757 ();
 FILLCELL_X1 FILLER_8_767 ();
 FILLCELL_X2 FILLER_8_772 ();
 FILLCELL_X1 FILLER_8_777 ();
 FILLCELL_X1 FILLER_8_789 ();
 FILLCELL_X1 FILLER_8_797 ();
 FILLCELL_X1 FILLER_8_802 ();
 FILLCELL_X2 FILLER_8_814 ();
 FILLCELL_X1 FILLER_8_816 ();
 FILLCELL_X4 FILLER_8_821 ();
 FILLCELL_X1 FILLER_8_825 ();
 FILLCELL_X8 FILLER_8_833 ();
 FILLCELL_X4 FILLER_8_841 ();
 FILLCELL_X8 FILLER_8_850 ();
 FILLCELL_X2 FILLER_8_858 ();
 FILLCELL_X4 FILLER_8_896 ();
 FILLCELL_X1 FILLER_8_900 ();
 FILLCELL_X2 FILLER_8_936 ();
 FILLCELL_X2 FILLER_8_955 ();
 FILLCELL_X32 FILLER_8_976 ();
 FILLCELL_X8 FILLER_8_1008 ();
 FILLCELL_X4 FILLER_8_1051 ();
 FILLCELL_X4 FILLER_8_1062 ();
 FILLCELL_X1 FILLER_8_1066 ();
 FILLCELL_X1 FILLER_8_1085 ();
 FILLCELL_X16 FILLER_8_1102 ();
 FILLCELL_X4 FILLER_8_1118 ();
 FILLCELL_X2 FILLER_8_1122 ();
 FILLCELL_X1 FILLER_8_1124 ();
 FILLCELL_X4 FILLER_8_1137 ();
 FILLCELL_X1 FILLER_8_1141 ();
 FILLCELL_X16 FILLER_8_1149 ();
 FILLCELL_X4 FILLER_8_1165 ();
 FILLCELL_X1 FILLER_8_1192 ();
 FILLCELL_X8 FILLER_8_1219 ();
 FILLCELL_X4 FILLER_8_1227 ();
 FILLCELL_X2 FILLER_8_1231 ();
 FILLCELL_X32 FILLER_8_1245 ();
 FILLCELL_X32 FILLER_8_1277 ();
 FILLCELL_X32 FILLER_8_1309 ();
 FILLCELL_X32 FILLER_8_1341 ();
 FILLCELL_X32 FILLER_8_1373 ();
 FILLCELL_X32 FILLER_8_1405 ();
 FILLCELL_X32 FILLER_8_1437 ();
 FILLCELL_X32 FILLER_8_1469 ();
 FILLCELL_X32 FILLER_8_1501 ();
 FILLCELL_X32 FILLER_8_1533 ();
 FILLCELL_X32 FILLER_8_1565 ();
 FILLCELL_X32 FILLER_8_1597 ();
 FILLCELL_X16 FILLER_8_1629 ();
 FILLCELL_X4 FILLER_8_1645 ();
 FILLCELL_X2 FILLER_8_1649 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X16 FILLER_9_161 ();
 FILLCELL_X8 FILLER_9_177 ();
 FILLCELL_X4 FILLER_9_194 ();
 FILLCELL_X2 FILLER_9_198 ();
 FILLCELL_X1 FILLER_9_200 ();
 FILLCELL_X4 FILLER_9_228 ();
 FILLCELL_X1 FILLER_9_263 ();
 FILLCELL_X4 FILLER_9_267 ();
 FILLCELL_X1 FILLER_9_271 ();
 FILLCELL_X2 FILLER_9_281 ();
 FILLCELL_X1 FILLER_9_283 ();
 FILLCELL_X8 FILLER_9_301 ();
 FILLCELL_X4 FILLER_9_309 ();
 FILLCELL_X4 FILLER_9_320 ();
 FILLCELL_X2 FILLER_9_324 ();
 FILLCELL_X4 FILLER_9_331 ();
 FILLCELL_X1 FILLER_9_335 ();
 FILLCELL_X4 FILLER_9_345 ();
 FILLCELL_X32 FILLER_9_411 ();
 FILLCELL_X8 FILLER_9_443 ();
 FILLCELL_X4 FILLER_9_451 ();
 FILLCELL_X2 FILLER_9_455 ();
 FILLCELL_X1 FILLER_9_457 ();
 FILLCELL_X1 FILLER_9_465 ();
 FILLCELL_X1 FILLER_9_495 ();
 FILLCELL_X2 FILLER_9_507 ();
 FILLCELL_X16 FILLER_9_529 ();
 FILLCELL_X8 FILLER_9_545 ();
 FILLCELL_X1 FILLER_9_553 ();
 FILLCELL_X8 FILLER_9_568 ();
 FILLCELL_X4 FILLER_9_576 ();
 FILLCELL_X2 FILLER_9_580 ();
 FILLCELL_X1 FILLER_9_582 ();
 FILLCELL_X4 FILLER_9_612 ();
 FILLCELL_X2 FILLER_9_621 ();
 FILLCELL_X4 FILLER_9_629 ();
 FILLCELL_X1 FILLER_9_633 ();
 FILLCELL_X2 FILLER_9_657 ();
 FILLCELL_X2 FILLER_9_664 ();
 FILLCELL_X1 FILLER_9_666 ();
 FILLCELL_X2 FILLER_9_671 ();
 FILLCELL_X1 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_678 ();
 FILLCELL_X16 FILLER_9_710 ();
 FILLCELL_X4 FILLER_9_726 ();
 FILLCELL_X1 FILLER_9_730 ();
 FILLCELL_X8 FILLER_9_740 ();
 FILLCELL_X4 FILLER_9_748 ();
 FILLCELL_X2 FILLER_9_752 ();
 FILLCELL_X1 FILLER_9_754 ();
 FILLCELL_X4 FILLER_9_773 ();
 FILLCELL_X2 FILLER_9_817 ();
 FILLCELL_X4 FILLER_9_824 ();
 FILLCELL_X2 FILLER_9_828 ();
 FILLCELL_X4 FILLER_9_875 ();
 FILLCELL_X1 FILLER_9_883 ();
 FILLCELL_X8 FILLER_9_896 ();
 FILLCELL_X4 FILLER_9_904 ();
 FILLCELL_X8 FILLER_9_944 ();
 FILLCELL_X1 FILLER_9_952 ();
 FILLCELL_X4 FILLER_9_960 ();
 FILLCELL_X2 FILLER_9_964 ();
 FILLCELL_X1 FILLER_9_966 ();
 FILLCELL_X32 FILLER_9_971 ();
 FILLCELL_X32 FILLER_9_1003 ();
 FILLCELL_X4 FILLER_9_1035 ();
 FILLCELL_X1 FILLER_9_1039 ();
 FILLCELL_X1 FILLER_9_1047 ();
 FILLCELL_X2 FILLER_9_1053 ();
 FILLCELL_X2 FILLER_9_1064 ();
 FILLCELL_X2 FILLER_9_1084 ();
 FILLCELL_X2 FILLER_9_1091 ();
 FILLCELL_X8 FILLER_9_1106 ();
 FILLCELL_X4 FILLER_9_1114 ();
 FILLCELL_X2 FILLER_9_1118 ();
 FILLCELL_X1 FILLER_9_1120 ();
 FILLCELL_X1 FILLER_9_1175 ();
 FILLCELL_X2 FILLER_9_1179 ();
 FILLCELL_X4 FILLER_9_1188 ();
 FILLCELL_X4 FILLER_9_1196 ();
 FILLCELL_X1 FILLER_9_1200 ();
 FILLCELL_X4 FILLER_9_1208 ();
 FILLCELL_X1 FILLER_9_1212 ();
 FILLCELL_X4 FILLER_9_1226 ();
 FILLCELL_X16 FILLER_9_1235 ();
 FILLCELL_X8 FILLER_9_1251 ();
 FILLCELL_X4 FILLER_9_1259 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X32 FILLER_9_1296 ();
 FILLCELL_X32 FILLER_9_1328 ();
 FILLCELL_X32 FILLER_9_1360 ();
 FILLCELL_X32 FILLER_9_1392 ();
 FILLCELL_X32 FILLER_9_1424 ();
 FILLCELL_X32 FILLER_9_1456 ();
 FILLCELL_X32 FILLER_9_1488 ();
 FILLCELL_X32 FILLER_9_1520 ();
 FILLCELL_X32 FILLER_9_1552 ();
 FILLCELL_X32 FILLER_9_1584 ();
 FILLCELL_X32 FILLER_9_1616 ();
 FILLCELL_X2 FILLER_9_1648 ();
 FILLCELL_X1 FILLER_9_1650 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X16 FILLER_10_161 ();
 FILLCELL_X8 FILLER_10_177 ();
 FILLCELL_X1 FILLER_10_185 ();
 FILLCELL_X4 FILLER_10_197 ();
 FILLCELL_X1 FILLER_10_201 ();
 FILLCELL_X1 FILLER_10_211 ();
 FILLCELL_X8 FILLER_10_216 ();
 FILLCELL_X2 FILLER_10_224 ();
 FILLCELL_X4 FILLER_10_230 ();
 FILLCELL_X4 FILLER_10_249 ();
 FILLCELL_X8 FILLER_10_299 ();
 FILLCELL_X1 FILLER_10_307 ();
 FILLCELL_X4 FILLER_10_313 ();
 FILLCELL_X1 FILLER_10_324 ();
 FILLCELL_X1 FILLER_10_332 ();
 FILLCELL_X1 FILLER_10_342 ();
 FILLCELL_X1 FILLER_10_350 ();
 FILLCELL_X1 FILLER_10_362 ();
 FILLCELL_X2 FILLER_10_377 ();
 FILLCELL_X2 FILLER_10_390 ();
 FILLCELL_X4 FILLER_10_401 ();
 FILLCELL_X16 FILLER_10_423 ();
 FILLCELL_X8 FILLER_10_439 ();
 FILLCELL_X4 FILLER_10_447 ();
 FILLCELL_X2 FILLER_10_451 ();
 FILLCELL_X4 FILLER_10_465 ();
 FILLCELL_X2 FILLER_10_469 ();
 FILLCELL_X1 FILLER_10_471 ();
 FILLCELL_X1 FILLER_10_485 ();
 FILLCELL_X4 FILLER_10_497 ();
 FILLCELL_X1 FILLER_10_501 ();
 FILLCELL_X4 FILLER_10_506 ();
 FILLCELL_X1 FILLER_10_510 ();
 FILLCELL_X4 FILLER_10_518 ();
 FILLCELL_X1 FILLER_10_531 ();
 FILLCELL_X2 FILLER_10_555 ();
 FILLCELL_X4 FILLER_10_571 ();
 FILLCELL_X2 FILLER_10_575 ();
 FILLCELL_X2 FILLER_10_595 ();
 FILLCELL_X1 FILLER_10_597 ();
 FILLCELL_X8 FILLER_10_601 ();
 FILLCELL_X4 FILLER_10_609 ();
 FILLCELL_X1 FILLER_10_613 ();
 FILLCELL_X4 FILLER_10_619 ();
 FILLCELL_X2 FILLER_10_623 ();
 FILLCELL_X1 FILLER_10_625 ();
 FILLCELL_X1 FILLER_10_630 ();
 FILLCELL_X2 FILLER_10_632 ();
 FILLCELL_X2 FILLER_10_651 ();
 FILLCELL_X1 FILLER_10_653 ();
 FILLCELL_X2 FILLER_10_663 ();
 FILLCELL_X1 FILLER_10_665 ();
 FILLCELL_X4 FILLER_10_673 ();
 FILLCELL_X2 FILLER_10_680 ();
 FILLCELL_X32 FILLER_10_689 ();
 FILLCELL_X4 FILLER_10_721 ();
 FILLCELL_X2 FILLER_10_725 ();
 FILLCELL_X1 FILLER_10_727 ();
 FILLCELL_X4 FILLER_10_755 ();
 FILLCELL_X2 FILLER_10_759 ();
 FILLCELL_X1 FILLER_10_761 ();
 FILLCELL_X2 FILLER_10_769 ();
 FILLCELL_X1 FILLER_10_771 ();
 FILLCELL_X2 FILLER_10_775 ();
 FILLCELL_X2 FILLER_10_794 ();
 FILLCELL_X1 FILLER_10_796 ();
 FILLCELL_X4 FILLER_10_812 ();
 FILLCELL_X4 FILLER_10_840 ();
 FILLCELL_X1 FILLER_10_844 ();
 FILLCELL_X2 FILLER_10_867 ();
 FILLCELL_X2 FILLER_10_882 ();
 FILLCELL_X1 FILLER_10_884 ();
 FILLCELL_X4 FILLER_10_889 ();
 FILLCELL_X2 FILLER_10_915 ();
 FILLCELL_X1 FILLER_10_921 ();
 FILLCELL_X4 FILLER_10_941 ();
 FILLCELL_X1 FILLER_10_945 ();
 FILLCELL_X4 FILLER_10_953 ();
 FILLCELL_X4 FILLER_10_964 ();
 FILLCELL_X32 FILLER_10_972 ();
 FILLCELL_X8 FILLER_10_1004 ();
 FILLCELL_X4 FILLER_10_1012 ();
 FILLCELL_X2 FILLER_10_1016 ();
 FILLCELL_X8 FILLER_10_1027 ();
 FILLCELL_X8 FILLER_10_1042 ();
 FILLCELL_X4 FILLER_10_1050 ();
 FILLCELL_X2 FILLER_10_1054 ();
 FILLCELL_X8 FILLER_10_1072 ();
 FILLCELL_X1 FILLER_10_1080 ();
 FILLCELL_X16 FILLER_10_1100 ();
 FILLCELL_X4 FILLER_10_1116 ();
 FILLCELL_X2 FILLER_10_1120 ();
 FILLCELL_X1 FILLER_10_1131 ();
 FILLCELL_X2 FILLER_10_1139 ();
 FILLCELL_X1 FILLER_10_1141 ();
 FILLCELL_X1 FILLER_10_1153 ();
 FILLCELL_X1 FILLER_10_1158 ();
 FILLCELL_X2 FILLER_10_1180 ();
 FILLCELL_X8 FILLER_10_1186 ();
 FILLCELL_X1 FILLER_10_1194 ();
 FILLCELL_X1 FILLER_10_1199 ();
 FILLCELL_X1 FILLER_10_1207 ();
 FILLCELL_X1 FILLER_10_1223 ();
 FILLCELL_X32 FILLER_10_1257 ();
 FILLCELL_X32 FILLER_10_1289 ();
 FILLCELL_X32 FILLER_10_1321 ();
 FILLCELL_X32 FILLER_10_1353 ();
 FILLCELL_X32 FILLER_10_1385 ();
 FILLCELL_X32 FILLER_10_1417 ();
 FILLCELL_X32 FILLER_10_1449 ();
 FILLCELL_X32 FILLER_10_1481 ();
 FILLCELL_X32 FILLER_10_1513 ();
 FILLCELL_X32 FILLER_10_1545 ();
 FILLCELL_X32 FILLER_10_1577 ();
 FILLCELL_X32 FILLER_10_1609 ();
 FILLCELL_X8 FILLER_10_1641 ();
 FILLCELL_X2 FILLER_10_1649 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X16 FILLER_11_161 ();
 FILLCELL_X4 FILLER_11_184 ();
 FILLCELL_X2 FILLER_11_188 ();
 FILLCELL_X2 FILLER_11_216 ();
 FILLCELL_X1 FILLER_11_218 ();
 FILLCELL_X4 FILLER_11_230 ();
 FILLCELL_X2 FILLER_11_234 ();
 FILLCELL_X1 FILLER_11_236 ();
 FILLCELL_X8 FILLER_11_255 ();
 FILLCELL_X2 FILLER_11_263 ();
 FILLCELL_X2 FILLER_11_286 ();
 FILLCELL_X2 FILLER_11_299 ();
 FILLCELL_X1 FILLER_11_316 ();
 FILLCELL_X2 FILLER_11_344 ();
 FILLCELL_X2 FILLER_11_355 ();
 FILLCELL_X1 FILLER_11_366 ();
 FILLCELL_X4 FILLER_11_383 ();
 FILLCELL_X32 FILLER_11_394 ();
 FILLCELL_X16 FILLER_11_426 ();
 FILLCELL_X8 FILLER_11_442 ();
 FILLCELL_X4 FILLER_11_450 ();
 FILLCELL_X2 FILLER_11_454 ();
 FILLCELL_X1 FILLER_11_463 ();
 FILLCELL_X2 FILLER_11_468 ();
 FILLCELL_X1 FILLER_11_474 ();
 FILLCELL_X4 FILLER_11_500 ();
 FILLCELL_X4 FILLER_11_512 ();
 FILLCELL_X2 FILLER_11_516 ();
 FILLCELL_X1 FILLER_11_527 ();
 FILLCELL_X2 FILLER_11_533 ();
 FILLCELL_X1 FILLER_11_535 ();
 FILLCELL_X2 FILLER_11_541 ();
 FILLCELL_X1 FILLER_11_543 ();
 FILLCELL_X1 FILLER_11_548 ();
 FILLCELL_X8 FILLER_11_571 ();
 FILLCELL_X4 FILLER_11_579 ();
 FILLCELL_X2 FILLER_11_583 ();
 FILLCELL_X1 FILLER_11_585 ();
 FILLCELL_X8 FILLER_11_593 ();
 FILLCELL_X4 FILLER_11_618 ();
 FILLCELL_X16 FILLER_11_632 ();
 FILLCELL_X2 FILLER_11_648 ();
 FILLCELL_X8 FILLER_11_659 ();
 FILLCELL_X2 FILLER_11_667 ();
 FILLCELL_X2 FILLER_11_680 ();
 FILLCELL_X1 FILLER_11_682 ();
 FILLCELL_X4 FILLER_11_688 ();
 FILLCELL_X32 FILLER_11_699 ();
 FILLCELL_X4 FILLER_11_731 ();
 FILLCELL_X2 FILLER_11_759 ();
 FILLCELL_X2 FILLER_11_775 ();
 FILLCELL_X1 FILLER_11_777 ();
 FILLCELL_X2 FILLER_11_784 ();
 FILLCELL_X1 FILLER_11_786 ();
 FILLCELL_X2 FILLER_11_802 ();
 FILLCELL_X2 FILLER_11_808 ();
 FILLCELL_X1 FILLER_11_823 ();
 FILLCELL_X1 FILLER_11_834 ();
 FILLCELL_X4 FILLER_11_844 ();
 FILLCELL_X1 FILLER_11_848 ();
 FILLCELL_X4 FILLER_11_852 ();
 FILLCELL_X4 FILLER_11_864 ();
 FILLCELL_X8 FILLER_11_877 ();
 FILLCELL_X4 FILLER_11_885 ();
 FILLCELL_X16 FILLER_11_902 ();
 FILLCELL_X4 FILLER_11_918 ();
 FILLCELL_X1 FILLER_11_922 ();
 FILLCELL_X1 FILLER_11_934 ();
 FILLCELL_X1 FILLER_11_946 ();
 FILLCELL_X1 FILLER_11_958 ();
 FILLCELL_X1 FILLER_11_970 ();
 FILLCELL_X8 FILLER_11_978 ();
 FILLCELL_X16 FILLER_11_993 ();
 FILLCELL_X8 FILLER_11_1009 ();
 FILLCELL_X2 FILLER_11_1017 ();
 FILLCELL_X1 FILLER_11_1019 ();
 FILLCELL_X1 FILLER_11_1038 ();
 FILLCELL_X2 FILLER_11_1049 ();
 FILLCELL_X4 FILLER_11_1063 ();
 FILLCELL_X1 FILLER_11_1067 ();
 FILLCELL_X8 FILLER_11_1098 ();
 FILLCELL_X2 FILLER_11_1135 ();
 FILLCELL_X1 FILLER_11_1137 ();
 FILLCELL_X1 FILLER_11_1145 ();
 FILLCELL_X4 FILLER_11_1150 ();
 FILLCELL_X1 FILLER_11_1154 ();
 FILLCELL_X4 FILLER_11_1158 ();
 FILLCELL_X2 FILLER_11_1162 ();
 FILLCELL_X4 FILLER_11_1170 ();
 FILLCELL_X2 FILLER_11_1174 ();
 FILLCELL_X8 FILLER_11_1180 ();
 FILLCELL_X1 FILLER_11_1188 ();
 FILLCELL_X4 FILLER_11_1203 ();
 FILLCELL_X2 FILLER_11_1215 ();
 FILLCELL_X1 FILLER_11_1217 ();
 FILLCELL_X1 FILLER_11_1221 ();
 FILLCELL_X1 FILLER_11_1229 ();
 FILLCELL_X8 FILLER_11_1235 ();
 FILLCELL_X2 FILLER_11_1243 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1257 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X32 FILLER_11_1296 ();
 FILLCELL_X32 FILLER_11_1328 ();
 FILLCELL_X32 FILLER_11_1360 ();
 FILLCELL_X32 FILLER_11_1392 ();
 FILLCELL_X32 FILLER_11_1424 ();
 FILLCELL_X32 FILLER_11_1456 ();
 FILLCELL_X32 FILLER_11_1488 ();
 FILLCELL_X32 FILLER_11_1520 ();
 FILLCELL_X32 FILLER_11_1552 ();
 FILLCELL_X32 FILLER_11_1584 ();
 FILLCELL_X32 FILLER_11_1616 ();
 FILLCELL_X2 FILLER_11_1648 ();
 FILLCELL_X1 FILLER_11_1650 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X2 FILLER_12_193 ();
 FILLCELL_X8 FILLER_12_205 ();
 FILLCELL_X4 FILLER_12_213 ();
 FILLCELL_X1 FILLER_12_259 ();
 FILLCELL_X4 FILLER_12_284 ();
 FILLCELL_X2 FILLER_12_288 ();
 FILLCELL_X1 FILLER_12_301 ();
 FILLCELL_X8 FILLER_12_307 ();
 FILLCELL_X4 FILLER_12_315 ();
 FILLCELL_X2 FILLER_12_339 ();
 FILLCELL_X1 FILLER_12_341 ();
 FILLCELL_X32 FILLER_12_358 ();
 FILLCELL_X2 FILLER_12_390 ();
 FILLCELL_X1 FILLER_12_392 ();
 FILLCELL_X8 FILLER_12_427 ();
 FILLCELL_X4 FILLER_12_435 ();
 FILLCELL_X2 FILLER_12_439 ();
 FILLCELL_X1 FILLER_12_441 ();
 FILLCELL_X2 FILLER_12_460 ();
 FILLCELL_X1 FILLER_12_462 ();
 FILLCELL_X2 FILLER_12_493 ();
 FILLCELL_X1 FILLER_12_495 ();
 FILLCELL_X4 FILLER_12_503 ();
 FILLCELL_X1 FILLER_12_534 ();
 FILLCELL_X1 FILLER_12_540 ();
 FILLCELL_X1 FILLER_12_557 ();
 FILLCELL_X8 FILLER_12_584 ();
 FILLCELL_X4 FILLER_12_592 ();
 FILLCELL_X8 FILLER_12_603 ();
 FILLCELL_X1 FILLER_12_616 ();
 FILLCELL_X2 FILLER_12_668 ();
 FILLCELL_X1 FILLER_12_670 ();
 FILLCELL_X32 FILLER_12_678 ();
 FILLCELL_X16 FILLER_12_710 ();
 FILLCELL_X8 FILLER_12_726 ();
 FILLCELL_X4 FILLER_12_734 ();
 FILLCELL_X2 FILLER_12_738 ();
 FILLCELL_X4 FILLER_12_758 ();
 FILLCELL_X2 FILLER_12_762 ();
 FILLCELL_X1 FILLER_12_764 ();
 FILLCELL_X4 FILLER_12_787 ();
 FILLCELL_X1 FILLER_12_791 ();
 FILLCELL_X2 FILLER_12_799 ();
 FILLCELL_X2 FILLER_12_806 ();
 FILLCELL_X1 FILLER_12_815 ();
 FILLCELL_X1 FILLER_12_819 ();
 FILLCELL_X4 FILLER_12_824 ();
 FILLCELL_X1 FILLER_12_828 ();
 FILLCELL_X2 FILLER_12_886 ();
 FILLCELL_X8 FILLER_12_899 ();
 FILLCELL_X2 FILLER_12_907 ();
 FILLCELL_X8 FILLER_12_921 ();
 FILLCELL_X4 FILLER_12_929 ();
 FILLCELL_X4 FILLER_12_979 ();
 FILLCELL_X2 FILLER_12_1001 ();
 FILLCELL_X2 FILLER_12_1010 ();
 FILLCELL_X1 FILLER_12_1012 ();
 FILLCELL_X4 FILLER_12_1056 ();
 FILLCELL_X4 FILLER_12_1069 ();
 FILLCELL_X2 FILLER_12_1080 ();
 FILLCELL_X8 FILLER_12_1095 ();
 FILLCELL_X1 FILLER_12_1103 ();
 FILLCELL_X4 FILLER_12_1133 ();
 FILLCELL_X2 FILLER_12_1148 ();
 FILLCELL_X1 FILLER_12_1150 ();
 FILLCELL_X1 FILLER_12_1158 ();
 FILLCELL_X2 FILLER_12_1178 ();
 FILLCELL_X1 FILLER_12_1180 ();
 FILLCELL_X8 FILLER_12_1204 ();
 FILLCELL_X4 FILLER_12_1212 ();
 FILLCELL_X2 FILLER_12_1235 ();
 FILLCELL_X1 FILLER_12_1237 ();
 FILLCELL_X32 FILLER_12_1255 ();
 FILLCELL_X32 FILLER_12_1287 ();
 FILLCELL_X32 FILLER_12_1319 ();
 FILLCELL_X32 FILLER_12_1351 ();
 FILLCELL_X32 FILLER_12_1383 ();
 FILLCELL_X32 FILLER_12_1415 ();
 FILLCELL_X32 FILLER_12_1447 ();
 FILLCELL_X32 FILLER_12_1479 ();
 FILLCELL_X32 FILLER_12_1511 ();
 FILLCELL_X32 FILLER_12_1543 ();
 FILLCELL_X32 FILLER_12_1575 ();
 FILLCELL_X32 FILLER_12_1607 ();
 FILLCELL_X8 FILLER_12_1639 ();
 FILLCELL_X4 FILLER_12_1647 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X16 FILLER_13_161 ();
 FILLCELL_X2 FILLER_13_177 ();
 FILLCELL_X1 FILLER_13_179 ();
 FILLCELL_X4 FILLER_13_198 ();
 FILLCELL_X2 FILLER_13_219 ();
 FILLCELL_X2 FILLER_13_239 ();
 FILLCELL_X1 FILLER_13_277 ();
 FILLCELL_X2 FILLER_13_291 ();
 FILLCELL_X1 FILLER_13_302 ();
 FILLCELL_X1 FILLER_13_321 ();
 FILLCELL_X1 FILLER_13_333 ();
 FILLCELL_X2 FILLER_13_338 ();
 FILLCELL_X4 FILLER_13_344 ();
 FILLCELL_X1 FILLER_13_348 ();
 FILLCELL_X4 FILLER_13_352 ();
 FILLCELL_X1 FILLER_13_356 ();
 FILLCELL_X2 FILLER_13_371 ();
 FILLCELL_X8 FILLER_13_391 ();
 FILLCELL_X4 FILLER_13_399 ();
 FILLCELL_X1 FILLER_13_403 ();
 FILLCELL_X32 FILLER_13_422 ();
 FILLCELL_X4 FILLER_13_454 ();
 FILLCELL_X1 FILLER_13_458 ();
 FILLCELL_X2 FILLER_13_471 ();
 FILLCELL_X1 FILLER_13_473 ();
 FILLCELL_X8 FILLER_13_477 ();
 FILLCELL_X4 FILLER_13_485 ();
 FILLCELL_X1 FILLER_13_489 ();
 FILLCELL_X4 FILLER_13_494 ();
 FILLCELL_X2 FILLER_13_498 ();
 FILLCELL_X4 FILLER_13_507 ();
 FILLCELL_X4 FILLER_13_518 ();
 FILLCELL_X2 FILLER_13_540 ();
 FILLCELL_X16 FILLER_13_557 ();
 FILLCELL_X4 FILLER_13_573 ();
 FILLCELL_X2 FILLER_13_617 ();
 FILLCELL_X1 FILLER_13_619 ();
 FILLCELL_X8 FILLER_13_631 ();
 FILLCELL_X2 FILLER_13_639 ();
 FILLCELL_X1 FILLER_13_641 ();
 FILLCELL_X4 FILLER_13_649 ();
 FILLCELL_X2 FILLER_13_653 ();
 FILLCELL_X1 FILLER_13_666 ();
 FILLCELL_X4 FILLER_13_674 ();
 FILLCELL_X2 FILLER_13_678 ();
 FILLCELL_X4 FILLER_13_684 ();
 FILLCELL_X1 FILLER_13_688 ();
 FILLCELL_X32 FILLER_13_695 ();
 FILLCELL_X8 FILLER_13_727 ();
 FILLCELL_X2 FILLER_13_735 ();
 FILLCELL_X1 FILLER_13_737 ();
 FILLCELL_X4 FILLER_13_763 ();
 FILLCELL_X2 FILLER_13_767 ();
 FILLCELL_X1 FILLER_13_769 ();
 FILLCELL_X8 FILLER_13_792 ();
 FILLCELL_X2 FILLER_13_800 ();
 FILLCELL_X1 FILLER_13_802 ();
 FILLCELL_X8 FILLER_13_807 ();
 FILLCELL_X8 FILLER_13_820 ();
 FILLCELL_X2 FILLER_13_828 ();
 FILLCELL_X16 FILLER_13_841 ();
 FILLCELL_X4 FILLER_13_857 ();
 FILLCELL_X4 FILLER_13_865 ();
 FILLCELL_X8 FILLER_13_876 ();
 FILLCELL_X2 FILLER_13_884 ();
 FILLCELL_X2 FILLER_13_889 ();
 FILLCELL_X2 FILLER_13_899 ();
 FILLCELL_X2 FILLER_13_908 ();
 FILLCELL_X8 FILLER_13_915 ();
 FILLCELL_X16 FILLER_13_932 ();
 FILLCELL_X8 FILLER_13_948 ();
 FILLCELL_X1 FILLER_13_960 ();
 FILLCELL_X4 FILLER_13_982 ();
 FILLCELL_X2 FILLER_13_1006 ();
 FILLCELL_X1 FILLER_13_1008 ();
 FILLCELL_X4 FILLER_13_1014 ();
 FILLCELL_X1 FILLER_13_1018 ();
 FILLCELL_X4 FILLER_13_1024 ();
 FILLCELL_X1 FILLER_13_1028 ();
 FILLCELL_X2 FILLER_13_1047 ();
 FILLCELL_X1 FILLER_13_1049 ();
 FILLCELL_X1 FILLER_13_1057 ();
 FILLCELL_X1 FILLER_13_1065 ();
 FILLCELL_X2 FILLER_13_1080 ();
 FILLCELL_X4 FILLER_13_1089 ();
 FILLCELL_X4 FILLER_13_1097 ();
 FILLCELL_X4 FILLER_13_1108 ();
 FILLCELL_X2 FILLER_13_1124 ();
 FILLCELL_X1 FILLER_13_1129 ();
 FILLCELL_X2 FILLER_13_1133 ();
 FILLCELL_X2 FILLER_13_1139 ();
 FILLCELL_X2 FILLER_13_1148 ();
 FILLCELL_X1 FILLER_13_1150 ();
 FILLCELL_X8 FILLER_13_1155 ();
 FILLCELL_X2 FILLER_13_1163 ();
 FILLCELL_X2 FILLER_13_1171 ();
 FILLCELL_X1 FILLER_13_1173 ();
 FILLCELL_X8 FILLER_13_1190 ();
 FILLCELL_X2 FILLER_13_1198 ();
 FILLCELL_X4 FILLER_13_1231 ();
 FILLCELL_X1 FILLER_13_1235 ();
 FILLCELL_X1 FILLER_13_1240 ();
 FILLCELL_X4 FILLER_13_1245 ();
 FILLCELL_X1 FILLER_13_1249 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X32 FILLER_13_1296 ();
 FILLCELL_X32 FILLER_13_1328 ();
 FILLCELL_X32 FILLER_13_1360 ();
 FILLCELL_X32 FILLER_13_1392 ();
 FILLCELL_X32 FILLER_13_1424 ();
 FILLCELL_X32 FILLER_13_1456 ();
 FILLCELL_X32 FILLER_13_1488 ();
 FILLCELL_X32 FILLER_13_1520 ();
 FILLCELL_X32 FILLER_13_1552 ();
 FILLCELL_X32 FILLER_13_1584 ();
 FILLCELL_X32 FILLER_13_1616 ();
 FILLCELL_X2 FILLER_13_1648 ();
 FILLCELL_X1 FILLER_13_1650 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X16 FILLER_14_161 ();
 FILLCELL_X4 FILLER_14_177 ();
 FILLCELL_X1 FILLER_14_197 ();
 FILLCELL_X2 FILLER_14_212 ();
 FILLCELL_X8 FILLER_14_218 ();
 FILLCELL_X4 FILLER_14_226 ();
 FILLCELL_X2 FILLER_14_230 ();
 FILLCELL_X2 FILLER_14_241 ();
 FILLCELL_X1 FILLER_14_243 ();
 FILLCELL_X4 FILLER_14_249 ();
 FILLCELL_X1 FILLER_14_253 ();
 FILLCELL_X4 FILLER_14_257 ();
 FILLCELL_X2 FILLER_14_261 ();
 FILLCELL_X1 FILLER_14_263 ();
 FILLCELL_X8 FILLER_14_268 ();
 FILLCELL_X4 FILLER_14_292 ();
 FILLCELL_X1 FILLER_14_300 ();
 FILLCELL_X1 FILLER_14_305 ();
 FILLCELL_X8 FILLER_14_309 ();
 FILLCELL_X4 FILLER_14_317 ();
 FILLCELL_X2 FILLER_14_321 ();
 FILLCELL_X1 FILLER_14_323 ();
 FILLCELL_X2 FILLER_14_331 ();
 FILLCELL_X4 FILLER_14_337 ();
 FILLCELL_X2 FILLER_14_344 ();
 FILLCELL_X1 FILLER_14_346 ();
 FILLCELL_X1 FILLER_14_369 ();
 FILLCELL_X1 FILLER_14_374 ();
 FILLCELL_X1 FILLER_14_382 ();
 FILLCELL_X1 FILLER_14_392 ();
 FILLCELL_X2 FILLER_14_400 ();
 FILLCELL_X32 FILLER_14_428 ();
 FILLCELL_X1 FILLER_14_460 ();
 FILLCELL_X8 FILLER_14_479 ();
 FILLCELL_X2 FILLER_14_487 ();
 FILLCELL_X1 FILLER_14_503 ();
 FILLCELL_X4 FILLER_14_508 ();
 FILLCELL_X2 FILLER_14_516 ();
 FILLCELL_X1 FILLER_14_518 ();
 FILLCELL_X2 FILLER_14_528 ();
 FILLCELL_X1 FILLER_14_530 ();
 FILLCELL_X4 FILLER_14_534 ();
 FILLCELL_X1 FILLER_14_538 ();
 FILLCELL_X1 FILLER_14_567 ();
 FILLCELL_X2 FILLER_14_577 ();
 FILLCELL_X1 FILLER_14_579 ();
 FILLCELL_X2 FILLER_14_585 ();
 FILLCELL_X8 FILLER_14_596 ();
 FILLCELL_X4 FILLER_14_604 ();
 FILLCELL_X1 FILLER_14_613 ();
 FILLCELL_X1 FILLER_14_621 ();
 FILLCELL_X4 FILLER_14_686 ();
 FILLCELL_X2 FILLER_14_690 ();
 FILLCELL_X2 FILLER_14_710 ();
 FILLCELL_X1 FILLER_14_712 ();
 FILLCELL_X4 FILLER_14_757 ();
 FILLCELL_X8 FILLER_14_765 ();
 FILLCELL_X4 FILLER_14_777 ();
 FILLCELL_X1 FILLER_14_781 ();
 FILLCELL_X4 FILLER_14_789 ();
 FILLCELL_X1 FILLER_14_793 ();
 FILLCELL_X2 FILLER_14_798 ();
 FILLCELL_X1 FILLER_14_800 ();
 FILLCELL_X1 FILLER_14_810 ();
 FILLCELL_X8 FILLER_14_820 ();
 FILLCELL_X2 FILLER_14_828 ();
 FILLCELL_X1 FILLER_14_830 ();
 FILLCELL_X8 FILLER_14_843 ();
 FILLCELL_X2 FILLER_14_851 ();
 FILLCELL_X1 FILLER_14_853 ();
 FILLCELL_X4 FILLER_14_866 ();
 FILLCELL_X1 FILLER_14_877 ();
 FILLCELL_X2 FILLER_14_881 ();
 FILLCELL_X8 FILLER_14_896 ();
 FILLCELL_X4 FILLER_14_904 ();
 FILLCELL_X1 FILLER_14_908 ();
 FILLCELL_X4 FILLER_14_913 ();
 FILLCELL_X2 FILLER_14_917 ();
 FILLCELL_X8 FILLER_14_923 ();
 FILLCELL_X2 FILLER_14_931 ();
 FILLCELL_X2 FILLER_14_945 ();
 FILLCELL_X1 FILLER_14_947 ();
 FILLCELL_X1 FILLER_14_956 ();
 FILLCELL_X32 FILLER_14_968 ();
 FILLCELL_X2 FILLER_14_1000 ();
 FILLCELL_X16 FILLER_14_1013 ();
 FILLCELL_X8 FILLER_14_1029 ();
 FILLCELL_X16 FILLER_14_1046 ();
 FILLCELL_X2 FILLER_14_1062 ();
 FILLCELL_X1 FILLER_14_1084 ();
 FILLCELL_X16 FILLER_14_1094 ();
 FILLCELL_X2 FILLER_14_1110 ();
 FILLCELL_X1 FILLER_14_1112 ();
 FILLCELL_X1 FILLER_14_1152 ();
 FILLCELL_X1 FILLER_14_1171 ();
 FILLCELL_X1 FILLER_14_1176 ();
 FILLCELL_X1 FILLER_14_1184 ();
 FILLCELL_X2 FILLER_14_1191 ();
 FILLCELL_X1 FILLER_14_1193 ();
 FILLCELL_X2 FILLER_14_1200 ();
 FILLCELL_X2 FILLER_14_1211 ();
 FILLCELL_X2 FILLER_14_1235 ();
 FILLCELL_X2 FILLER_14_1257 ();
 FILLCELL_X1 FILLER_14_1259 ();
 FILLCELL_X32 FILLER_14_1267 ();
 FILLCELL_X32 FILLER_14_1299 ();
 FILLCELL_X32 FILLER_14_1331 ();
 FILLCELL_X16 FILLER_14_1363 ();
 FILLCELL_X2 FILLER_14_1379 ();
 FILLCELL_X8 FILLER_14_1391 ();
 FILLCELL_X32 FILLER_14_1406 ();
 FILLCELL_X32 FILLER_14_1438 ();
 FILLCELL_X32 FILLER_14_1470 ();
 FILLCELL_X32 FILLER_14_1502 ();
 FILLCELL_X32 FILLER_14_1534 ();
 FILLCELL_X32 FILLER_14_1566 ();
 FILLCELL_X32 FILLER_14_1598 ();
 FILLCELL_X16 FILLER_14_1630 ();
 FILLCELL_X4 FILLER_14_1646 ();
 FILLCELL_X1 FILLER_14_1650 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_161 ();
 FILLCELL_X4 FILLER_15_169 ();
 FILLCELL_X2 FILLER_15_173 ();
 FILLCELL_X1 FILLER_15_185 ();
 FILLCELL_X1 FILLER_15_191 ();
 FILLCELL_X1 FILLER_15_196 ();
 FILLCELL_X1 FILLER_15_202 ();
 FILLCELL_X1 FILLER_15_213 ();
 FILLCELL_X8 FILLER_15_219 ();
 FILLCELL_X1 FILLER_15_227 ();
 FILLCELL_X1 FILLER_15_244 ();
 FILLCELL_X8 FILLER_15_257 ();
 FILLCELL_X2 FILLER_15_265 ();
 FILLCELL_X1 FILLER_15_267 ();
 FILLCELL_X8 FILLER_15_273 ();
 FILLCELL_X2 FILLER_15_285 ();
 FILLCELL_X2 FILLER_15_296 ();
 FILLCELL_X1 FILLER_15_298 ();
 FILLCELL_X2 FILLER_15_315 ();
 FILLCELL_X16 FILLER_15_328 ();
 FILLCELL_X8 FILLER_15_396 ();
 FILLCELL_X2 FILLER_15_404 ();
 FILLCELL_X1 FILLER_15_406 ();
 FILLCELL_X32 FILLER_15_438 ();
 FILLCELL_X16 FILLER_15_474 ();
 FILLCELL_X2 FILLER_15_490 ();
 FILLCELL_X1 FILLER_15_492 ();
 FILLCELL_X4 FILLER_15_498 ();
 FILLCELL_X4 FILLER_15_514 ();
 FILLCELL_X2 FILLER_15_518 ();
 FILLCELL_X1 FILLER_15_528 ();
 FILLCELL_X2 FILLER_15_533 ();
 FILLCELL_X1 FILLER_15_535 ();
 FILLCELL_X1 FILLER_15_582 ();
 FILLCELL_X4 FILLER_15_600 ();
 FILLCELL_X2 FILLER_15_604 ();
 FILLCELL_X8 FILLER_15_613 ();
 FILLCELL_X2 FILLER_15_621 ();
 FILLCELL_X1 FILLER_15_630 ();
 FILLCELL_X4 FILLER_15_638 ();
 FILLCELL_X2 FILLER_15_642 ();
 FILLCELL_X1 FILLER_15_644 ();
 FILLCELL_X8 FILLER_15_656 ();
 FILLCELL_X1 FILLER_15_664 ();
 FILLCELL_X32 FILLER_15_681 ();
 FILLCELL_X16 FILLER_15_713 ();
 FILLCELL_X4 FILLER_15_729 ();
 FILLCELL_X2 FILLER_15_733 ();
 FILLCELL_X2 FILLER_15_740 ();
 FILLCELL_X1 FILLER_15_742 ();
 FILLCELL_X1 FILLER_15_761 ();
 FILLCELL_X2 FILLER_15_788 ();
 FILLCELL_X1 FILLER_15_793 ();
 FILLCELL_X4 FILLER_15_798 ();
 FILLCELL_X1 FILLER_15_802 ();
 FILLCELL_X1 FILLER_15_819 ();
 FILLCELL_X1 FILLER_15_829 ();
 FILLCELL_X1 FILLER_15_841 ();
 FILLCELL_X2 FILLER_15_860 ();
 FILLCELL_X1 FILLER_15_866 ();
 FILLCELL_X2 FILLER_15_884 ();
 FILLCELL_X8 FILLER_15_895 ();
 FILLCELL_X1 FILLER_15_903 ();
 FILLCELL_X1 FILLER_15_937 ();
 FILLCELL_X1 FILLER_15_941 ();
 FILLCELL_X1 FILLER_15_953 ();
 FILLCELL_X32 FILLER_15_958 ();
 FILLCELL_X4 FILLER_15_990 ();
 FILLCELL_X2 FILLER_15_1018 ();
 FILLCELL_X4 FILLER_15_1029 ();
 FILLCELL_X2 FILLER_15_1060 ();
 FILLCELL_X1 FILLER_15_1062 ();
 FILLCELL_X2 FILLER_15_1066 ();
 FILLCELL_X4 FILLER_15_1090 ();
 FILLCELL_X2 FILLER_15_1098 ();
 FILLCELL_X1 FILLER_15_1104 ();
 FILLCELL_X1 FILLER_15_1112 ();
 FILLCELL_X1 FILLER_15_1117 ();
 FILLCELL_X8 FILLER_15_1123 ();
 FILLCELL_X4 FILLER_15_1131 ();
 FILLCELL_X2 FILLER_15_1135 ();
 FILLCELL_X1 FILLER_15_1137 ();
 FILLCELL_X16 FILLER_15_1158 ();
 FILLCELL_X8 FILLER_15_1174 ();
 FILLCELL_X1 FILLER_15_1182 ();
 FILLCELL_X16 FILLER_15_1194 ();
 FILLCELL_X2 FILLER_15_1227 ();
 FILLCELL_X1 FILLER_15_1247 ();
 FILLCELL_X8 FILLER_15_1255 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X8 FILLER_15_1296 ();
 FILLCELL_X2 FILLER_15_1304 ();
 FILLCELL_X1 FILLER_15_1306 ();
 FILLCELL_X2 FILLER_15_1312 ();
 FILLCELL_X1 FILLER_15_1317 ();
 FILLCELL_X4 FILLER_15_1340 ();
 FILLCELL_X2 FILLER_15_1344 ();
 FILLCELL_X8 FILLER_15_1350 ();
 FILLCELL_X8 FILLER_15_1362 ();
 FILLCELL_X4 FILLER_15_1370 ();
 FILLCELL_X2 FILLER_15_1374 ();
 FILLCELL_X1 FILLER_15_1379 ();
 FILLCELL_X2 FILLER_15_1396 ();
 FILLCELL_X4 FILLER_15_1401 ();
 FILLCELL_X1 FILLER_15_1405 ();
 FILLCELL_X4 FILLER_15_1413 ();
 FILLCELL_X2 FILLER_15_1417 ();
 FILLCELL_X1 FILLER_15_1419 ();
 FILLCELL_X2 FILLER_15_1424 ();
 FILLCELL_X32 FILLER_15_1431 ();
 FILLCELL_X32 FILLER_15_1463 ();
 FILLCELL_X32 FILLER_15_1495 ();
 FILLCELL_X32 FILLER_15_1527 ();
 FILLCELL_X32 FILLER_15_1559 ();
 FILLCELL_X32 FILLER_15_1591 ();
 FILLCELL_X16 FILLER_15_1623 ();
 FILLCELL_X8 FILLER_15_1639 ();
 FILLCELL_X4 FILLER_15_1647 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X2 FILLER_16_161 ();
 FILLCELL_X1 FILLER_16_163 ();
 FILLCELL_X1 FILLER_16_171 ();
 FILLCELL_X1 FILLER_16_176 ();
 FILLCELL_X1 FILLER_16_184 ();
 FILLCELL_X2 FILLER_16_191 ();
 FILLCELL_X1 FILLER_16_193 ();
 FILLCELL_X2 FILLER_16_199 ();
 FILLCELL_X8 FILLER_16_212 ();
 FILLCELL_X4 FILLER_16_220 ();
 FILLCELL_X2 FILLER_16_224 ();
 FILLCELL_X2 FILLER_16_233 ();
 FILLCELL_X2 FILLER_16_239 ();
 FILLCELL_X1 FILLER_16_241 ();
 FILLCELL_X2 FILLER_16_249 ();
 FILLCELL_X1 FILLER_16_251 ();
 FILLCELL_X2 FILLER_16_264 ();
 FILLCELL_X1 FILLER_16_266 ();
 FILLCELL_X4 FILLER_16_283 ();
 FILLCELL_X2 FILLER_16_287 ();
 FILLCELL_X1 FILLER_16_319 ();
 FILLCELL_X2 FILLER_16_325 ();
 FILLCELL_X8 FILLER_16_334 ();
 FILLCELL_X1 FILLER_16_342 ();
 FILLCELL_X4 FILLER_16_348 ();
 FILLCELL_X2 FILLER_16_352 ();
 FILLCELL_X1 FILLER_16_354 ();
 FILLCELL_X2 FILLER_16_362 ();
 FILLCELL_X4 FILLER_16_381 ();
 FILLCELL_X16 FILLER_16_392 ();
 FILLCELL_X2 FILLER_16_408 ();
 FILLCELL_X16 FILLER_16_430 ();
 FILLCELL_X8 FILLER_16_446 ();
 FILLCELL_X4 FILLER_16_454 ();
 FILLCELL_X8 FILLER_16_467 ();
 FILLCELL_X1 FILLER_16_475 ();
 FILLCELL_X4 FILLER_16_486 ();
 FILLCELL_X1 FILLER_16_490 ();
 FILLCELL_X4 FILLER_16_500 ();
 FILLCELL_X8 FILLER_16_512 ();
 FILLCELL_X16 FILLER_16_534 ();
 FILLCELL_X1 FILLER_16_550 ();
 FILLCELL_X4 FILLER_16_569 ();
 FILLCELL_X1 FILLER_16_573 ();
 FILLCELL_X2 FILLER_16_588 ();
 FILLCELL_X8 FILLER_16_597 ();
 FILLCELL_X2 FILLER_16_605 ();
 FILLCELL_X1 FILLER_16_630 ();
 FILLCELL_X4 FILLER_16_632 ();
 FILLCELL_X2 FILLER_16_636 ();
 FILLCELL_X1 FILLER_16_638 ();
 FILLCELL_X2 FILLER_16_648 ();
 FILLCELL_X1 FILLER_16_664 ();
 FILLCELL_X8 FILLER_16_672 ();
 FILLCELL_X1 FILLER_16_680 ();
 FILLCELL_X32 FILLER_16_698 ();
 FILLCELL_X16 FILLER_16_730 ();
 FILLCELL_X2 FILLER_16_746 ();
 FILLCELL_X8 FILLER_16_752 ();
 FILLCELL_X2 FILLER_16_760 ();
 FILLCELL_X1 FILLER_16_762 ();
 FILLCELL_X4 FILLER_16_769 ();
 FILLCELL_X8 FILLER_16_780 ();
 FILLCELL_X1 FILLER_16_799 ();
 FILLCELL_X1 FILLER_16_804 ();
 FILLCELL_X1 FILLER_16_815 ();
 FILLCELL_X2 FILLER_16_827 ();
 FILLCELL_X1 FILLER_16_829 ();
 FILLCELL_X2 FILLER_16_851 ();
 FILLCELL_X16 FILLER_16_862 ();
 FILLCELL_X1 FILLER_16_878 ();
 FILLCELL_X16 FILLER_16_891 ();
 FILLCELL_X4 FILLER_16_916 ();
 FILLCELL_X1 FILLER_16_920 ();
 FILLCELL_X1 FILLER_16_925 ();
 FILLCELL_X2 FILLER_16_931 ();
 FILLCELL_X1 FILLER_16_937 ();
 FILLCELL_X2 FILLER_16_947 ();
 FILLCELL_X1 FILLER_16_961 ();
 FILLCELL_X8 FILLER_16_979 ();
 FILLCELL_X4 FILLER_16_987 ();
 FILLCELL_X2 FILLER_16_991 ();
 FILLCELL_X2 FILLER_16_1027 ();
 FILLCELL_X4 FILLER_16_1038 ();
 FILLCELL_X1 FILLER_16_1042 ();
 FILLCELL_X1 FILLER_16_1059 ();
 FILLCELL_X2 FILLER_16_1080 ();
 FILLCELL_X8 FILLER_16_1100 ();
 FILLCELL_X2 FILLER_16_1108 ();
 FILLCELL_X8 FILLER_16_1128 ();
 FILLCELL_X1 FILLER_16_1136 ();
 FILLCELL_X8 FILLER_16_1142 ();
 FILLCELL_X8 FILLER_16_1171 ();
 FILLCELL_X2 FILLER_16_1179 ();
 FILLCELL_X1 FILLER_16_1181 ();
 FILLCELL_X8 FILLER_16_1193 ();
 FILLCELL_X2 FILLER_16_1201 ();
 FILLCELL_X4 FILLER_16_1206 ();
 FILLCELL_X2 FILLER_16_1219 ();
 FILLCELL_X1 FILLER_16_1221 ();
 FILLCELL_X4 FILLER_16_1233 ();
 FILLCELL_X1 FILLER_16_1237 ();
 FILLCELL_X32 FILLER_16_1243 ();
 FILLCELL_X16 FILLER_16_1275 ();
 FILLCELL_X8 FILLER_16_1291 ();
 FILLCELL_X2 FILLER_16_1299 ();
 FILLCELL_X1 FILLER_16_1301 ();
 FILLCELL_X1 FILLER_16_1322 ();
 FILLCELL_X1 FILLER_16_1334 ();
 FILLCELL_X4 FILLER_16_1349 ();
 FILLCELL_X4 FILLER_16_1373 ();
 FILLCELL_X2 FILLER_16_1377 ();
 FILLCELL_X1 FILLER_16_1379 ();
 FILLCELL_X4 FILLER_16_1385 ();
 FILLCELL_X1 FILLER_16_1389 ();
 FILLCELL_X8 FILLER_16_1397 ();
 FILLCELL_X2 FILLER_16_1405 ();
 FILLCELL_X2 FILLER_16_1418 ();
 FILLCELL_X16 FILLER_16_1424 ();
 FILLCELL_X1 FILLER_16_1440 ();
 FILLCELL_X32 FILLER_16_1448 ();
 FILLCELL_X32 FILLER_16_1480 ();
 FILLCELL_X32 FILLER_16_1512 ();
 FILLCELL_X32 FILLER_16_1544 ();
 FILLCELL_X32 FILLER_16_1576 ();
 FILLCELL_X32 FILLER_16_1608 ();
 FILLCELL_X8 FILLER_16_1640 ();
 FILLCELL_X2 FILLER_16_1648 ();
 FILLCELL_X1 FILLER_16_1650 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X4 FILLER_17_161 ();
 FILLCELL_X2 FILLER_17_193 ();
 FILLCELL_X2 FILLER_17_236 ();
 FILLCELL_X2 FILLER_17_247 ();
 FILLCELL_X1 FILLER_17_249 ();
 FILLCELL_X1 FILLER_17_273 ();
 FILLCELL_X1 FILLER_17_285 ();
 FILLCELL_X4 FILLER_17_293 ();
 FILLCELL_X2 FILLER_17_297 ();
 FILLCELL_X1 FILLER_17_314 ();
 FILLCELL_X8 FILLER_17_326 ();
 FILLCELL_X1 FILLER_17_334 ();
 FILLCELL_X1 FILLER_17_346 ();
 FILLCELL_X1 FILLER_17_354 ();
 FILLCELL_X1 FILLER_17_364 ();
 FILLCELL_X8 FILLER_17_368 ();
 FILLCELL_X2 FILLER_17_376 ();
 FILLCELL_X1 FILLER_17_387 ();
 FILLCELL_X32 FILLER_17_398 ();
 FILLCELL_X2 FILLER_17_430 ();
 FILLCELL_X1 FILLER_17_432 ();
 FILLCELL_X32 FILLER_17_436 ();
 FILLCELL_X4 FILLER_17_468 ();
 FILLCELL_X2 FILLER_17_472 ();
 FILLCELL_X1 FILLER_17_474 ();
 FILLCELL_X4 FILLER_17_493 ();
 FILLCELL_X1 FILLER_17_497 ();
 FILLCELL_X2 FILLER_17_516 ();
 FILLCELL_X4 FILLER_17_521 ();
 FILLCELL_X1 FILLER_17_525 ();
 FILLCELL_X2 FILLER_17_535 ();
 FILLCELL_X1 FILLER_17_537 ();
 FILLCELL_X2 FILLER_17_554 ();
 FILLCELL_X2 FILLER_17_580 ();
 FILLCELL_X4 FILLER_17_586 ();
 FILLCELL_X2 FILLER_17_590 ();
 FILLCELL_X1 FILLER_17_592 ();
 FILLCELL_X8 FILLER_17_600 ();
 FILLCELL_X2 FILLER_17_608 ();
 FILLCELL_X1 FILLER_17_610 ();
 FILLCELL_X1 FILLER_17_625 ();
 FILLCELL_X2 FILLER_17_633 ();
 FILLCELL_X1 FILLER_17_638 ();
 FILLCELL_X2 FILLER_17_660 ();
 FILLCELL_X1 FILLER_17_662 ();
 FILLCELL_X4 FILLER_17_677 ();
 FILLCELL_X1 FILLER_17_681 ();
 FILLCELL_X32 FILLER_17_699 ();
 FILLCELL_X4 FILLER_17_731 ();
 FILLCELL_X1 FILLER_17_735 ();
 FILLCELL_X1 FILLER_17_747 ();
 FILLCELL_X4 FILLER_17_772 ();
 FILLCELL_X2 FILLER_17_776 ();
 FILLCELL_X1 FILLER_17_778 ();
 FILLCELL_X2 FILLER_17_800 ();
 FILLCELL_X1 FILLER_17_802 ();
 FILLCELL_X8 FILLER_17_834 ();
 FILLCELL_X4 FILLER_17_842 ();
 FILLCELL_X2 FILLER_17_846 ();
 FILLCELL_X4 FILLER_17_859 ();
 FILLCELL_X1 FILLER_17_874 ();
 FILLCELL_X8 FILLER_17_901 ();
 FILLCELL_X1 FILLER_17_909 ();
 FILLCELL_X4 FILLER_17_915 ();
 FILLCELL_X2 FILLER_17_928 ();
 FILLCELL_X1 FILLER_17_930 ();
 FILLCELL_X8 FILLER_17_941 ();
 FILLCELL_X2 FILLER_17_952 ();
 FILLCELL_X1 FILLER_17_954 ();
 FILLCELL_X32 FILLER_17_959 ();
 FILLCELL_X8 FILLER_17_991 ();
 FILLCELL_X8 FILLER_17_1021 ();
 FILLCELL_X4 FILLER_17_1041 ();
 FILLCELL_X1 FILLER_17_1045 ();
 FILLCELL_X4 FILLER_17_1049 ();
 FILLCELL_X2 FILLER_17_1080 ();
 FILLCELL_X1 FILLER_17_1082 ();
 FILLCELL_X2 FILLER_17_1098 ();
 FILLCELL_X1 FILLER_17_1100 ();
 FILLCELL_X4 FILLER_17_1104 ();
 FILLCELL_X2 FILLER_17_1172 ();
 FILLCELL_X1 FILLER_17_1174 ();
 FILLCELL_X2 FILLER_17_1198 ();
 FILLCELL_X1 FILLER_17_1209 ();
 FILLCELL_X2 FILLER_17_1226 ();
 FILLCELL_X2 FILLER_17_1232 ();
 FILLCELL_X4 FILLER_17_1247 ();
 FILLCELL_X4 FILLER_17_1258 ();
 FILLCELL_X1 FILLER_17_1262 ();
 FILLCELL_X16 FILLER_17_1264 ();
 FILLCELL_X8 FILLER_17_1280 ();
 FILLCELL_X4 FILLER_17_1288 ();
 FILLCELL_X2 FILLER_17_1292 ();
 FILLCELL_X1 FILLER_17_1294 ();
 FILLCELL_X1 FILLER_17_1302 ();
 FILLCELL_X2 FILLER_17_1307 ();
 FILLCELL_X1 FILLER_17_1316 ();
 FILLCELL_X8 FILLER_17_1348 ();
 FILLCELL_X1 FILLER_17_1356 ();
 FILLCELL_X4 FILLER_17_1372 ();
 FILLCELL_X1 FILLER_17_1376 ();
 FILLCELL_X8 FILLER_17_1381 ();
 FILLCELL_X1 FILLER_17_1395 ();
 FILLCELL_X4 FILLER_17_1401 ();
 FILLCELL_X1 FILLER_17_1405 ();
 FILLCELL_X8 FILLER_17_1416 ();
 FILLCELL_X1 FILLER_17_1424 ();
 FILLCELL_X4 FILLER_17_1437 ();
 FILLCELL_X8 FILLER_17_1448 ();
 FILLCELL_X32 FILLER_17_1460 ();
 FILLCELL_X32 FILLER_17_1492 ();
 FILLCELL_X32 FILLER_17_1524 ();
 FILLCELL_X32 FILLER_17_1556 ();
 FILLCELL_X32 FILLER_17_1588 ();
 FILLCELL_X16 FILLER_17_1620 ();
 FILLCELL_X8 FILLER_17_1636 ();
 FILLCELL_X4 FILLER_17_1644 ();
 FILLCELL_X2 FILLER_17_1648 ();
 FILLCELL_X1 FILLER_17_1650 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X8 FILLER_18_161 ();
 FILLCELL_X2 FILLER_18_169 ();
 FILLCELL_X1 FILLER_18_171 ();
 FILLCELL_X1 FILLER_18_179 ();
 FILLCELL_X2 FILLER_18_184 ();
 FILLCELL_X2 FILLER_18_193 ();
 FILLCELL_X1 FILLER_18_195 ();
 FILLCELL_X8 FILLER_18_209 ();
 FILLCELL_X2 FILLER_18_217 ();
 FILLCELL_X1 FILLER_18_219 ();
 FILLCELL_X8 FILLER_18_224 ();
 FILLCELL_X2 FILLER_18_232 ();
 FILLCELL_X16 FILLER_18_273 ();
 FILLCELL_X8 FILLER_18_289 ();
 FILLCELL_X1 FILLER_18_297 ();
 FILLCELL_X8 FILLER_18_305 ();
 FILLCELL_X2 FILLER_18_313 ();
 FILLCELL_X4 FILLER_18_340 ();
 FILLCELL_X2 FILLER_18_344 ();
 FILLCELL_X1 FILLER_18_346 ();
 FILLCELL_X8 FILLER_18_354 ();
 FILLCELL_X4 FILLER_18_362 ();
 FILLCELL_X1 FILLER_18_366 ();
 FILLCELL_X2 FILLER_18_378 ();
 FILLCELL_X16 FILLER_18_391 ();
 FILLCELL_X4 FILLER_18_407 ();
 FILLCELL_X2 FILLER_18_411 ();
 FILLCELL_X4 FILLER_18_420 ();
 FILLCELL_X2 FILLER_18_424 ();
 FILLCELL_X16 FILLER_18_442 ();
 FILLCELL_X8 FILLER_18_458 ();
 FILLCELL_X1 FILLER_18_466 ();
 FILLCELL_X2 FILLER_18_471 ();
 FILLCELL_X1 FILLER_18_493 ();
 FILLCELL_X2 FILLER_18_499 ();
 FILLCELL_X1 FILLER_18_504 ();
 FILLCELL_X2 FILLER_18_512 ();
 FILLCELL_X2 FILLER_18_517 ();
 FILLCELL_X1 FILLER_18_519 ();
 FILLCELL_X4 FILLER_18_538 ();
 FILLCELL_X2 FILLER_18_546 ();
 FILLCELL_X1 FILLER_18_548 ();
 FILLCELL_X1 FILLER_18_561 ();
 FILLCELL_X16 FILLER_18_589 ();
 FILLCELL_X4 FILLER_18_605 ();
 FILLCELL_X1 FILLER_18_630 ();
 FILLCELL_X1 FILLER_18_632 ();
 FILLCELL_X8 FILLER_18_637 ();
 FILLCELL_X2 FILLER_18_652 ();
 FILLCELL_X16 FILLER_18_676 ();
 FILLCELL_X2 FILLER_18_692 ();
 FILLCELL_X8 FILLER_18_711 ();
 FILLCELL_X2 FILLER_18_719 ();
 FILLCELL_X1 FILLER_18_721 ();
 FILLCELL_X2 FILLER_18_741 ();
 FILLCELL_X1 FILLER_18_743 ();
 FILLCELL_X2 FILLER_18_747 ();
 FILLCELL_X4 FILLER_18_767 ();
 FILLCELL_X1 FILLER_18_771 ();
 FILLCELL_X4 FILLER_18_775 ();
 FILLCELL_X2 FILLER_18_779 ();
 FILLCELL_X4 FILLER_18_799 ();
 FILLCELL_X1 FILLER_18_803 ();
 FILLCELL_X4 FILLER_18_832 ();
 FILLCELL_X1 FILLER_18_836 ();
 FILLCELL_X8 FILLER_18_840 ();
 FILLCELL_X2 FILLER_18_848 ();
 FILLCELL_X2 FILLER_18_853 ();
 FILLCELL_X1 FILLER_18_865 ();
 FILLCELL_X8 FILLER_18_870 ();
 FILLCELL_X4 FILLER_18_878 ();
 FILLCELL_X2 FILLER_18_886 ();
 FILLCELL_X1 FILLER_18_914 ();
 FILLCELL_X4 FILLER_18_926 ();
 FILLCELL_X2 FILLER_18_939 ();
 FILLCELL_X1 FILLER_18_941 ();
 FILLCELL_X8 FILLER_18_958 ();
 FILLCELL_X2 FILLER_18_966 ();
 FILLCELL_X16 FILLER_18_985 ();
 FILLCELL_X1 FILLER_18_1001 ();
 FILLCELL_X8 FILLER_18_1011 ();
 FILLCELL_X2 FILLER_18_1019 ();
 FILLCELL_X1 FILLER_18_1021 ();
 FILLCELL_X1 FILLER_18_1031 ();
 FILLCELL_X4 FILLER_18_1039 ();
 FILLCELL_X1 FILLER_18_1043 ();
 FILLCELL_X2 FILLER_18_1055 ();
 FILLCELL_X2 FILLER_18_1061 ();
 FILLCELL_X1 FILLER_18_1063 ();
 FILLCELL_X1 FILLER_18_1075 ();
 FILLCELL_X4 FILLER_18_1085 ();
 FILLCELL_X2 FILLER_18_1089 ();
 FILLCELL_X1 FILLER_18_1091 ();
 FILLCELL_X8 FILLER_18_1096 ();
 FILLCELL_X1 FILLER_18_1104 ();
 FILLCELL_X2 FILLER_18_1117 ();
 FILLCELL_X4 FILLER_18_1146 ();
 FILLCELL_X2 FILLER_18_1150 ();
 FILLCELL_X1 FILLER_18_1152 ();
 FILLCELL_X1 FILLER_18_1156 ();
 FILLCELL_X1 FILLER_18_1161 ();
 FILLCELL_X1 FILLER_18_1166 ();
 FILLCELL_X2 FILLER_18_1171 ();
 FILLCELL_X4 FILLER_18_1176 ();
 FILLCELL_X2 FILLER_18_1187 ();
 FILLCELL_X4 FILLER_18_1218 ();
 FILLCELL_X2 FILLER_18_1222 ();
 FILLCELL_X1 FILLER_18_1224 ();
 FILLCELL_X1 FILLER_18_1228 ();
 FILLCELL_X1 FILLER_18_1232 ();
 FILLCELL_X1 FILLER_18_1237 ();
 FILLCELL_X1 FILLER_18_1247 ();
 FILLCELL_X32 FILLER_18_1252 ();
 FILLCELL_X4 FILLER_18_1284 ();
 FILLCELL_X1 FILLER_18_1288 ();
 FILLCELL_X8 FILLER_18_1292 ();
 FILLCELL_X4 FILLER_18_1300 ();
 FILLCELL_X4 FILLER_18_1308 ();
 FILLCELL_X1 FILLER_18_1312 ();
 FILLCELL_X2 FILLER_18_1337 ();
 FILLCELL_X4 FILLER_18_1351 ();
 FILLCELL_X2 FILLER_18_1377 ();
 FILLCELL_X1 FILLER_18_1379 ();
 FILLCELL_X2 FILLER_18_1385 ();
 FILLCELL_X2 FILLER_18_1398 ();
 FILLCELL_X1 FILLER_18_1400 ();
 FILLCELL_X2 FILLER_18_1411 ();
 FILLCELL_X1 FILLER_18_1413 ();
 FILLCELL_X2 FILLER_18_1427 ();
 FILLCELL_X1 FILLER_18_1429 ();
 FILLCELL_X2 FILLER_18_1435 ();
 FILLCELL_X1 FILLER_18_1437 ();
 FILLCELL_X32 FILLER_18_1446 ();
 FILLCELL_X32 FILLER_18_1478 ();
 FILLCELL_X32 FILLER_18_1510 ();
 FILLCELL_X32 FILLER_18_1542 ();
 FILLCELL_X32 FILLER_18_1574 ();
 FILLCELL_X32 FILLER_18_1606 ();
 FILLCELL_X8 FILLER_18_1638 ();
 FILLCELL_X4 FILLER_18_1646 ();
 FILLCELL_X1 FILLER_18_1650 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X8 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_169 ();
 FILLCELL_X2 FILLER_19_173 ();
 FILLCELL_X1 FILLER_19_175 ();
 FILLCELL_X4 FILLER_19_180 ();
 FILLCELL_X1 FILLER_19_184 ();
 FILLCELL_X4 FILLER_19_192 ();
 FILLCELL_X2 FILLER_19_196 ();
 FILLCELL_X4 FILLER_19_222 ();
 FILLCELL_X1 FILLER_19_226 ();
 FILLCELL_X2 FILLER_19_232 ();
 FILLCELL_X2 FILLER_19_266 ();
 FILLCELL_X8 FILLER_19_289 ();
 FILLCELL_X4 FILLER_19_301 ();
 FILLCELL_X2 FILLER_19_312 ();
 FILLCELL_X4 FILLER_19_321 ();
 FILLCELL_X4 FILLER_19_343 ();
 FILLCELL_X2 FILLER_19_351 ();
 FILLCELL_X1 FILLER_19_357 ();
 FILLCELL_X4 FILLER_19_396 ();
 FILLCELL_X2 FILLER_19_400 ();
 FILLCELL_X1 FILLER_19_402 ();
 FILLCELL_X2 FILLER_19_410 ();
 FILLCELL_X32 FILLER_19_430 ();
 FILLCELL_X4 FILLER_19_462 ();
 FILLCELL_X2 FILLER_19_470 ();
 FILLCELL_X2 FILLER_19_489 ();
 FILLCELL_X1 FILLER_19_491 ();
 FILLCELL_X2 FILLER_19_508 ();
 FILLCELL_X2 FILLER_19_513 ();
 FILLCELL_X1 FILLER_19_515 ();
 FILLCELL_X4 FILLER_19_525 ();
 FILLCELL_X2 FILLER_19_529 ();
 FILLCELL_X8 FILLER_19_559 ();
 FILLCELL_X1 FILLER_19_585 ();
 FILLCELL_X4 FILLER_19_590 ();
 FILLCELL_X2 FILLER_19_594 ();
 FILLCELL_X1 FILLER_19_601 ();
 FILLCELL_X4 FILLER_19_634 ();
 FILLCELL_X2 FILLER_19_638 ();
 FILLCELL_X1 FILLER_19_640 ();
 FILLCELL_X1 FILLER_19_645 ();
 FILLCELL_X2 FILLER_19_653 ();
 FILLCELL_X1 FILLER_19_664 ();
 FILLCELL_X32 FILLER_19_677 ();
 FILLCELL_X32 FILLER_19_709 ();
 FILLCELL_X1 FILLER_19_741 ();
 FILLCELL_X4 FILLER_19_756 ();
 FILLCELL_X2 FILLER_19_760 ();
 FILLCELL_X1 FILLER_19_762 ();
 FILLCELL_X4 FILLER_19_786 ();
 FILLCELL_X2 FILLER_19_790 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X4 FILLER_19_845 ();
 FILLCELL_X1 FILLER_19_849 ();
 FILLCELL_X2 FILLER_19_855 ();
 FILLCELL_X8 FILLER_19_903 ();
 FILLCELL_X2 FILLER_19_911 ();
 FILLCELL_X2 FILLER_19_933 ();
 FILLCELL_X1 FILLER_19_935 ();
 FILLCELL_X2 FILLER_19_943 ();
 FILLCELL_X2 FILLER_19_949 ();
 FILLCELL_X1 FILLER_19_951 ();
 FILLCELL_X32 FILLER_19_959 ();
 FILLCELL_X2 FILLER_19_991 ();
 FILLCELL_X1 FILLER_19_993 ();
 FILLCELL_X8 FILLER_19_1072 ();
 FILLCELL_X4 FILLER_19_1080 ();
 FILLCELL_X1 FILLER_19_1084 ();
 FILLCELL_X16 FILLER_19_1092 ();
 FILLCELL_X2 FILLER_19_1108 ();
 FILLCELL_X1 FILLER_19_1110 ();
 FILLCELL_X4 FILLER_19_1125 ();
 FILLCELL_X8 FILLER_19_1147 ();
 FILLCELL_X1 FILLER_19_1188 ();
 FILLCELL_X4 FILLER_19_1205 ();
 FILLCELL_X1 FILLER_19_1209 ();
 FILLCELL_X2 FILLER_19_1214 ();
 FILLCELL_X1 FILLER_19_1216 ();
 FILLCELL_X2 FILLER_19_1243 ();
 FILLCELL_X16 FILLER_19_1264 ();
 FILLCELL_X4 FILLER_19_1280 ();
 FILLCELL_X1 FILLER_19_1284 ();
 FILLCELL_X2 FILLER_19_1298 ();
 FILLCELL_X2 FILLER_19_1312 ();
 FILLCELL_X1 FILLER_19_1323 ();
 FILLCELL_X1 FILLER_19_1333 ();
 FILLCELL_X2 FILLER_19_1338 ();
 FILLCELL_X1 FILLER_19_1340 ();
 FILLCELL_X1 FILLER_19_1345 ();
 FILLCELL_X8 FILLER_19_1350 ();
 FILLCELL_X2 FILLER_19_1370 ();
 FILLCELL_X2 FILLER_19_1378 ();
 FILLCELL_X1 FILLER_19_1380 ();
 FILLCELL_X1 FILLER_19_1391 ();
 FILLCELL_X4 FILLER_19_1412 ();
 FILLCELL_X32 FILLER_19_1434 ();
 FILLCELL_X32 FILLER_19_1466 ();
 FILLCELL_X32 FILLER_19_1498 ();
 FILLCELL_X32 FILLER_19_1530 ();
 FILLCELL_X32 FILLER_19_1562 ();
 FILLCELL_X32 FILLER_19_1594 ();
 FILLCELL_X16 FILLER_19_1626 ();
 FILLCELL_X8 FILLER_19_1642 ();
 FILLCELL_X1 FILLER_19_1650 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_169 ();
 FILLCELL_X2 FILLER_20_173 ();
 FILLCELL_X1 FILLER_20_192 ();
 FILLCELL_X1 FILLER_20_210 ();
 FILLCELL_X1 FILLER_20_237 ();
 FILLCELL_X1 FILLER_20_243 ();
 FILLCELL_X8 FILLER_20_283 ();
 FILLCELL_X4 FILLER_20_291 ();
 FILLCELL_X4 FILLER_20_309 ();
 FILLCELL_X2 FILLER_20_313 ();
 FILLCELL_X8 FILLER_20_335 ();
 FILLCELL_X2 FILLER_20_343 ();
 FILLCELL_X1 FILLER_20_345 ();
 FILLCELL_X1 FILLER_20_353 ();
 FILLCELL_X4 FILLER_20_357 ();
 FILLCELL_X2 FILLER_20_361 ();
 FILLCELL_X1 FILLER_20_372 ();
 FILLCELL_X1 FILLER_20_378 ();
 FILLCELL_X2 FILLER_20_392 ();
 FILLCELL_X8 FILLER_20_398 ();
 FILLCELL_X2 FILLER_20_406 ();
 FILLCELL_X1 FILLER_20_408 ();
 FILLCELL_X2 FILLER_20_426 ();
 FILLCELL_X8 FILLER_20_446 ();
 FILLCELL_X4 FILLER_20_454 ();
 FILLCELL_X2 FILLER_20_458 ();
 FILLCELL_X2 FILLER_20_467 ();
 FILLCELL_X1 FILLER_20_469 ();
 FILLCELL_X2 FILLER_20_477 ();
 FILLCELL_X8 FILLER_20_490 ();
 FILLCELL_X4 FILLER_20_498 ();
 FILLCELL_X1 FILLER_20_502 ();
 FILLCELL_X1 FILLER_20_553 ();
 FILLCELL_X2 FILLER_20_601 ();
 FILLCELL_X1 FILLER_20_603 ();
 FILLCELL_X1 FILLER_20_615 ();
 FILLCELL_X2 FILLER_20_621 ();
 FILLCELL_X1 FILLER_20_623 ();
 FILLCELL_X1 FILLER_20_654 ();
 FILLCELL_X4 FILLER_20_662 ();
 FILLCELL_X2 FILLER_20_666 ();
 FILLCELL_X2 FILLER_20_677 ();
 FILLCELL_X32 FILLER_20_694 ();
 FILLCELL_X8 FILLER_20_726 ();
 FILLCELL_X4 FILLER_20_734 ();
 FILLCELL_X4 FILLER_20_745 ();
 FILLCELL_X2 FILLER_20_756 ();
 FILLCELL_X1 FILLER_20_772 ();
 FILLCELL_X1 FILLER_20_780 ();
 FILLCELL_X2 FILLER_20_790 ();
 FILLCELL_X2 FILLER_20_797 ();
 FILLCELL_X8 FILLER_20_806 ();
 FILLCELL_X1 FILLER_20_814 ();
 FILLCELL_X2 FILLER_20_819 ();
 FILLCELL_X1 FILLER_20_829 ();
 FILLCELL_X4 FILLER_20_837 ();
 FILLCELL_X1 FILLER_20_841 ();
 FILLCELL_X4 FILLER_20_846 ();
 FILLCELL_X2 FILLER_20_850 ();
 FILLCELL_X4 FILLER_20_861 ();
 FILLCELL_X1 FILLER_20_865 ();
 FILLCELL_X4 FILLER_20_873 ();
 FILLCELL_X1 FILLER_20_877 ();
 FILLCELL_X4 FILLER_20_893 ();
 FILLCELL_X4 FILLER_20_902 ();
 FILLCELL_X1 FILLER_20_906 ();
 FILLCELL_X4 FILLER_20_912 ();
 FILLCELL_X4 FILLER_20_928 ();
 FILLCELL_X1 FILLER_20_932 ();
 FILLCELL_X8 FILLER_20_947 ();
 FILLCELL_X4 FILLER_20_955 ();
 FILLCELL_X2 FILLER_20_959 ();
 FILLCELL_X8 FILLER_20_974 ();
 FILLCELL_X2 FILLER_20_982 ();
 FILLCELL_X1 FILLER_20_984 ();
 FILLCELL_X1 FILLER_20_1014 ();
 FILLCELL_X2 FILLER_20_1024 ();
 FILLCELL_X2 FILLER_20_1040 ();
 FILLCELL_X1 FILLER_20_1049 ();
 FILLCELL_X2 FILLER_20_1078 ();
 FILLCELL_X1 FILLER_20_1080 ();
 FILLCELL_X16 FILLER_20_1092 ();
 FILLCELL_X2 FILLER_20_1108 ();
 FILLCELL_X1 FILLER_20_1118 ();
 FILLCELL_X4 FILLER_20_1130 ();
 FILLCELL_X1 FILLER_20_1134 ();
 FILLCELL_X4 FILLER_20_1142 ();
 FILLCELL_X2 FILLER_20_1160 ();
 FILLCELL_X8 FILLER_20_1169 ();
 FILLCELL_X2 FILLER_20_1177 ();
 FILLCELL_X8 FILLER_20_1184 ();
 FILLCELL_X4 FILLER_20_1192 ();
 FILLCELL_X1 FILLER_20_1196 ();
 FILLCELL_X4 FILLER_20_1206 ();
 FILLCELL_X2 FILLER_20_1219 ();
 FILLCELL_X1 FILLER_20_1221 ();
 FILLCELL_X32 FILLER_20_1244 ();
 FILLCELL_X8 FILLER_20_1276 ();
 FILLCELL_X2 FILLER_20_1298 ();
 FILLCELL_X8 FILLER_20_1311 ();
 FILLCELL_X4 FILLER_20_1319 ();
 FILLCELL_X4 FILLER_20_1333 ();
 FILLCELL_X2 FILLER_20_1348 ();
 FILLCELL_X1 FILLER_20_1353 ();
 FILLCELL_X2 FILLER_20_1364 ();
 FILLCELL_X2 FILLER_20_1377 ();
 FILLCELL_X2 FILLER_20_1383 ();
 FILLCELL_X1 FILLER_20_1388 ();
 FILLCELL_X2 FILLER_20_1405 ();
 FILLCELL_X1 FILLER_20_1407 ();
 FILLCELL_X16 FILLER_20_1412 ();
 FILLCELL_X8 FILLER_20_1428 ();
 FILLCELL_X4 FILLER_20_1436 ();
 FILLCELL_X2 FILLER_20_1440 ();
 FILLCELL_X4 FILLER_20_1446 ();
 FILLCELL_X32 FILLER_20_1457 ();
 FILLCELL_X32 FILLER_20_1489 ();
 FILLCELL_X32 FILLER_20_1521 ();
 FILLCELL_X32 FILLER_20_1553 ();
 FILLCELL_X32 FILLER_20_1585 ();
 FILLCELL_X32 FILLER_20_1617 ();
 FILLCELL_X2 FILLER_20_1649 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X8 FILLER_21_161 ();
 FILLCELL_X2 FILLER_21_169 ();
 FILLCELL_X1 FILLER_21_171 ();
 FILLCELL_X2 FILLER_21_175 ();
 FILLCELL_X2 FILLER_21_190 ();
 FILLCELL_X1 FILLER_21_192 ();
 FILLCELL_X1 FILLER_21_207 ();
 FILLCELL_X8 FILLER_21_232 ();
 FILLCELL_X4 FILLER_21_240 ();
 FILLCELL_X2 FILLER_21_244 ();
 FILLCELL_X1 FILLER_21_246 ();
 FILLCELL_X16 FILLER_21_251 ();
 FILLCELL_X8 FILLER_21_267 ();
 FILLCELL_X8 FILLER_21_278 ();
 FILLCELL_X4 FILLER_21_299 ();
 FILLCELL_X16 FILLER_21_307 ();
 FILLCELL_X1 FILLER_21_323 ();
 FILLCELL_X8 FILLER_21_327 ();
 FILLCELL_X2 FILLER_21_335 ();
 FILLCELL_X2 FILLER_21_341 ();
 FILLCELL_X2 FILLER_21_352 ();
 FILLCELL_X8 FILLER_21_363 ();
 FILLCELL_X4 FILLER_21_371 ();
 FILLCELL_X2 FILLER_21_375 ();
 FILLCELL_X1 FILLER_21_377 ();
 FILLCELL_X8 FILLER_21_401 ();
 FILLCELL_X16 FILLER_21_444 ();
 FILLCELL_X4 FILLER_21_477 ();
 FILLCELL_X1 FILLER_21_485 ();
 FILLCELL_X8 FILLER_21_489 ();
 FILLCELL_X2 FILLER_21_497 ();
 FILLCELL_X16 FILLER_21_535 ();
 FILLCELL_X8 FILLER_21_551 ();
 FILLCELL_X2 FILLER_21_559 ();
 FILLCELL_X8 FILLER_21_570 ();
 FILLCELL_X1 FILLER_21_578 ();
 FILLCELL_X2 FILLER_21_584 ();
 FILLCELL_X2 FILLER_21_593 ();
 FILLCELL_X1 FILLER_21_595 ();
 FILLCELL_X1 FILLER_21_621 ();
 FILLCELL_X8 FILLER_21_626 ();
 FILLCELL_X1 FILLER_21_634 ();
 FILLCELL_X1 FILLER_21_648 ();
 FILLCELL_X1 FILLER_21_654 ();
 FILLCELL_X8 FILLER_21_680 ();
 FILLCELL_X2 FILLER_21_688 ();
 FILLCELL_X1 FILLER_21_690 ();
 FILLCELL_X32 FILLER_21_708 ();
 FILLCELL_X2 FILLER_21_747 ();
 FILLCELL_X1 FILLER_21_754 ();
 FILLCELL_X2 FILLER_21_760 ();
 FILLCELL_X4 FILLER_21_767 ();
 FILLCELL_X1 FILLER_21_771 ();
 FILLCELL_X4 FILLER_21_784 ();
 FILLCELL_X1 FILLER_21_788 ();
 FILLCELL_X2 FILLER_21_797 ();
 FILLCELL_X1 FILLER_21_799 ();
 FILLCELL_X4 FILLER_21_809 ();
 FILLCELL_X1 FILLER_21_813 ();
 FILLCELL_X4 FILLER_21_817 ();
 FILLCELL_X1 FILLER_21_821 ();
 FILLCELL_X8 FILLER_21_839 ();
 FILLCELL_X2 FILLER_21_847 ();
 FILLCELL_X2 FILLER_21_865 ();
 FILLCELL_X4 FILLER_21_872 ();
 FILLCELL_X2 FILLER_21_876 ();
 FILLCELL_X2 FILLER_21_906 ();
 FILLCELL_X1 FILLER_21_944 ();
 FILLCELL_X32 FILLER_21_950 ();
 FILLCELL_X16 FILLER_21_982 ();
 FILLCELL_X2 FILLER_21_998 ();
 FILLCELL_X1 FILLER_21_1000 ();
 FILLCELL_X16 FILLER_21_1012 ();
 FILLCELL_X4 FILLER_21_1028 ();
 FILLCELL_X2 FILLER_21_1032 ();
 FILLCELL_X2 FILLER_21_1052 ();
 FILLCELL_X4 FILLER_21_1063 ();
 FILLCELL_X4 FILLER_21_1088 ();
 FILLCELL_X4 FILLER_21_1106 ();
 FILLCELL_X2 FILLER_21_1121 ();
 FILLCELL_X2 FILLER_21_1127 ();
 FILLCELL_X1 FILLER_21_1143 ();
 FILLCELL_X1 FILLER_21_1155 ();
 FILLCELL_X1 FILLER_21_1160 ();
 FILLCELL_X8 FILLER_21_1182 ();
 FILLCELL_X1 FILLER_21_1190 ();
 FILLCELL_X8 FILLER_21_1196 ();
 FILLCELL_X2 FILLER_21_1204 ();
 FILLCELL_X1 FILLER_21_1213 ();
 FILLCELL_X2 FILLER_21_1231 ();
 FILLCELL_X1 FILLER_21_1240 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X2 FILLER_21_1296 ();
 FILLCELL_X2 FILLER_21_1307 ();
 FILLCELL_X1 FILLER_21_1316 ();
 FILLCELL_X4 FILLER_21_1324 ();
 FILLCELL_X2 FILLER_21_1328 ();
 FILLCELL_X1 FILLER_21_1330 ();
 FILLCELL_X4 FILLER_21_1336 ();
 FILLCELL_X1 FILLER_21_1340 ();
 FILLCELL_X1 FILLER_21_1354 ();
 FILLCELL_X8 FILLER_21_1369 ();
 FILLCELL_X1 FILLER_21_1381 ();
 FILLCELL_X2 FILLER_21_1386 ();
 FILLCELL_X1 FILLER_21_1392 ();
 FILLCELL_X8 FILLER_21_1396 ();
 FILLCELL_X2 FILLER_21_1412 ();
 FILLCELL_X1 FILLER_21_1422 ();
 FILLCELL_X1 FILLER_21_1427 ();
 FILLCELL_X2 FILLER_21_1445 ();
 FILLCELL_X1 FILLER_21_1447 ();
 FILLCELL_X32 FILLER_21_1455 ();
 FILLCELL_X32 FILLER_21_1487 ();
 FILLCELL_X32 FILLER_21_1519 ();
 FILLCELL_X32 FILLER_21_1551 ();
 FILLCELL_X32 FILLER_21_1583 ();
 FILLCELL_X32 FILLER_21_1615 ();
 FILLCELL_X4 FILLER_21_1647 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X16 FILLER_22_161 ();
 FILLCELL_X2 FILLER_22_189 ();
 FILLCELL_X1 FILLER_22_198 ();
 FILLCELL_X1 FILLER_22_203 ();
 FILLCELL_X2 FILLER_22_209 ();
 FILLCELL_X1 FILLER_22_211 ();
 FILLCELL_X4 FILLER_22_221 ();
 FILLCELL_X1 FILLER_22_225 ();
 FILLCELL_X2 FILLER_22_233 ();
 FILLCELL_X1 FILLER_22_235 ();
 FILLCELL_X2 FILLER_22_240 ();
 FILLCELL_X4 FILLER_22_249 ();
 FILLCELL_X8 FILLER_22_258 ();
 FILLCELL_X4 FILLER_22_300 ();
 FILLCELL_X2 FILLER_22_304 ();
 FILLCELL_X1 FILLER_22_312 ();
 FILLCELL_X4 FILLER_22_324 ();
 FILLCELL_X2 FILLER_22_328 ();
 FILLCELL_X2 FILLER_22_334 ();
 FILLCELL_X1 FILLER_22_336 ();
 FILLCELL_X4 FILLER_22_344 ();
 FILLCELL_X1 FILLER_22_357 ();
 FILLCELL_X2 FILLER_22_365 ();
 FILLCELL_X1 FILLER_22_379 ();
 FILLCELL_X1 FILLER_22_387 ();
 FILLCELL_X16 FILLER_22_392 ();
 FILLCELL_X2 FILLER_22_408 ();
 FILLCELL_X2 FILLER_22_419 ();
 FILLCELL_X1 FILLER_22_421 ();
 FILLCELL_X16 FILLER_22_448 ();
 FILLCELL_X2 FILLER_22_464 ();
 FILLCELL_X1 FILLER_22_477 ();
 FILLCELL_X1 FILLER_22_491 ();
 FILLCELL_X2 FILLER_22_499 ();
 FILLCELL_X2 FILLER_22_519 ();
 FILLCELL_X2 FILLER_22_535 ();
 FILLCELL_X1 FILLER_22_537 ();
 FILLCELL_X8 FILLER_22_558 ();
 FILLCELL_X2 FILLER_22_566 ();
 FILLCELL_X1 FILLER_22_568 ();
 FILLCELL_X4 FILLER_22_573 ();
 FILLCELL_X4 FILLER_22_590 ();
 FILLCELL_X1 FILLER_22_594 ();
 FILLCELL_X4 FILLER_22_613 ();
 FILLCELL_X4 FILLER_22_627 ();
 FILLCELL_X2 FILLER_22_659 ();
 FILLCELL_X2 FILLER_22_670 ();
 FILLCELL_X4 FILLER_22_681 ();
 FILLCELL_X16 FILLER_22_714 ();
 FILLCELL_X4 FILLER_22_730 ();
 FILLCELL_X2 FILLER_22_734 ();
 FILLCELL_X1 FILLER_22_736 ();
 FILLCELL_X1 FILLER_22_751 ();
 FILLCELL_X2 FILLER_22_756 ();
 FILLCELL_X8 FILLER_22_781 ();
 FILLCELL_X4 FILLER_22_789 ();
 FILLCELL_X2 FILLER_22_800 ();
 FILLCELL_X1 FILLER_22_802 ();
 FILLCELL_X1 FILLER_22_812 ();
 FILLCELL_X4 FILLER_22_820 ();
 FILLCELL_X2 FILLER_22_824 ();
 FILLCELL_X1 FILLER_22_826 ();
 FILLCELL_X1 FILLER_22_831 ();
 FILLCELL_X16 FILLER_22_859 ();
 FILLCELL_X2 FILLER_22_875 ();
 FILLCELL_X1 FILLER_22_877 ();
 FILLCELL_X2 FILLER_22_908 ();
 FILLCELL_X1 FILLER_22_941 ();
 FILLCELL_X32 FILLER_22_953 ();
 FILLCELL_X1 FILLER_22_1020 ();
 FILLCELL_X1 FILLER_22_1090 ();
 FILLCELL_X1 FILLER_22_1100 ();
 FILLCELL_X1 FILLER_22_1108 ();
 FILLCELL_X2 FILLER_22_1120 ();
 FILLCELL_X1 FILLER_22_1129 ();
 FILLCELL_X1 FILLER_22_1135 ();
 FILLCELL_X1 FILLER_22_1147 ();
 FILLCELL_X1 FILLER_22_1155 ();
 FILLCELL_X1 FILLER_22_1160 ();
 FILLCELL_X8 FILLER_22_1165 ();
 FILLCELL_X2 FILLER_22_1181 ();
 FILLCELL_X4 FILLER_22_1204 ();
 FILLCELL_X2 FILLER_22_1208 ();
 FILLCELL_X1 FILLER_22_1234 ();
 FILLCELL_X4 FILLER_22_1244 ();
 FILLCELL_X2 FILLER_22_1248 ();
 FILLCELL_X16 FILLER_22_1257 ();
 FILLCELL_X8 FILLER_22_1273 ();
 FILLCELL_X1 FILLER_22_1281 ();
 FILLCELL_X1 FILLER_22_1289 ();
 FILLCELL_X1 FILLER_22_1299 ();
 FILLCELL_X1 FILLER_22_1304 ();
 FILLCELL_X1 FILLER_22_1316 ();
 FILLCELL_X2 FILLER_22_1321 ();
 FILLCELL_X4 FILLER_22_1327 ();
 FILLCELL_X2 FILLER_22_1336 ();
 FILLCELL_X2 FILLER_22_1341 ();
 FILLCELL_X1 FILLER_22_1343 ();
 FILLCELL_X2 FILLER_22_1347 ();
 FILLCELL_X2 FILLER_22_1366 ();
 FILLCELL_X4 FILLER_22_1385 ();
 FILLCELL_X2 FILLER_22_1389 ();
 FILLCELL_X4 FILLER_22_1395 ();
 FILLCELL_X2 FILLER_22_1402 ();
 FILLCELL_X1 FILLER_22_1404 ();
 FILLCELL_X4 FILLER_22_1423 ();
 FILLCELL_X1 FILLER_22_1434 ();
 FILLCELL_X2 FILLER_22_1439 ();
 FILLCELL_X8 FILLER_22_1449 ();
 FILLCELL_X1 FILLER_22_1457 ();
 FILLCELL_X32 FILLER_22_1465 ();
 FILLCELL_X32 FILLER_22_1497 ();
 FILLCELL_X32 FILLER_22_1529 ();
 FILLCELL_X32 FILLER_22_1561 ();
 FILLCELL_X32 FILLER_22_1593 ();
 FILLCELL_X16 FILLER_22_1625 ();
 FILLCELL_X8 FILLER_22_1641 ();
 FILLCELL_X2 FILLER_22_1649 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X8 FILLER_23_161 ();
 FILLCELL_X4 FILLER_23_169 ();
 FILLCELL_X4 FILLER_23_205 ();
 FILLCELL_X2 FILLER_23_209 ();
 FILLCELL_X1 FILLER_23_211 ();
 FILLCELL_X8 FILLER_23_225 ();
 FILLCELL_X1 FILLER_23_233 ();
 FILLCELL_X1 FILLER_23_238 ();
 FILLCELL_X2 FILLER_23_242 ();
 FILLCELL_X1 FILLER_23_244 ();
 FILLCELL_X2 FILLER_23_248 ();
 FILLCELL_X2 FILLER_23_254 ();
 FILLCELL_X4 FILLER_23_263 ();
 FILLCELL_X1 FILLER_23_267 ();
 FILLCELL_X2 FILLER_23_302 ();
 FILLCELL_X2 FILLER_23_311 ();
 FILLCELL_X1 FILLER_23_313 ();
 FILLCELL_X2 FILLER_23_321 ();
 FILLCELL_X4 FILLER_23_341 ();
 FILLCELL_X2 FILLER_23_345 ();
 FILLCELL_X1 FILLER_23_347 ();
 FILLCELL_X1 FILLER_23_355 ();
 FILLCELL_X4 FILLER_23_368 ();
 FILLCELL_X1 FILLER_23_385 ();
 FILLCELL_X1 FILLER_23_393 ();
 FILLCELL_X1 FILLER_23_411 ();
 FILLCELL_X1 FILLER_23_425 ();
 FILLCELL_X16 FILLER_23_437 ();
 FILLCELL_X8 FILLER_23_453 ();
 FILLCELL_X4 FILLER_23_461 ();
 FILLCELL_X2 FILLER_23_465 ();
 FILLCELL_X1 FILLER_23_467 ();
 FILLCELL_X4 FILLER_23_484 ();
 FILLCELL_X2 FILLER_23_488 ();
 FILLCELL_X4 FILLER_23_497 ();
 FILLCELL_X2 FILLER_23_508 ();
 FILLCELL_X1 FILLER_23_510 ();
 FILLCELL_X2 FILLER_23_514 ();
 FILLCELL_X4 FILLER_23_525 ();
 FILLCELL_X2 FILLER_23_529 ();
 FILLCELL_X1 FILLER_23_531 ();
 FILLCELL_X8 FILLER_23_536 ();
 FILLCELL_X4 FILLER_23_544 ();
 FILLCELL_X1 FILLER_23_552 ();
 FILLCELL_X16 FILLER_23_557 ();
 FILLCELL_X4 FILLER_23_593 ();
 FILLCELL_X1 FILLER_23_611 ();
 FILLCELL_X4 FILLER_23_621 ();
 FILLCELL_X4 FILLER_23_629 ();
 FILLCELL_X1 FILLER_23_633 ();
 FILLCELL_X1 FILLER_23_645 ();
 FILLCELL_X2 FILLER_23_653 ();
 FILLCELL_X2 FILLER_23_662 ();
 FILLCELL_X2 FILLER_23_678 ();
 FILLCELL_X2 FILLER_23_683 ();
 FILLCELL_X1 FILLER_23_685 ();
 FILLCELL_X32 FILLER_23_703 ();
 FILLCELL_X2 FILLER_23_735 ();
 FILLCELL_X1 FILLER_23_737 ();
 FILLCELL_X1 FILLER_23_762 ();
 FILLCELL_X1 FILLER_23_770 ();
 FILLCELL_X1 FILLER_23_780 ();
 FILLCELL_X1 FILLER_23_788 ();
 FILLCELL_X1 FILLER_23_796 ();
 FILLCELL_X1 FILLER_23_813 ();
 FILLCELL_X8 FILLER_23_818 ();
 FILLCELL_X2 FILLER_23_826 ();
 FILLCELL_X1 FILLER_23_828 ();
 FILLCELL_X8 FILLER_23_842 ();
 FILLCELL_X2 FILLER_23_850 ();
 FILLCELL_X1 FILLER_23_861 ();
 FILLCELL_X1 FILLER_23_865 ();
 FILLCELL_X2 FILLER_23_887 ();
 FILLCELL_X1 FILLER_23_889 ();
 FILLCELL_X4 FILLER_23_905 ();
 FILLCELL_X16 FILLER_23_927 ();
 FILLCELL_X8 FILLER_23_943 ();
 FILLCELL_X2 FILLER_23_951 ();
 FILLCELL_X1 FILLER_23_953 ();
 FILLCELL_X8 FILLER_23_970 ();
 FILLCELL_X2 FILLER_23_978 ();
 FILLCELL_X2 FILLER_23_996 ();
 FILLCELL_X2 FILLER_23_1007 ();
 FILLCELL_X1 FILLER_23_1009 ();
 FILLCELL_X2 FILLER_23_1020 ();
 FILLCELL_X4 FILLER_23_1048 ();
 FILLCELL_X2 FILLER_23_1052 ();
 FILLCELL_X1 FILLER_23_1054 ();
 FILLCELL_X1 FILLER_23_1073 ();
 FILLCELL_X1 FILLER_23_1115 ();
 FILLCELL_X2 FILLER_23_1151 ();
 FILLCELL_X1 FILLER_23_1153 ();
 FILLCELL_X4 FILLER_23_1165 ();
 FILLCELL_X2 FILLER_23_1173 ();
 FILLCELL_X16 FILLER_23_1185 ();
 FILLCELL_X2 FILLER_23_1201 ();
 FILLCELL_X1 FILLER_23_1203 ();
 FILLCELL_X1 FILLER_23_1208 ();
 FILLCELL_X8 FILLER_23_1213 ();
 FILLCELL_X4 FILLER_23_1221 ();
 FILLCELL_X2 FILLER_23_1240 ();
 FILLCELL_X1 FILLER_23_1242 ();
 FILLCELL_X8 FILLER_23_1250 ();
 FILLCELL_X4 FILLER_23_1258 ();
 FILLCELL_X1 FILLER_23_1262 ();
 FILLCELL_X8 FILLER_23_1264 ();
 FILLCELL_X4 FILLER_23_1272 ();
 FILLCELL_X2 FILLER_23_1285 ();
 FILLCELL_X8 FILLER_23_1296 ();
 FILLCELL_X4 FILLER_23_1308 ();
 FILLCELL_X2 FILLER_23_1317 ();
 FILLCELL_X4 FILLER_23_1324 ();
 FILLCELL_X2 FILLER_23_1331 ();
 FILLCELL_X8 FILLER_23_1346 ();
 FILLCELL_X4 FILLER_23_1354 ();
 FILLCELL_X2 FILLER_23_1358 ();
 FILLCELL_X1 FILLER_23_1360 ();
 FILLCELL_X1 FILLER_23_1373 ();
 FILLCELL_X4 FILLER_23_1378 ();
 FILLCELL_X1 FILLER_23_1382 ();
 FILLCELL_X2 FILLER_23_1407 ();
 FILLCELL_X1 FILLER_23_1419 ();
 FILLCELL_X1 FILLER_23_1439 ();
 FILLCELL_X32 FILLER_23_1451 ();
 FILLCELL_X32 FILLER_23_1483 ();
 FILLCELL_X32 FILLER_23_1515 ();
 FILLCELL_X32 FILLER_23_1547 ();
 FILLCELL_X32 FILLER_23_1579 ();
 FILLCELL_X32 FILLER_23_1611 ();
 FILLCELL_X8 FILLER_23_1643 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X8 FILLER_24_161 ();
 FILLCELL_X2 FILLER_24_169 ();
 FILLCELL_X1 FILLER_24_171 ();
 FILLCELL_X1 FILLER_24_179 ();
 FILLCELL_X1 FILLER_24_189 ();
 FILLCELL_X2 FILLER_24_194 ();
 FILLCELL_X4 FILLER_24_216 ();
 FILLCELL_X2 FILLER_24_220 ();
 FILLCELL_X4 FILLER_24_227 ();
 FILLCELL_X2 FILLER_24_231 ();
 FILLCELL_X2 FILLER_24_243 ();
 FILLCELL_X16 FILLER_24_265 ();
 FILLCELL_X2 FILLER_24_281 ();
 FILLCELL_X2 FILLER_24_287 ();
 FILLCELL_X4 FILLER_24_299 ();
 FILLCELL_X1 FILLER_24_303 ();
 FILLCELL_X16 FILLER_24_338 ();
 FILLCELL_X4 FILLER_24_354 ();
 FILLCELL_X2 FILLER_24_358 ();
 FILLCELL_X4 FILLER_24_378 ();
 FILLCELL_X4 FILLER_24_391 ();
 FILLCELL_X2 FILLER_24_395 ();
 FILLCELL_X1 FILLER_24_397 ();
 FILLCELL_X4 FILLER_24_429 ();
 FILLCELL_X2 FILLER_24_433 ();
 FILLCELL_X1 FILLER_24_435 ();
 FILLCELL_X16 FILLER_24_454 ();
 FILLCELL_X8 FILLER_24_470 ();
 FILLCELL_X1 FILLER_24_478 ();
 FILLCELL_X1 FILLER_24_486 ();
 FILLCELL_X4 FILLER_24_494 ();
 FILLCELL_X2 FILLER_24_498 ();
 FILLCELL_X4 FILLER_24_504 ();
 FILLCELL_X1 FILLER_24_521 ();
 FILLCELL_X1 FILLER_24_549 ();
 FILLCELL_X8 FILLER_24_566 ();
 FILLCELL_X4 FILLER_24_574 ();
 FILLCELL_X1 FILLER_24_578 ();
 FILLCELL_X16 FILLER_24_597 ();
 FILLCELL_X2 FILLER_24_613 ();
 FILLCELL_X1 FILLER_24_630 ();
 FILLCELL_X1 FILLER_24_644 ();
 FILLCELL_X2 FILLER_24_650 ();
 FILLCELL_X1 FILLER_24_673 ();
 FILLCELL_X4 FILLER_24_683 ();
 FILLCELL_X8 FILLER_24_694 ();
 FILLCELL_X2 FILLER_24_702 ();
 FILLCELL_X1 FILLER_24_704 ();
 FILLCELL_X2 FILLER_24_723 ();
 FILLCELL_X1 FILLER_24_725 ();
 FILLCELL_X2 FILLER_24_740 ();
 FILLCELL_X1 FILLER_24_742 ();
 FILLCELL_X4 FILLER_24_750 ();
 FILLCELL_X2 FILLER_24_754 ();
 FILLCELL_X4 FILLER_24_774 ();
 FILLCELL_X4 FILLER_24_787 ();
 FILLCELL_X2 FILLER_24_791 ();
 FILLCELL_X2 FILLER_24_820 ();
 FILLCELL_X1 FILLER_24_822 ();
 FILLCELL_X1 FILLER_24_830 ();
 FILLCELL_X2 FILLER_24_834 ();
 FILLCELL_X1 FILLER_24_842 ();
 FILLCELL_X4 FILLER_24_850 ();
 FILLCELL_X1 FILLER_24_854 ();
 FILLCELL_X2 FILLER_24_858 ();
 FILLCELL_X1 FILLER_24_878 ();
 FILLCELL_X8 FILLER_24_896 ();
 FILLCELL_X8 FILLER_24_917 ();
 FILLCELL_X4 FILLER_24_925 ();
 FILLCELL_X1 FILLER_24_929 ();
 FILLCELL_X2 FILLER_24_937 ();
 FILLCELL_X16 FILLER_24_963 ();
 FILLCELL_X4 FILLER_24_979 ();
 FILLCELL_X1 FILLER_24_983 ();
 FILLCELL_X4 FILLER_24_1013 ();
 FILLCELL_X4 FILLER_24_1024 ();
 FILLCELL_X2 FILLER_24_1028 ();
 FILLCELL_X1 FILLER_24_1030 ();
 FILLCELL_X8 FILLER_24_1049 ();
 FILLCELL_X1 FILLER_24_1057 ();
 FILLCELL_X4 FILLER_24_1086 ();
 FILLCELL_X1 FILLER_24_1104 ();
 FILLCELL_X4 FILLER_24_1109 ();
 FILLCELL_X2 FILLER_24_1113 ();
 FILLCELL_X4 FILLER_24_1124 ();
 FILLCELL_X2 FILLER_24_1128 ();
 FILLCELL_X4 FILLER_24_1153 ();
 FILLCELL_X2 FILLER_24_1157 ();
 FILLCELL_X2 FILLER_24_1168 ();
 FILLCELL_X8 FILLER_24_1177 ();
 FILLCELL_X1 FILLER_24_1185 ();
 FILLCELL_X8 FILLER_24_1190 ();
 FILLCELL_X2 FILLER_24_1214 ();
 FILLCELL_X1 FILLER_24_1216 ();
 FILLCELL_X4 FILLER_24_1237 ();
 FILLCELL_X2 FILLER_24_1241 ();
 FILLCELL_X1 FILLER_24_1243 ();
 FILLCELL_X8 FILLER_24_1262 ();
 FILLCELL_X4 FILLER_24_1270 ();
 FILLCELL_X2 FILLER_24_1274 ();
 FILLCELL_X8 FILLER_24_1285 ();
 FILLCELL_X4 FILLER_24_1293 ();
 FILLCELL_X2 FILLER_24_1297 ();
 FILLCELL_X1 FILLER_24_1299 ();
 FILLCELL_X2 FILLER_24_1308 ();
 FILLCELL_X1 FILLER_24_1310 ();
 FILLCELL_X2 FILLER_24_1319 ();
 FILLCELL_X2 FILLER_24_1332 ();
 FILLCELL_X1 FILLER_24_1334 ();
 FILLCELL_X2 FILLER_24_1350 ();
 FILLCELL_X8 FILLER_24_1355 ();
 FILLCELL_X2 FILLER_24_1363 ();
 FILLCELL_X1 FILLER_24_1365 ();
 FILLCELL_X8 FILLER_24_1379 ();
 FILLCELL_X2 FILLER_24_1387 ();
 FILLCELL_X1 FILLER_24_1389 ();
 FILLCELL_X2 FILLER_24_1404 ();
 FILLCELL_X2 FILLER_24_1410 ();
 FILLCELL_X2 FILLER_24_1417 ();
 FILLCELL_X1 FILLER_24_1419 ();
 FILLCELL_X2 FILLER_24_1439 ();
 FILLCELL_X4 FILLER_24_1446 ();
 FILLCELL_X2 FILLER_24_1450 ();
 FILLCELL_X1 FILLER_24_1452 ();
 FILLCELL_X32 FILLER_24_1457 ();
 FILLCELL_X32 FILLER_24_1489 ();
 FILLCELL_X32 FILLER_24_1521 ();
 FILLCELL_X32 FILLER_24_1553 ();
 FILLCELL_X32 FILLER_24_1585 ();
 FILLCELL_X32 FILLER_24_1617 ();
 FILLCELL_X2 FILLER_24_1649 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X4 FILLER_25_161 ();
 FILLCELL_X2 FILLER_25_165 ();
 FILLCELL_X1 FILLER_25_167 ();
 FILLCELL_X4 FILLER_25_189 ();
 FILLCELL_X1 FILLER_25_193 ();
 FILLCELL_X1 FILLER_25_198 ();
 FILLCELL_X8 FILLER_25_203 ();
 FILLCELL_X4 FILLER_25_211 ();
 FILLCELL_X2 FILLER_25_222 ();
 FILLCELL_X2 FILLER_25_243 ();
 FILLCELL_X2 FILLER_25_261 ();
 FILLCELL_X2 FILLER_25_269 ();
 FILLCELL_X8 FILLER_25_280 ();
 FILLCELL_X1 FILLER_25_288 ();
 FILLCELL_X4 FILLER_25_292 ();
 FILLCELL_X2 FILLER_25_296 ();
 FILLCELL_X4 FILLER_25_305 ();
 FILLCELL_X2 FILLER_25_309 ();
 FILLCELL_X1 FILLER_25_311 ();
 FILLCELL_X16 FILLER_25_327 ();
 FILLCELL_X8 FILLER_25_343 ();
 FILLCELL_X2 FILLER_25_351 ();
 FILLCELL_X2 FILLER_25_362 ();
 FILLCELL_X1 FILLER_25_364 ();
 FILLCELL_X4 FILLER_25_381 ();
 FILLCELL_X1 FILLER_25_385 ();
 FILLCELL_X2 FILLER_25_400 ();
 FILLCELL_X1 FILLER_25_402 ();
 FILLCELL_X2 FILLER_25_414 ();
 FILLCELL_X32 FILLER_25_436 ();
 FILLCELL_X8 FILLER_25_468 ();
 FILLCELL_X4 FILLER_25_476 ();
 FILLCELL_X1 FILLER_25_480 ();
 FILLCELL_X2 FILLER_25_508 ();
 FILLCELL_X4 FILLER_25_515 ();
 FILLCELL_X2 FILLER_25_528 ();
 FILLCELL_X4 FILLER_25_533 ();
 FILLCELL_X8 FILLER_25_551 ();
 FILLCELL_X4 FILLER_25_559 ();
 FILLCELL_X2 FILLER_25_563 ();
 FILLCELL_X4 FILLER_25_573 ();
 FILLCELL_X1 FILLER_25_577 ();
 FILLCELL_X1 FILLER_25_594 ();
 FILLCELL_X4 FILLER_25_600 ();
 FILLCELL_X2 FILLER_25_604 ();
 FILLCELL_X1 FILLER_25_606 ();
 FILLCELL_X4 FILLER_25_610 ();
 FILLCELL_X2 FILLER_25_614 ();
 FILLCELL_X2 FILLER_25_621 ();
 FILLCELL_X1 FILLER_25_623 ();
 FILLCELL_X4 FILLER_25_636 ();
 FILLCELL_X2 FILLER_25_640 ();
 FILLCELL_X2 FILLER_25_645 ();
 FILLCELL_X1 FILLER_25_647 ();
 FILLCELL_X4 FILLER_25_664 ();
 FILLCELL_X1 FILLER_25_668 ();
 FILLCELL_X1 FILLER_25_676 ();
 FILLCELL_X1 FILLER_25_701 ();
 FILLCELL_X8 FILLER_25_720 ();
 FILLCELL_X2 FILLER_25_728 ();
 FILLCELL_X4 FILLER_25_761 ();
 FILLCELL_X1 FILLER_25_765 ();
 FILLCELL_X8 FILLER_25_784 ();
 FILLCELL_X1 FILLER_25_792 ();
 FILLCELL_X4 FILLER_25_800 ();
 FILLCELL_X2 FILLER_25_804 ();
 FILLCELL_X1 FILLER_25_806 ();
 FILLCELL_X4 FILLER_25_812 ();
 FILLCELL_X4 FILLER_25_823 ();
 FILLCELL_X2 FILLER_25_827 ();
 FILLCELL_X1 FILLER_25_846 ();
 FILLCELL_X1 FILLER_25_851 ();
 FILLCELL_X2 FILLER_25_870 ();
 FILLCELL_X1 FILLER_25_883 ();
 FILLCELL_X2 FILLER_25_887 ();
 FILLCELL_X4 FILLER_25_892 ();
 FILLCELL_X2 FILLER_25_896 ();
 FILLCELL_X1 FILLER_25_912 ();
 FILLCELL_X2 FILLER_25_918 ();
 FILLCELL_X2 FILLER_25_927 ();
 FILLCELL_X1 FILLER_25_929 ();
 FILLCELL_X4 FILLER_25_933 ();
 FILLCELL_X1 FILLER_25_953 ();
 FILLCELL_X8 FILLER_25_967 ();
 FILLCELL_X2 FILLER_25_975 ();
 FILLCELL_X2 FILLER_25_985 ();
 FILLCELL_X2 FILLER_25_1000 ();
 FILLCELL_X16 FILLER_25_1015 ();
 FILLCELL_X2 FILLER_25_1031 ();
 FILLCELL_X2 FILLER_25_1042 ();
 FILLCELL_X2 FILLER_25_1061 ();
 FILLCELL_X1 FILLER_25_1063 ();
 FILLCELL_X32 FILLER_25_1082 ();
 FILLCELL_X16 FILLER_25_1114 ();
 FILLCELL_X1 FILLER_25_1130 ();
 FILLCELL_X8 FILLER_25_1138 ();
 FILLCELL_X4 FILLER_25_1149 ();
 FILLCELL_X2 FILLER_25_1153 ();
 FILLCELL_X1 FILLER_25_1166 ();
 FILLCELL_X4 FILLER_25_1170 ();
 FILLCELL_X1 FILLER_25_1174 ();
 FILLCELL_X1 FILLER_25_1209 ();
 FILLCELL_X2 FILLER_25_1227 ();
 FILLCELL_X8 FILLER_25_1236 ();
 FILLCELL_X1 FILLER_25_1244 ();
 FILLCELL_X8 FILLER_25_1248 ();
 FILLCELL_X4 FILLER_25_1256 ();
 FILLCELL_X2 FILLER_25_1260 ();
 FILLCELL_X1 FILLER_25_1262 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X2 FILLER_25_1296 ();
 FILLCELL_X1 FILLER_25_1312 ();
 FILLCELL_X4 FILLER_25_1322 ();
 FILLCELL_X2 FILLER_25_1334 ();
 FILLCELL_X4 FILLER_25_1346 ();
 FILLCELL_X2 FILLER_25_1373 ();
 FILLCELL_X2 FILLER_25_1380 ();
 FILLCELL_X1 FILLER_25_1382 ();
 FILLCELL_X4 FILLER_25_1386 ();
 FILLCELL_X2 FILLER_25_1390 ();
 FILLCELL_X1 FILLER_25_1392 ();
 FILLCELL_X16 FILLER_25_1397 ();
 FILLCELL_X8 FILLER_25_1413 ();
 FILLCELL_X1 FILLER_25_1421 ();
 FILLCELL_X4 FILLER_25_1425 ();
 FILLCELL_X2 FILLER_25_1434 ();
 FILLCELL_X1 FILLER_25_1436 ();
 FILLCELL_X8 FILLER_25_1444 ();
 FILLCELL_X32 FILLER_25_1464 ();
 FILLCELL_X32 FILLER_25_1496 ();
 FILLCELL_X32 FILLER_25_1528 ();
 FILLCELL_X32 FILLER_25_1560 ();
 FILLCELL_X32 FILLER_25_1592 ();
 FILLCELL_X16 FILLER_25_1624 ();
 FILLCELL_X8 FILLER_25_1640 ();
 FILLCELL_X2 FILLER_25_1648 ();
 FILLCELL_X1 FILLER_25_1650 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X16 FILLER_26_161 ();
 FILLCELL_X8 FILLER_26_177 ();
 FILLCELL_X2 FILLER_26_185 ();
 FILLCELL_X2 FILLER_26_190 ();
 FILLCELL_X1 FILLER_26_192 ();
 FILLCELL_X4 FILLER_26_228 ();
 FILLCELL_X1 FILLER_26_232 ();
 FILLCELL_X1 FILLER_26_241 ();
 FILLCELL_X2 FILLER_26_246 ();
 FILLCELL_X8 FILLER_26_252 ();
 FILLCELL_X4 FILLER_26_260 ();
 FILLCELL_X1 FILLER_26_270 ();
 FILLCELL_X1 FILLER_26_275 ();
 FILLCELL_X4 FILLER_26_283 ();
 FILLCELL_X2 FILLER_26_287 ();
 FILLCELL_X1 FILLER_26_289 ();
 FILLCELL_X8 FILLER_26_298 ();
 FILLCELL_X4 FILLER_26_306 ();
 FILLCELL_X1 FILLER_26_310 ();
 FILLCELL_X8 FILLER_26_318 ();
 FILLCELL_X2 FILLER_26_326 ();
 FILLCELL_X1 FILLER_26_328 ();
 FILLCELL_X4 FILLER_26_407 ();
 FILLCELL_X16 FILLER_26_438 ();
 FILLCELL_X2 FILLER_26_454 ();
 FILLCELL_X4 FILLER_26_474 ();
 FILLCELL_X2 FILLER_26_478 ();
 FILLCELL_X2 FILLER_26_487 ();
 FILLCELL_X1 FILLER_26_489 ();
 FILLCELL_X4 FILLER_26_514 ();
 FILLCELL_X1 FILLER_26_518 ();
 FILLCELL_X2 FILLER_26_526 ();
 FILLCELL_X4 FILLER_26_535 ();
 FILLCELL_X4 FILLER_26_546 ();
 FILLCELL_X4 FILLER_26_555 ();
 FILLCELL_X1 FILLER_26_576 ();
 FILLCELL_X2 FILLER_26_593 ();
 FILLCELL_X2 FILLER_26_599 ();
 FILLCELL_X1 FILLER_26_601 ();
 FILLCELL_X1 FILLER_26_625 ();
 FILLCELL_X1 FILLER_26_630 ();
 FILLCELL_X2 FILLER_26_632 ();
 FILLCELL_X1 FILLER_26_634 ();
 FILLCELL_X4 FILLER_26_651 ();
 FILLCELL_X1 FILLER_26_655 ();
 FILLCELL_X8 FILLER_26_665 ();
 FILLCELL_X2 FILLER_26_673 ();
 FILLCELL_X1 FILLER_26_675 ();
 FILLCELL_X4 FILLER_26_694 ();
 FILLCELL_X1 FILLER_26_698 ();
 FILLCELL_X32 FILLER_26_706 ();
 FILLCELL_X8 FILLER_26_738 ();
 FILLCELL_X4 FILLER_26_746 ();
 FILLCELL_X16 FILLER_26_757 ();
 FILLCELL_X4 FILLER_26_773 ();
 FILLCELL_X1 FILLER_26_777 ();
 FILLCELL_X2 FILLER_26_785 ();
 FILLCELL_X4 FILLER_26_800 ();
 FILLCELL_X16 FILLER_26_822 ();
 FILLCELL_X2 FILLER_26_838 ();
 FILLCELL_X1 FILLER_26_840 ();
 FILLCELL_X4 FILLER_26_890 ();
 FILLCELL_X1 FILLER_26_894 ();
 FILLCELL_X1 FILLER_26_929 ();
 FILLCELL_X2 FILLER_26_935 ();
 FILLCELL_X8 FILLER_26_967 ();
 FILLCELL_X4 FILLER_26_975 ();
 FILLCELL_X4 FILLER_26_1006 ();
 FILLCELL_X1 FILLER_26_1010 ();
 FILLCELL_X1 FILLER_26_1040 ();
 FILLCELL_X4 FILLER_26_1050 ();
 FILLCELL_X2 FILLER_26_1054 ();
 FILLCELL_X1 FILLER_26_1074 ();
 FILLCELL_X4 FILLER_26_1078 ();
 FILLCELL_X2 FILLER_26_1082 ();
 FILLCELL_X4 FILLER_26_1123 ();
 FILLCELL_X2 FILLER_26_1127 ();
 FILLCELL_X8 FILLER_26_1141 ();
 FILLCELL_X2 FILLER_26_1149 ();
 FILLCELL_X2 FILLER_26_1177 ();
 FILLCELL_X1 FILLER_26_1179 ();
 FILLCELL_X4 FILLER_26_1185 ();
 FILLCELL_X2 FILLER_26_1211 ();
 FILLCELL_X2 FILLER_26_1217 ();
 FILLCELL_X1 FILLER_26_1219 ();
 FILLCELL_X2 FILLER_26_1228 ();
 FILLCELL_X1 FILLER_26_1230 ();
 FILLCELL_X2 FILLER_26_1238 ();
 FILLCELL_X1 FILLER_26_1244 ();
 FILLCELL_X32 FILLER_26_1252 ();
 FILLCELL_X2 FILLER_26_1284 ();
 FILLCELL_X1 FILLER_26_1286 ();
 FILLCELL_X4 FILLER_26_1291 ();
 FILLCELL_X1 FILLER_26_1295 ();
 FILLCELL_X4 FILLER_26_1302 ();
 FILLCELL_X1 FILLER_26_1306 ();
 FILLCELL_X2 FILLER_26_1317 ();
 FILLCELL_X4 FILLER_26_1329 ();
 FILLCELL_X1 FILLER_26_1333 ();
 FILLCELL_X4 FILLER_26_1340 ();
 FILLCELL_X2 FILLER_26_1344 ();
 FILLCELL_X1 FILLER_26_1363 ();
 FILLCELL_X4 FILLER_26_1388 ();
 FILLCELL_X2 FILLER_26_1392 ();
 FILLCELL_X8 FILLER_26_1398 ();
 FILLCELL_X2 FILLER_26_1411 ();
 FILLCELL_X1 FILLER_26_1413 ();
 FILLCELL_X4 FILLER_26_1418 ();
 FILLCELL_X2 FILLER_26_1426 ();
 FILLCELL_X32 FILLER_26_1451 ();
 FILLCELL_X32 FILLER_26_1483 ();
 FILLCELL_X32 FILLER_26_1515 ();
 FILLCELL_X32 FILLER_26_1547 ();
 FILLCELL_X32 FILLER_26_1579 ();
 FILLCELL_X32 FILLER_26_1611 ();
 FILLCELL_X8 FILLER_26_1643 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X8 FILLER_27_161 ();
 FILLCELL_X4 FILLER_27_169 ();
 FILLCELL_X2 FILLER_27_173 ();
 FILLCELL_X8 FILLER_27_189 ();
 FILLCELL_X1 FILLER_27_197 ();
 FILLCELL_X8 FILLER_27_205 ();
 FILLCELL_X2 FILLER_27_213 ();
 FILLCELL_X2 FILLER_27_226 ();
 FILLCELL_X1 FILLER_27_228 ();
 FILLCELL_X4 FILLER_27_233 ();
 FILLCELL_X2 FILLER_27_237 ();
 FILLCELL_X8 FILLER_27_246 ();
 FILLCELL_X4 FILLER_27_254 ();
 FILLCELL_X2 FILLER_27_258 ();
 FILLCELL_X4 FILLER_27_267 ();
 FILLCELL_X2 FILLER_27_280 ();
 FILLCELL_X2 FILLER_27_287 ();
 FILLCELL_X1 FILLER_27_289 ();
 FILLCELL_X4 FILLER_27_293 ();
 FILLCELL_X2 FILLER_27_309 ();
 FILLCELL_X1 FILLER_27_311 ();
 FILLCELL_X1 FILLER_27_326 ();
 FILLCELL_X8 FILLER_27_331 ();
 FILLCELL_X2 FILLER_27_339 ();
 FILLCELL_X2 FILLER_27_357 ();
 FILLCELL_X4 FILLER_27_368 ();
 FILLCELL_X2 FILLER_27_372 ();
 FILLCELL_X1 FILLER_27_374 ();
 FILLCELL_X2 FILLER_27_391 ();
 FILLCELL_X8 FILLER_27_404 ();
 FILLCELL_X1 FILLER_27_412 ();
 FILLCELL_X8 FILLER_27_424 ();
 FILLCELL_X4 FILLER_27_432 ();
 FILLCELL_X16 FILLER_27_445 ();
 FILLCELL_X4 FILLER_27_461 ();
 FILLCELL_X1 FILLER_27_483 ();
 FILLCELL_X1 FILLER_27_515 ();
 FILLCELL_X1 FILLER_27_527 ();
 FILLCELL_X2 FILLER_27_546 ();
 FILLCELL_X4 FILLER_27_565 ();
 FILLCELL_X1 FILLER_27_569 ();
 FILLCELL_X2 FILLER_27_601 ();
 FILLCELL_X2 FILLER_27_648 ();
 FILLCELL_X1 FILLER_27_650 ();
 FILLCELL_X1 FILLER_27_660 ();
 FILLCELL_X4 FILLER_27_670 ();
 FILLCELL_X1 FILLER_27_674 ();
 FILLCELL_X4 FILLER_27_686 ();
 FILLCELL_X16 FILLER_27_712 ();
 FILLCELL_X8 FILLER_27_728 ();
 FILLCELL_X2 FILLER_27_743 ();
 FILLCELL_X1 FILLER_27_745 ();
 FILLCELL_X8 FILLER_27_766 ();
 FILLCELL_X4 FILLER_27_781 ();
 FILLCELL_X2 FILLER_27_785 ();
 FILLCELL_X1 FILLER_27_816 ();
 FILLCELL_X1 FILLER_27_820 ();
 FILLCELL_X1 FILLER_27_828 ();
 FILLCELL_X1 FILLER_27_835 ();
 FILLCELL_X2 FILLER_27_850 ();
 FILLCELL_X1 FILLER_27_852 ();
 FILLCELL_X1 FILLER_27_857 ();
 FILLCELL_X4 FILLER_27_863 ();
 FILLCELL_X4 FILLER_27_885 ();
 FILLCELL_X32 FILLER_27_893 ();
 FILLCELL_X8 FILLER_27_925 ();
 FILLCELL_X1 FILLER_27_933 ();
 FILLCELL_X4 FILLER_27_943 ();
 FILLCELL_X1 FILLER_27_947 ();
 FILLCELL_X16 FILLER_27_961 ();
 FILLCELL_X8 FILLER_27_977 ();
 FILLCELL_X2 FILLER_27_994 ();
 FILLCELL_X4 FILLER_27_1014 ();
 FILLCELL_X2 FILLER_27_1018 ();
 FILLCELL_X1 FILLER_27_1020 ();
 FILLCELL_X8 FILLER_27_1032 ();
 FILLCELL_X2 FILLER_27_1040 ();
 FILLCELL_X4 FILLER_27_1051 ();
 FILLCELL_X2 FILLER_27_1064 ();
 FILLCELL_X1 FILLER_27_1066 ();
 FILLCELL_X4 FILLER_27_1092 ();
 FILLCELL_X2 FILLER_27_1096 ();
 FILLCELL_X16 FILLER_27_1115 ();
 FILLCELL_X1 FILLER_27_1131 ();
 FILLCELL_X2 FILLER_27_1150 ();
 FILLCELL_X1 FILLER_27_1152 ();
 FILLCELL_X4 FILLER_27_1171 ();
 FILLCELL_X2 FILLER_27_1175 ();
 FILLCELL_X2 FILLER_27_1181 ();
 FILLCELL_X4 FILLER_27_1188 ();
 FILLCELL_X2 FILLER_27_1192 ();
 FILLCELL_X4 FILLER_27_1205 ();
 FILLCELL_X8 FILLER_27_1218 ();
 FILLCELL_X2 FILLER_27_1226 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X16 FILLER_27_1264 ();
 FILLCELL_X4 FILLER_27_1280 ();
 FILLCELL_X1 FILLER_27_1284 ();
 FILLCELL_X4 FILLER_27_1289 ();
 FILLCELL_X2 FILLER_27_1293 ();
 FILLCELL_X1 FILLER_27_1303 ();
 FILLCELL_X4 FILLER_27_1315 ();
 FILLCELL_X2 FILLER_27_1326 ();
 FILLCELL_X1 FILLER_27_1333 ();
 FILLCELL_X1 FILLER_27_1338 ();
 FILLCELL_X1 FILLER_27_1348 ();
 FILLCELL_X2 FILLER_27_1358 ();
 FILLCELL_X4 FILLER_27_1369 ();
 FILLCELL_X2 FILLER_27_1389 ();
 FILLCELL_X1 FILLER_27_1403 ();
 FILLCELL_X4 FILLER_27_1411 ();
 FILLCELL_X1 FILLER_27_1415 ();
 FILLCELL_X32 FILLER_27_1470 ();
 FILLCELL_X32 FILLER_27_1502 ();
 FILLCELL_X32 FILLER_27_1534 ();
 FILLCELL_X32 FILLER_27_1566 ();
 FILLCELL_X32 FILLER_27_1598 ();
 FILLCELL_X16 FILLER_27_1630 ();
 FILLCELL_X4 FILLER_27_1646 ();
 FILLCELL_X1 FILLER_27_1650 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X8 FILLER_28_161 ();
 FILLCELL_X4 FILLER_28_169 ();
 FILLCELL_X1 FILLER_28_173 ();
 FILLCELL_X4 FILLER_28_192 ();
 FILLCELL_X4 FILLER_28_203 ();
 FILLCELL_X1 FILLER_28_207 ();
 FILLCELL_X4 FILLER_28_226 ();
 FILLCELL_X1 FILLER_28_230 ();
 FILLCELL_X1 FILLER_28_235 ();
 FILLCELL_X1 FILLER_28_240 ();
 FILLCELL_X1 FILLER_28_246 ();
 FILLCELL_X8 FILLER_28_265 ();
 FILLCELL_X2 FILLER_28_280 ();
 FILLCELL_X1 FILLER_28_282 ();
 FILLCELL_X4 FILLER_28_286 ();
 FILLCELL_X1 FILLER_28_290 ();
 FILLCELL_X4 FILLER_28_314 ();
 FILLCELL_X2 FILLER_28_318 ();
 FILLCELL_X1 FILLER_28_320 ();
 FILLCELL_X1 FILLER_28_325 ();
 FILLCELL_X8 FILLER_28_334 ();
 FILLCELL_X2 FILLER_28_342 ();
 FILLCELL_X2 FILLER_28_358 ();
 FILLCELL_X1 FILLER_28_360 ();
 FILLCELL_X4 FILLER_28_379 ();
 FILLCELL_X2 FILLER_28_383 ();
 FILLCELL_X4 FILLER_28_403 ();
 FILLCELL_X1 FILLER_28_407 ();
 FILLCELL_X1 FILLER_28_422 ();
 FILLCELL_X2 FILLER_28_443 ();
 FILLCELL_X1 FILLER_28_445 ();
 FILLCELL_X16 FILLER_28_455 ();
 FILLCELL_X8 FILLER_28_471 ();
 FILLCELL_X4 FILLER_28_479 ();
 FILLCELL_X2 FILLER_28_483 ();
 FILLCELL_X1 FILLER_28_485 ();
 FILLCELL_X16 FILLER_28_490 ();
 FILLCELL_X8 FILLER_28_506 ();
 FILLCELL_X4 FILLER_28_514 ();
 FILLCELL_X2 FILLER_28_518 ();
 FILLCELL_X4 FILLER_28_537 ();
 FILLCELL_X2 FILLER_28_541 ();
 FILLCELL_X1 FILLER_28_547 ();
 FILLCELL_X2 FILLER_28_600 ();
 FILLCELL_X2 FILLER_28_607 ();
 FILLCELL_X2 FILLER_28_620 ();
 FILLCELL_X2 FILLER_28_632 ();
 FILLCELL_X2 FILLER_28_650 ();
 FILLCELL_X4 FILLER_28_661 ();
 FILLCELL_X2 FILLER_28_665 ();
 FILLCELL_X1 FILLER_28_667 ();
 FILLCELL_X4 FILLER_28_688 ();
 FILLCELL_X4 FILLER_28_701 ();
 FILLCELL_X2 FILLER_28_705 ();
 FILLCELL_X1 FILLER_28_707 ();
 FILLCELL_X8 FILLER_28_725 ();
 FILLCELL_X4 FILLER_28_733 ();
 FILLCELL_X2 FILLER_28_737 ();
 FILLCELL_X1 FILLER_28_739 ();
 FILLCELL_X16 FILLER_28_768 ();
 FILLCELL_X1 FILLER_28_784 ();
 FILLCELL_X4 FILLER_28_799 ();
 FILLCELL_X16 FILLER_28_815 ();
 FILLCELL_X4 FILLER_28_831 ();
 FILLCELL_X8 FILLER_28_842 ();
 FILLCELL_X4 FILLER_28_850 ();
 FILLCELL_X2 FILLER_28_869 ();
 FILLCELL_X8 FILLER_28_878 ();
 FILLCELL_X4 FILLER_28_886 ();
 FILLCELL_X2 FILLER_28_890 ();
 FILLCELL_X1 FILLER_28_892 ();
 FILLCELL_X2 FILLER_28_928 ();
 FILLCELL_X1 FILLER_28_930 ();
 FILLCELL_X8 FILLER_28_940 ();
 FILLCELL_X8 FILLER_28_955 ();
 FILLCELL_X2 FILLER_28_963 ();
 FILLCELL_X16 FILLER_28_978 ();
 FILLCELL_X4 FILLER_28_994 ();
 FILLCELL_X1 FILLER_28_998 ();
 FILLCELL_X1 FILLER_28_1010 ();
 FILLCELL_X2 FILLER_28_1018 ();
 FILLCELL_X1 FILLER_28_1020 ();
 FILLCELL_X16 FILLER_28_1037 ();
 FILLCELL_X8 FILLER_28_1053 ();
 FILLCELL_X4 FILLER_28_1061 ();
 FILLCELL_X4 FILLER_28_1082 ();
 FILLCELL_X2 FILLER_28_1086 ();
 FILLCELL_X1 FILLER_28_1088 ();
 FILLCELL_X4 FILLER_28_1109 ();
 FILLCELL_X2 FILLER_28_1113 ();
 FILLCELL_X1 FILLER_28_1137 ();
 FILLCELL_X2 FILLER_28_1141 ();
 FILLCELL_X2 FILLER_28_1152 ();
 FILLCELL_X1 FILLER_28_1154 ();
 FILLCELL_X1 FILLER_28_1159 ();
 FILLCELL_X1 FILLER_28_1164 ();
 FILLCELL_X4 FILLER_28_1198 ();
 FILLCELL_X2 FILLER_28_1202 ();
 FILLCELL_X1 FILLER_28_1204 ();
 FILLCELL_X2 FILLER_28_1210 ();
 FILLCELL_X2 FILLER_28_1218 ();
 FILLCELL_X4 FILLER_28_1223 ();
 FILLCELL_X1 FILLER_28_1227 ();
 FILLCELL_X32 FILLER_28_1233 ();
 FILLCELL_X32 FILLER_28_1265 ();
 FILLCELL_X2 FILLER_28_1297 ();
 FILLCELL_X1 FILLER_28_1303 ();
 FILLCELL_X2 FILLER_28_1323 ();
 FILLCELL_X4 FILLER_28_1329 ();
 FILLCELL_X1 FILLER_28_1333 ();
 FILLCELL_X1 FILLER_28_1338 ();
 FILLCELL_X1 FILLER_28_1367 ();
 FILLCELL_X4 FILLER_28_1375 ();
 FILLCELL_X1 FILLER_28_1379 ();
 FILLCELL_X2 FILLER_28_1384 ();
 FILLCELL_X1 FILLER_28_1386 ();
 FILLCELL_X16 FILLER_28_1392 ();
 FILLCELL_X4 FILLER_28_1408 ();
 FILLCELL_X1 FILLER_28_1412 ();
 FILLCELL_X1 FILLER_28_1451 ();
 FILLCELL_X4 FILLER_28_1455 ();
 FILLCELL_X32 FILLER_28_1466 ();
 FILLCELL_X32 FILLER_28_1498 ();
 FILLCELL_X32 FILLER_28_1530 ();
 FILLCELL_X32 FILLER_28_1562 ();
 FILLCELL_X32 FILLER_28_1594 ();
 FILLCELL_X16 FILLER_28_1626 ();
 FILLCELL_X8 FILLER_28_1642 ();
 FILLCELL_X1 FILLER_28_1650 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X8 FILLER_29_161 ();
 FILLCELL_X4 FILLER_29_169 ();
 FILLCELL_X2 FILLER_29_173 ();
 FILLCELL_X1 FILLER_29_178 ();
 FILLCELL_X8 FILLER_29_193 ();
 FILLCELL_X4 FILLER_29_201 ();
 FILLCELL_X4 FILLER_29_212 ();
 FILLCELL_X1 FILLER_29_216 ();
 FILLCELL_X2 FILLER_29_237 ();
 FILLCELL_X2 FILLER_29_248 ();
 FILLCELL_X1 FILLER_29_250 ();
 FILLCELL_X1 FILLER_29_255 ();
 FILLCELL_X2 FILLER_29_267 ();
 FILLCELL_X1 FILLER_29_269 ();
 FILLCELL_X1 FILLER_29_282 ();
 FILLCELL_X4 FILLER_29_288 ();
 FILLCELL_X1 FILLER_29_300 ();
 FILLCELL_X4 FILLER_29_305 ();
 FILLCELL_X2 FILLER_29_309 ();
 FILLCELL_X1 FILLER_29_316 ();
 FILLCELL_X2 FILLER_29_321 ();
 FILLCELL_X1 FILLER_29_323 ();
 FILLCELL_X8 FILLER_29_335 ();
 FILLCELL_X1 FILLER_29_343 ();
 FILLCELL_X2 FILLER_29_361 ();
 FILLCELL_X1 FILLER_29_363 ();
 FILLCELL_X8 FILLER_29_367 ();
 FILLCELL_X4 FILLER_29_375 ();
 FILLCELL_X2 FILLER_29_379 ();
 FILLCELL_X1 FILLER_29_381 ();
 FILLCELL_X2 FILLER_29_393 ();
 FILLCELL_X4 FILLER_29_428 ();
 FILLCELL_X16 FILLER_29_445 ();
 FILLCELL_X2 FILLER_29_461 ();
 FILLCELL_X1 FILLER_29_463 ();
 FILLCELL_X4 FILLER_29_478 ();
 FILLCELL_X2 FILLER_29_482 ();
 FILLCELL_X1 FILLER_29_484 ();
 FILLCELL_X16 FILLER_29_492 ();
 FILLCELL_X4 FILLER_29_508 ();
 FILLCELL_X1 FILLER_29_512 ();
 FILLCELL_X16 FILLER_29_526 ();
 FILLCELL_X1 FILLER_29_542 ();
 FILLCELL_X4 FILLER_29_552 ();
 FILLCELL_X1 FILLER_29_556 ();
 FILLCELL_X2 FILLER_29_562 ();
 FILLCELL_X1 FILLER_29_606 ();
 FILLCELL_X4 FILLER_29_629 ();
 FILLCELL_X4 FILLER_29_640 ();
 FILLCELL_X4 FILLER_29_651 ();
 FILLCELL_X4 FILLER_29_686 ();
 FILLCELL_X1 FILLER_29_690 ();
 FILLCELL_X32 FILLER_29_716 ();
 FILLCELL_X4 FILLER_29_748 ();
 FILLCELL_X8 FILLER_29_759 ();
 FILLCELL_X4 FILLER_29_767 ();
 FILLCELL_X8 FILLER_29_780 ();
 FILLCELL_X4 FILLER_29_788 ();
 FILLCELL_X4 FILLER_29_797 ();
 FILLCELL_X8 FILLER_29_815 ();
 FILLCELL_X4 FILLER_29_823 ();
 FILLCELL_X8 FILLER_29_836 ();
 FILLCELL_X2 FILLER_29_844 ();
 FILLCELL_X16 FILLER_29_852 ();
 FILLCELL_X4 FILLER_29_868 ();
 FILLCELL_X2 FILLER_29_872 ();
 FILLCELL_X1 FILLER_29_874 ();
 FILLCELL_X4 FILLER_29_893 ();
 FILLCELL_X2 FILLER_29_897 ();
 FILLCELL_X1 FILLER_29_899 ();
 FILLCELL_X32 FILLER_29_924 ();
 FILLCELL_X32 FILLER_29_956 ();
 FILLCELL_X4 FILLER_29_988 ();
 FILLCELL_X1 FILLER_29_992 ();
 FILLCELL_X4 FILLER_29_1011 ();
 FILLCELL_X1 FILLER_29_1015 ();
 FILLCELL_X2 FILLER_29_1045 ();
 FILLCELL_X4 FILLER_29_1131 ();
 FILLCELL_X2 FILLER_29_1135 ();
 FILLCELL_X4 FILLER_29_1148 ();
 FILLCELL_X2 FILLER_29_1152 ();
 FILLCELL_X1 FILLER_29_1154 ();
 FILLCELL_X1 FILLER_29_1157 ();
 FILLCELL_X8 FILLER_29_1171 ();
 FILLCELL_X2 FILLER_29_1179 ();
 FILLCELL_X1 FILLER_29_1181 ();
 FILLCELL_X4 FILLER_29_1189 ();
 FILLCELL_X1 FILLER_29_1193 ();
 FILLCELL_X2 FILLER_29_1219 ();
 FILLCELL_X16 FILLER_29_1232 ();
 FILLCELL_X8 FILLER_29_1248 ();
 FILLCELL_X4 FILLER_29_1256 ();
 FILLCELL_X2 FILLER_29_1260 ();
 FILLCELL_X1 FILLER_29_1262 ();
 FILLCELL_X16 FILLER_29_1264 ();
 FILLCELL_X4 FILLER_29_1280 ();
 FILLCELL_X4 FILLER_29_1291 ();
 FILLCELL_X2 FILLER_29_1299 ();
 FILLCELL_X1 FILLER_29_1305 ();
 FILLCELL_X1 FILLER_29_1313 ();
 FILLCELL_X2 FILLER_29_1318 ();
 FILLCELL_X1 FILLER_29_1329 ();
 FILLCELL_X16 FILLER_29_1358 ();
 FILLCELL_X2 FILLER_29_1374 ();
 FILLCELL_X1 FILLER_29_1376 ();
 FILLCELL_X1 FILLER_29_1380 ();
 FILLCELL_X1 FILLER_29_1393 ();
 FILLCELL_X4 FILLER_29_1401 ();
 FILLCELL_X2 FILLER_29_1405 ();
 FILLCELL_X1 FILLER_29_1407 ();
 FILLCELL_X2 FILLER_29_1416 ();
 FILLCELL_X4 FILLER_29_1424 ();
 FILLCELL_X2 FILLER_29_1428 ();
 FILLCELL_X2 FILLER_29_1439 ();
 FILLCELL_X1 FILLER_29_1441 ();
 FILLCELL_X4 FILLER_29_1454 ();
 FILLCELL_X32 FILLER_29_1465 ();
 FILLCELL_X32 FILLER_29_1497 ();
 FILLCELL_X32 FILLER_29_1529 ();
 FILLCELL_X32 FILLER_29_1561 ();
 FILLCELL_X32 FILLER_29_1593 ();
 FILLCELL_X16 FILLER_29_1625 ();
 FILLCELL_X8 FILLER_29_1641 ();
 FILLCELL_X2 FILLER_29_1649 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X8 FILLER_30_193 ();
 FILLCELL_X1 FILLER_30_225 ();
 FILLCELL_X4 FILLER_30_233 ();
 FILLCELL_X2 FILLER_30_237 ();
 FILLCELL_X1 FILLER_30_239 ();
 FILLCELL_X8 FILLER_30_244 ();
 FILLCELL_X2 FILLER_30_252 ();
 FILLCELL_X1 FILLER_30_258 ();
 FILLCELL_X2 FILLER_30_264 ();
 FILLCELL_X4 FILLER_30_284 ();
 FILLCELL_X2 FILLER_30_288 ();
 FILLCELL_X2 FILLER_30_296 ();
 FILLCELL_X4 FILLER_30_315 ();
 FILLCELL_X1 FILLER_30_319 ();
 FILLCELL_X8 FILLER_30_332 ();
 FILLCELL_X2 FILLER_30_340 ();
 FILLCELL_X1 FILLER_30_342 ();
 FILLCELL_X1 FILLER_30_382 ();
 FILLCELL_X1 FILLER_30_386 ();
 FILLCELL_X1 FILLER_30_396 ();
 FILLCELL_X2 FILLER_30_408 ();
 FILLCELL_X1 FILLER_30_410 ();
 FILLCELL_X4 FILLER_30_429 ();
 FILLCELL_X1 FILLER_30_433 ();
 FILLCELL_X16 FILLER_30_445 ();
 FILLCELL_X8 FILLER_30_461 ();
 FILLCELL_X4 FILLER_30_469 ();
 FILLCELL_X1 FILLER_30_473 ();
 FILLCELL_X1 FILLER_30_485 ();
 FILLCELL_X16 FILLER_30_493 ();
 FILLCELL_X2 FILLER_30_509 ();
 FILLCELL_X8 FILLER_30_529 ();
 FILLCELL_X1 FILLER_30_537 ();
 FILLCELL_X2 FILLER_30_554 ();
 FILLCELL_X4 FILLER_30_569 ();
 FILLCELL_X2 FILLER_30_573 ();
 FILLCELL_X1 FILLER_30_575 ();
 FILLCELL_X4 FILLER_30_592 ();
 FILLCELL_X8 FILLER_30_622 ();
 FILLCELL_X1 FILLER_30_630 ();
 FILLCELL_X2 FILLER_30_632 ();
 FILLCELL_X1 FILLER_30_672 ();
 FILLCELL_X4 FILLER_30_691 ();
 FILLCELL_X2 FILLER_30_704 ();
 FILLCELL_X1 FILLER_30_706 ();
 FILLCELL_X4 FILLER_30_714 ();
 FILLCELL_X2 FILLER_30_718 ();
 FILLCELL_X4 FILLER_30_727 ();
 FILLCELL_X2 FILLER_30_731 ();
 FILLCELL_X1 FILLER_30_733 ();
 FILLCELL_X8 FILLER_30_741 ();
 FILLCELL_X2 FILLER_30_749 ();
 FILLCELL_X8 FILLER_30_775 ();
 FILLCELL_X1 FILLER_30_783 ();
 FILLCELL_X8 FILLER_30_807 ();
 FILLCELL_X2 FILLER_30_815 ();
 FILLCELL_X1 FILLER_30_817 ();
 FILLCELL_X8 FILLER_30_836 ();
 FILLCELL_X8 FILLER_30_855 ();
 FILLCELL_X2 FILLER_30_863 ();
 FILLCELL_X1 FILLER_30_865 ();
 FILLCELL_X4 FILLER_30_871 ();
 FILLCELL_X2 FILLER_30_875 ();
 FILLCELL_X8 FILLER_30_891 ();
 FILLCELL_X4 FILLER_30_917 ();
 FILLCELL_X4 FILLER_30_939 ();
 FILLCELL_X2 FILLER_30_943 ();
 FILLCELL_X1 FILLER_30_945 ();
 FILLCELL_X4 FILLER_30_959 ();
 FILLCELL_X1 FILLER_30_963 ();
 FILLCELL_X4 FILLER_30_989 ();
 FILLCELL_X2 FILLER_30_993 ();
 FILLCELL_X1 FILLER_30_995 ();
 FILLCELL_X4 FILLER_30_1005 ();
 FILLCELL_X2 FILLER_30_1009 ();
 FILLCELL_X1 FILLER_30_1011 ();
 FILLCELL_X2 FILLER_30_1039 ();
 FILLCELL_X1 FILLER_30_1041 ();
 FILLCELL_X16 FILLER_30_1105 ();
 FILLCELL_X1 FILLER_30_1121 ();
 FILLCELL_X2 FILLER_30_1132 ();
 FILLCELL_X2 FILLER_30_1141 ();
 FILLCELL_X2 FILLER_30_1158 ();
 FILLCELL_X8 FILLER_30_1169 ();
 FILLCELL_X1 FILLER_30_1177 ();
 FILLCELL_X1 FILLER_30_1191 ();
 FILLCELL_X8 FILLER_30_1196 ();
 FILLCELL_X16 FILLER_30_1208 ();
 FILLCELL_X4 FILLER_30_1224 ();
 FILLCELL_X32 FILLER_30_1237 ();
 FILLCELL_X8 FILLER_30_1269 ();
 FILLCELL_X2 FILLER_30_1277 ();
 FILLCELL_X1 FILLER_30_1303 ();
 FILLCELL_X4 FILLER_30_1309 ();
 FILLCELL_X2 FILLER_30_1313 ();
 FILLCELL_X1 FILLER_30_1323 ();
 FILLCELL_X1 FILLER_30_1342 ();
 FILLCELL_X4 FILLER_30_1351 ();
 FILLCELL_X2 FILLER_30_1355 ();
 FILLCELL_X1 FILLER_30_1357 ();
 FILLCELL_X2 FILLER_30_1361 ();
 FILLCELL_X1 FILLER_30_1363 ();
 FILLCELL_X4 FILLER_30_1370 ();
 FILLCELL_X2 FILLER_30_1374 ();
 FILLCELL_X2 FILLER_30_1383 ();
 FILLCELL_X1 FILLER_30_1385 ();
 FILLCELL_X2 FILLER_30_1400 ();
 FILLCELL_X1 FILLER_30_1402 ();
 FILLCELL_X2 FILLER_30_1408 ();
 FILLCELL_X4 FILLER_30_1413 ();
 FILLCELL_X8 FILLER_30_1420 ();
 FILLCELL_X2 FILLER_30_1428 ();
 FILLCELL_X1 FILLER_30_1430 ();
 FILLCELL_X1 FILLER_30_1434 ();
 FILLCELL_X8 FILLER_30_1446 ();
 FILLCELL_X4 FILLER_30_1461 ();
 FILLCELL_X2 FILLER_30_1465 ();
 FILLCELL_X32 FILLER_30_1474 ();
 FILLCELL_X32 FILLER_30_1506 ();
 FILLCELL_X32 FILLER_30_1538 ();
 FILLCELL_X32 FILLER_30_1570 ();
 FILLCELL_X32 FILLER_30_1602 ();
 FILLCELL_X16 FILLER_30_1634 ();
 FILLCELL_X1 FILLER_30_1650 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X16 FILLER_31_193 ();
 FILLCELL_X4 FILLER_31_209 ();
 FILLCELL_X1 FILLER_31_213 ();
 FILLCELL_X2 FILLER_31_221 ();
 FILLCELL_X2 FILLER_31_232 ();
 FILLCELL_X1 FILLER_31_234 ();
 FILLCELL_X2 FILLER_31_238 ();
 FILLCELL_X4 FILLER_31_249 ();
 FILLCELL_X2 FILLER_31_265 ();
 FILLCELL_X2 FILLER_31_276 ();
 FILLCELL_X2 FILLER_31_285 ();
 FILLCELL_X2 FILLER_31_294 ();
 FILLCELL_X8 FILLER_31_309 ();
 FILLCELL_X2 FILLER_31_317 ();
 FILLCELL_X1 FILLER_31_319 ();
 FILLCELL_X1 FILLER_31_332 ();
 FILLCELL_X4 FILLER_31_342 ();
 FILLCELL_X1 FILLER_31_369 ();
 FILLCELL_X1 FILLER_31_384 ();
 FILLCELL_X2 FILLER_31_396 ();
 FILLCELL_X8 FILLER_31_400 ();
 FILLCELL_X4 FILLER_31_408 ();
 FILLCELL_X2 FILLER_31_412 ();
 FILLCELL_X4 FILLER_31_427 ();
 FILLCELL_X2 FILLER_31_431 ();
 FILLCELL_X16 FILLER_31_450 ();
 FILLCELL_X8 FILLER_31_466 ();
 FILLCELL_X8 FILLER_31_505 ();
 FILLCELL_X2 FILLER_31_513 ();
 FILLCELL_X1 FILLER_31_515 ();
 FILLCELL_X2 FILLER_31_523 ();
 FILLCELL_X1 FILLER_31_525 ();
 FILLCELL_X1 FILLER_31_589 ();
 FILLCELL_X1 FILLER_31_601 ();
 FILLCELL_X2 FILLER_31_605 ();
 FILLCELL_X1 FILLER_31_607 ();
 FILLCELL_X2 FILLER_31_616 ();
 FILLCELL_X1 FILLER_31_630 ();
 FILLCELL_X1 FILLER_31_656 ();
 FILLCELL_X1 FILLER_31_659 ();
 FILLCELL_X32 FILLER_31_710 ();
 FILLCELL_X8 FILLER_31_742 ();
 FILLCELL_X1 FILLER_31_750 ();
 FILLCELL_X2 FILLER_31_758 ();
 FILLCELL_X1 FILLER_31_785 ();
 FILLCELL_X4 FILLER_31_793 ();
 FILLCELL_X2 FILLER_31_823 ();
 FILLCELL_X1 FILLER_31_825 ();
 FILLCELL_X2 FILLER_31_837 ();
 FILLCELL_X2 FILLER_31_844 ();
 FILLCELL_X1 FILLER_31_846 ();
 FILLCELL_X2 FILLER_31_858 ();
 FILLCELL_X1 FILLER_31_860 ();
 FILLCELL_X1 FILLER_31_879 ();
 FILLCELL_X1 FILLER_31_886 ();
 FILLCELL_X2 FILLER_31_894 ();
 FILLCELL_X1 FILLER_31_907 ();
 FILLCELL_X2 FILLER_31_919 ();
 FILLCELL_X16 FILLER_31_930 ();
 FILLCELL_X4 FILLER_31_946 ();
 FILLCELL_X1 FILLER_31_950 ();
 FILLCELL_X16 FILLER_31_997 ();
 FILLCELL_X2 FILLER_31_1046 ();
 FILLCELL_X2 FILLER_31_1061 ();
 FILLCELL_X1 FILLER_31_1063 ();
 FILLCELL_X1 FILLER_31_1073 ();
 FILLCELL_X8 FILLER_31_1115 ();
 FILLCELL_X4 FILLER_31_1123 ();
 FILLCELL_X2 FILLER_31_1127 ();
 FILLCELL_X2 FILLER_31_1132 ();
 FILLCELL_X1 FILLER_31_1148 ();
 FILLCELL_X2 FILLER_31_1154 ();
 FILLCELL_X8 FILLER_31_1174 ();
 FILLCELL_X2 FILLER_31_1182 ();
 FILLCELL_X1 FILLER_31_1191 ();
 FILLCELL_X16 FILLER_31_1195 ();
 FILLCELL_X2 FILLER_31_1211 ();
 FILLCELL_X1 FILLER_31_1213 ();
 FILLCELL_X32 FILLER_31_1218 ();
 FILLCELL_X8 FILLER_31_1250 ();
 FILLCELL_X4 FILLER_31_1258 ();
 FILLCELL_X1 FILLER_31_1262 ();
 FILLCELL_X16 FILLER_31_1264 ();
 FILLCELL_X8 FILLER_31_1280 ();
 FILLCELL_X4 FILLER_31_1288 ();
 FILLCELL_X2 FILLER_31_1292 ();
 FILLCELL_X1 FILLER_31_1306 ();
 FILLCELL_X2 FILLER_31_1320 ();
 FILLCELL_X1 FILLER_31_1325 ();
 FILLCELL_X16 FILLER_31_1330 ();
 FILLCELL_X8 FILLER_31_1349 ();
 FILLCELL_X1 FILLER_31_1362 ();
 FILLCELL_X1 FILLER_31_1374 ();
 FILLCELL_X1 FILLER_31_1384 ();
 FILLCELL_X1 FILLER_31_1389 ();
 FILLCELL_X4 FILLER_31_1410 ();
 FILLCELL_X1 FILLER_31_1417 ();
 FILLCELL_X1 FILLER_31_1421 ();
 FILLCELL_X2 FILLER_31_1429 ();
 FILLCELL_X2 FILLER_31_1438 ();
 FILLCELL_X1 FILLER_31_1449 ();
 FILLCELL_X2 FILLER_31_1459 ();
 FILLCELL_X32 FILLER_31_1475 ();
 FILLCELL_X32 FILLER_31_1507 ();
 FILLCELL_X32 FILLER_31_1539 ();
 FILLCELL_X32 FILLER_31_1571 ();
 FILLCELL_X32 FILLER_31_1603 ();
 FILLCELL_X16 FILLER_31_1635 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X16 FILLER_32_193 ();
 FILLCELL_X8 FILLER_32_209 ();
 FILLCELL_X4 FILLER_32_217 ();
 FILLCELL_X4 FILLER_32_250 ();
 FILLCELL_X2 FILLER_32_254 ();
 FILLCELL_X1 FILLER_32_256 ();
 FILLCELL_X4 FILLER_32_275 ();
 FILLCELL_X16 FILLER_32_285 ();
 FILLCELL_X4 FILLER_32_319 ();
 FILLCELL_X2 FILLER_32_323 ();
 FILLCELL_X1 FILLER_32_325 ();
 FILLCELL_X8 FILLER_32_348 ();
 FILLCELL_X2 FILLER_32_356 ();
 FILLCELL_X1 FILLER_32_358 ();
 FILLCELL_X2 FILLER_32_415 ();
 FILLCELL_X8 FILLER_32_426 ();
 FILLCELL_X2 FILLER_32_434 ();
 FILLCELL_X1 FILLER_32_436 ();
 FILLCELL_X16 FILLER_32_447 ();
 FILLCELL_X8 FILLER_32_463 ();
 FILLCELL_X2 FILLER_32_471 ();
 FILLCELL_X1 FILLER_32_480 ();
 FILLCELL_X2 FILLER_32_488 ();
 FILLCELL_X2 FILLER_32_494 ();
 FILLCELL_X1 FILLER_32_496 ();
 FILLCELL_X8 FILLER_32_499 ();
 FILLCELL_X4 FILLER_32_507 ();
 FILLCELL_X1 FILLER_32_511 ();
 FILLCELL_X2 FILLER_32_526 ();
 FILLCELL_X1 FILLER_32_528 ();
 FILLCELL_X2 FILLER_32_536 ();
 FILLCELL_X32 FILLER_32_543 ();
 FILLCELL_X4 FILLER_32_575 ();
 FILLCELL_X2 FILLER_32_579 ();
 FILLCELL_X1 FILLER_32_581 ();
 FILLCELL_X8 FILLER_32_591 ();
 FILLCELL_X2 FILLER_32_599 ();
 FILLCELL_X4 FILLER_32_632 ();
 FILLCELL_X2 FILLER_32_636 ();
 FILLCELL_X8 FILLER_32_665 ();
 FILLCELL_X4 FILLER_32_673 ();
 FILLCELL_X2 FILLER_32_677 ();
 FILLCELL_X1 FILLER_32_679 ();
 FILLCELL_X2 FILLER_32_691 ();
 FILLCELL_X1 FILLER_32_695 ();
 FILLCELL_X2 FILLER_32_701 ();
 FILLCELL_X2 FILLER_32_714 ();
 FILLCELL_X8 FILLER_32_776 ();
 FILLCELL_X16 FILLER_32_809 ();
 FILLCELL_X4 FILLER_32_825 ();
 FILLCELL_X1 FILLER_32_829 ();
 FILLCELL_X4 FILLER_32_839 ();
 FILLCELL_X1 FILLER_32_854 ();
 FILLCELL_X1 FILLER_32_901 ();
 FILLCELL_X2 FILLER_32_913 ();
 FILLCELL_X1 FILLER_32_915 ();
 FILLCELL_X8 FILLER_32_927 ();
 FILLCELL_X4 FILLER_32_935 ();
 FILLCELL_X1 FILLER_32_939 ();
 FILLCELL_X8 FILLER_32_953 ();
 FILLCELL_X2 FILLER_32_961 ();
 FILLCELL_X1 FILLER_32_963 ();
 FILLCELL_X4 FILLER_32_982 ();
 FILLCELL_X4 FILLER_32_999 ();
 FILLCELL_X2 FILLER_32_1008 ();
 FILLCELL_X1 FILLER_32_1010 ();
 FILLCELL_X4 FILLER_32_1025 ();
 FILLCELL_X1 FILLER_32_1029 ();
 FILLCELL_X1 FILLER_32_1037 ();
 FILLCELL_X4 FILLER_32_1051 ();
 FILLCELL_X1 FILLER_32_1055 ();
 FILLCELL_X8 FILLER_32_1063 ();
 FILLCELL_X4 FILLER_32_1071 ();
 FILLCELL_X1 FILLER_32_1075 ();
 FILLCELL_X32 FILLER_32_1100 ();
 FILLCELL_X16 FILLER_32_1132 ();
 FILLCELL_X8 FILLER_32_1150 ();
 FILLCELL_X4 FILLER_32_1158 ();
 FILLCELL_X2 FILLER_32_1162 ();
 FILLCELL_X2 FILLER_32_1182 ();
 FILLCELL_X1 FILLER_32_1184 ();
 FILLCELL_X4 FILLER_32_1188 ();
 FILLCELL_X1 FILLER_32_1192 ();
 FILLCELL_X1 FILLER_32_1206 ();
 FILLCELL_X32 FILLER_32_1235 ();
 FILLCELL_X16 FILLER_32_1267 ();
 FILLCELL_X2 FILLER_32_1283 ();
 FILLCELL_X8 FILLER_32_1292 ();
 FILLCELL_X4 FILLER_32_1300 ();
 FILLCELL_X1 FILLER_32_1316 ();
 FILLCELL_X2 FILLER_32_1328 ();
 FILLCELL_X4 FILLER_32_1334 ();
 FILLCELL_X2 FILLER_32_1338 ();
 FILLCELL_X16 FILLER_32_1360 ();
 FILLCELL_X1 FILLER_32_1376 ();
 FILLCELL_X2 FILLER_32_1382 ();
 FILLCELL_X8 FILLER_32_1392 ();
 FILLCELL_X2 FILLER_32_1400 ();
 FILLCELL_X2 FILLER_32_1406 ();
 FILLCELL_X2 FILLER_32_1430 ();
 FILLCELL_X1 FILLER_32_1432 ();
 FILLCELL_X2 FILLER_32_1442 ();
 FILLCELL_X4 FILLER_32_1458 ();
 FILLCELL_X1 FILLER_32_1462 ();
 FILLCELL_X32 FILLER_32_1477 ();
 FILLCELL_X32 FILLER_32_1509 ();
 FILLCELL_X32 FILLER_32_1541 ();
 FILLCELL_X32 FILLER_32_1573 ();
 FILLCELL_X32 FILLER_32_1605 ();
 FILLCELL_X8 FILLER_32_1637 ();
 FILLCELL_X4 FILLER_32_1645 ();
 FILLCELL_X2 FILLER_32_1649 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X8 FILLER_33_225 ();
 FILLCELL_X4 FILLER_33_233 ();
 FILLCELL_X1 FILLER_33_237 ();
 FILLCELL_X8 FILLER_33_242 ();
 FILLCELL_X4 FILLER_33_274 ();
 FILLCELL_X8 FILLER_33_293 ();
 FILLCELL_X1 FILLER_33_301 ();
 FILLCELL_X4 FILLER_33_319 ();
 FILLCELL_X2 FILLER_33_323 ();
 FILLCELL_X1 FILLER_33_325 ();
 FILLCELL_X8 FILLER_33_335 ();
 FILLCELL_X1 FILLER_33_343 ();
 FILLCELL_X2 FILLER_33_362 ();
 FILLCELL_X1 FILLER_33_364 ();
 FILLCELL_X1 FILLER_33_399 ();
 FILLCELL_X16 FILLER_33_428 ();
 FILLCELL_X8 FILLER_33_444 ();
 FILLCELL_X4 FILLER_33_452 ();
 FILLCELL_X2 FILLER_33_479 ();
 FILLCELL_X1 FILLER_33_481 ();
 FILLCELL_X8 FILLER_33_495 ();
 FILLCELL_X4 FILLER_33_503 ();
 FILLCELL_X1 FILLER_33_507 ();
 FILLCELL_X2 FILLER_33_521 ();
 FILLCELL_X1 FILLER_33_523 ();
 FILLCELL_X4 FILLER_33_552 ();
 FILLCELL_X2 FILLER_33_556 ();
 FILLCELL_X4 FILLER_33_562 ();
 FILLCELL_X1 FILLER_33_566 ();
 FILLCELL_X16 FILLER_33_579 ();
 FILLCELL_X1 FILLER_33_628 ();
 FILLCELL_X1 FILLER_33_640 ();
 FILLCELL_X1 FILLER_33_646 ();
 FILLCELL_X1 FILLER_33_652 ();
 FILLCELL_X1 FILLER_33_671 ();
 FILLCELL_X2 FILLER_33_681 ();
 FILLCELL_X4 FILLER_33_692 ();
 FILLCELL_X2 FILLER_33_709 ();
 FILLCELL_X1 FILLER_33_711 ();
 FILLCELL_X32 FILLER_33_721 ();
 FILLCELL_X16 FILLER_33_791 ();
 FILLCELL_X4 FILLER_33_807 ();
 FILLCELL_X4 FILLER_33_836 ();
 FILLCELL_X2 FILLER_33_840 ();
 FILLCELL_X2 FILLER_33_851 ();
 FILLCELL_X2 FILLER_33_856 ();
 FILLCELL_X4 FILLER_33_896 ();
 FILLCELL_X2 FILLER_33_900 ();
 FILLCELL_X2 FILLER_33_911 ();
 FILLCELL_X4 FILLER_33_922 ();
 FILLCELL_X1 FILLER_33_926 ();
 FILLCELL_X8 FILLER_33_952 ();
 FILLCELL_X1 FILLER_33_960 ();
 FILLCELL_X4 FILLER_33_971 ();
 FILLCELL_X4 FILLER_33_1015 ();
 FILLCELL_X2 FILLER_33_1019 ();
 FILLCELL_X1 FILLER_33_1032 ();
 FILLCELL_X1 FILLER_33_1064 ();
 FILLCELL_X8 FILLER_33_1078 ();
 FILLCELL_X4 FILLER_33_1104 ();
 FILLCELL_X2 FILLER_33_1108 ();
 FILLCELL_X16 FILLER_33_1136 ();
 FILLCELL_X8 FILLER_33_1152 ();
 FILLCELL_X2 FILLER_33_1160 ();
 FILLCELL_X1 FILLER_33_1162 ();
 FILLCELL_X4 FILLER_33_1197 ();
 FILLCELL_X2 FILLER_33_1201 ();
 FILLCELL_X1 FILLER_33_1203 ();
 FILLCELL_X16 FILLER_33_1209 ();
 FILLCELL_X8 FILLER_33_1225 ();
 FILLCELL_X1 FILLER_33_1233 ();
 FILLCELL_X8 FILLER_33_1252 ();
 FILLCELL_X2 FILLER_33_1260 ();
 FILLCELL_X1 FILLER_33_1262 ();
 FILLCELL_X16 FILLER_33_1264 ();
 FILLCELL_X8 FILLER_33_1280 ();
 FILLCELL_X1 FILLER_33_1288 ();
 FILLCELL_X4 FILLER_33_1293 ();
 FILLCELL_X2 FILLER_33_1297 ();
 FILLCELL_X4 FILLER_33_1326 ();
 FILLCELL_X1 FILLER_33_1330 ();
 FILLCELL_X2 FILLER_33_1356 ();
 FILLCELL_X4 FILLER_33_1362 ();
 FILLCELL_X1 FILLER_33_1366 ();
 FILLCELL_X2 FILLER_33_1376 ();
 FILLCELL_X1 FILLER_33_1378 ();
 FILLCELL_X2 FILLER_33_1396 ();
 FILLCELL_X4 FILLER_33_1407 ();
 FILLCELL_X2 FILLER_33_1422 ();
 FILLCELL_X2 FILLER_33_1428 ();
 FILLCELL_X4 FILLER_33_1439 ();
 FILLCELL_X1 FILLER_33_1443 ();
 FILLCELL_X8 FILLER_33_1447 ();
 FILLCELL_X1 FILLER_33_1455 ();
 FILLCELL_X32 FILLER_33_1465 ();
 FILLCELL_X32 FILLER_33_1497 ();
 FILLCELL_X32 FILLER_33_1529 ();
 FILLCELL_X32 FILLER_33_1561 ();
 FILLCELL_X32 FILLER_33_1593 ();
 FILLCELL_X16 FILLER_33_1625 ();
 FILLCELL_X8 FILLER_33_1641 ();
 FILLCELL_X2 FILLER_33_1649 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X8 FILLER_34_225 ();
 FILLCELL_X4 FILLER_34_233 ();
 FILLCELL_X2 FILLER_34_237 ();
 FILLCELL_X8 FILLER_34_263 ();
 FILLCELL_X8 FILLER_34_297 ();
 FILLCELL_X2 FILLER_34_320 ();
 FILLCELL_X1 FILLER_34_327 ();
 FILLCELL_X2 FILLER_34_334 ();
 FILLCELL_X2 FILLER_34_363 ();
 FILLCELL_X1 FILLER_34_365 ();
 FILLCELL_X2 FILLER_34_375 ();
 FILLCELL_X1 FILLER_34_377 ();
 FILLCELL_X8 FILLER_34_390 ();
 FILLCELL_X1 FILLER_34_398 ();
 FILLCELL_X8 FILLER_34_408 ();
 FILLCELL_X4 FILLER_34_416 ();
 FILLCELL_X1 FILLER_34_420 ();
 FILLCELL_X4 FILLER_34_428 ();
 FILLCELL_X2 FILLER_34_432 ();
 FILLCELL_X2 FILLER_34_441 ();
 FILLCELL_X1 FILLER_34_443 ();
 FILLCELL_X8 FILLER_34_463 ();
 FILLCELL_X8 FILLER_34_494 ();
 FILLCELL_X2 FILLER_34_502 ();
 FILLCELL_X1 FILLER_34_504 ();
 FILLCELL_X4 FILLER_34_537 ();
 FILLCELL_X1 FILLER_34_541 ();
 FILLCELL_X1 FILLER_34_564 ();
 FILLCELL_X1 FILLER_34_569 ();
 FILLCELL_X4 FILLER_34_579 ();
 FILLCELL_X1 FILLER_34_592 ();
 FILLCELL_X2 FILLER_34_628 ();
 FILLCELL_X1 FILLER_34_630 ();
 FILLCELL_X2 FILLER_34_632 ();
 FILLCELL_X2 FILLER_34_648 ();
 FILLCELL_X1 FILLER_34_661 ();
 FILLCELL_X1 FILLER_34_671 ();
 FILLCELL_X1 FILLER_34_683 ();
 FILLCELL_X1 FILLER_34_686 ();
 FILLCELL_X16 FILLER_34_696 ();
 FILLCELL_X2 FILLER_34_712 ();
 FILLCELL_X1 FILLER_34_714 ();
 FILLCELL_X2 FILLER_34_722 ();
 FILLCELL_X4 FILLER_34_731 ();
 FILLCELL_X8 FILLER_34_742 ();
 FILLCELL_X2 FILLER_34_750 ();
 FILLCELL_X1 FILLER_34_759 ();
 FILLCELL_X1 FILLER_34_780 ();
 FILLCELL_X2 FILLER_34_784 ();
 FILLCELL_X2 FILLER_34_797 ();
 FILLCELL_X2 FILLER_34_808 ();
 FILLCELL_X4 FILLER_34_821 ();
 FILLCELL_X2 FILLER_34_825 ();
 FILLCELL_X1 FILLER_34_855 ();
 FILLCELL_X4 FILLER_34_867 ();
 FILLCELL_X2 FILLER_34_897 ();
 FILLCELL_X1 FILLER_34_899 ();
 FILLCELL_X4 FILLER_34_913 ();
 FILLCELL_X1 FILLER_34_917 ();
 FILLCELL_X4 FILLER_34_985 ();
 FILLCELL_X2 FILLER_34_989 ();
 FILLCELL_X1 FILLER_34_991 ();
 FILLCELL_X8 FILLER_34_1009 ();
 FILLCELL_X2 FILLER_34_1017 ();
 FILLCELL_X1 FILLER_34_1019 ();
 FILLCELL_X8 FILLER_34_1038 ();
 FILLCELL_X4 FILLER_34_1046 ();
 FILLCELL_X2 FILLER_34_1050 ();
 FILLCELL_X2 FILLER_34_1061 ();
 FILLCELL_X32 FILLER_34_1081 ();
 FILLCELL_X8 FILLER_34_1122 ();
 FILLCELL_X4 FILLER_34_1130 ();
 FILLCELL_X2 FILLER_34_1134 ();
 FILLCELL_X1 FILLER_34_1136 ();
 FILLCELL_X16 FILLER_34_1157 ();
 FILLCELL_X8 FILLER_34_1173 ();
 FILLCELL_X2 FILLER_34_1181 ();
 FILLCELL_X32 FILLER_34_1201 ();
 FILLCELL_X32 FILLER_34_1233 ();
 FILLCELL_X16 FILLER_34_1265 ();
 FILLCELL_X2 FILLER_34_1281 ();
 FILLCELL_X1 FILLER_34_1283 ();
 FILLCELL_X4 FILLER_34_1287 ();
 FILLCELL_X1 FILLER_34_1291 ();
 FILLCELL_X1 FILLER_34_1300 ();
 FILLCELL_X1 FILLER_34_1315 ();
 FILLCELL_X1 FILLER_34_1320 ();
 FILLCELL_X4 FILLER_34_1330 ();
 FILLCELL_X2 FILLER_34_1334 ();
 FILLCELL_X16 FILLER_34_1349 ();
 FILLCELL_X8 FILLER_34_1365 ();
 FILLCELL_X2 FILLER_34_1373 ();
 FILLCELL_X1 FILLER_34_1375 ();
 FILLCELL_X2 FILLER_34_1392 ();
 FILLCELL_X1 FILLER_34_1398 ();
 FILLCELL_X4 FILLER_34_1412 ();
 FILLCELL_X8 FILLER_34_1429 ();
 FILLCELL_X2 FILLER_34_1437 ();
 FILLCELL_X1 FILLER_34_1459 ();
 FILLCELL_X1 FILLER_34_1478 ();
 FILLCELL_X32 FILLER_34_1483 ();
 FILLCELL_X32 FILLER_34_1515 ();
 FILLCELL_X32 FILLER_34_1547 ();
 FILLCELL_X32 FILLER_34_1579 ();
 FILLCELL_X32 FILLER_34_1611 ();
 FILLCELL_X8 FILLER_34_1643 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X16 FILLER_35_257 ();
 FILLCELL_X4 FILLER_35_273 ();
 FILLCELL_X8 FILLER_35_284 ();
 FILLCELL_X2 FILLER_35_292 ();
 FILLCELL_X8 FILLER_35_299 ();
 FILLCELL_X4 FILLER_35_307 ();
 FILLCELL_X16 FILLER_35_324 ();
 FILLCELL_X8 FILLER_35_340 ();
 FILLCELL_X2 FILLER_35_348 ();
 FILLCELL_X1 FILLER_35_350 ();
 FILLCELL_X8 FILLER_35_365 ();
 FILLCELL_X2 FILLER_35_373 ();
 FILLCELL_X1 FILLER_35_375 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X8 FILLER_35_513 ();
 FILLCELL_X2 FILLER_35_532 ();
 FILLCELL_X1 FILLER_35_543 ();
 FILLCELL_X8 FILLER_35_551 ();
 FILLCELL_X4 FILLER_35_559 ();
 FILLCELL_X2 FILLER_35_595 ();
 FILLCELL_X1 FILLER_35_637 ();
 FILLCELL_X2 FILLER_35_665 ();
 FILLCELL_X1 FILLER_35_667 ();
 FILLCELL_X1 FILLER_35_677 ();
 FILLCELL_X16 FILLER_35_685 ();
 FILLCELL_X4 FILLER_35_701 ();
 FILLCELL_X2 FILLER_35_710 ();
 FILLCELL_X2 FILLER_35_723 ();
 FILLCELL_X1 FILLER_35_725 ();
 FILLCELL_X2 FILLER_35_736 ();
 FILLCELL_X2 FILLER_35_751 ();
 FILLCELL_X1 FILLER_35_753 ();
 FILLCELL_X1 FILLER_35_768 ();
 FILLCELL_X1 FILLER_35_778 ();
 FILLCELL_X1 FILLER_35_791 ();
 FILLCELL_X2 FILLER_35_812 ();
 FILLCELL_X16 FILLER_35_821 ();
 FILLCELL_X2 FILLER_35_855 ();
 FILLCELL_X1 FILLER_35_857 ();
 FILLCELL_X32 FILLER_35_877 ();
 FILLCELL_X4 FILLER_35_909 ();
 FILLCELL_X2 FILLER_35_913 ();
 FILLCELL_X1 FILLER_35_940 ();
 FILLCELL_X1 FILLER_35_947 ();
 FILLCELL_X1 FILLER_35_961 ();
 FILLCELL_X8 FILLER_35_969 ();
 FILLCELL_X1 FILLER_35_977 ();
 FILLCELL_X2 FILLER_35_985 ();
 FILLCELL_X2 FILLER_35_1010 ();
 FILLCELL_X1 FILLER_35_1012 ();
 FILLCELL_X8 FILLER_35_1043 ();
 FILLCELL_X1 FILLER_35_1051 ();
 FILLCELL_X32 FILLER_35_1070 ();
 FILLCELL_X8 FILLER_35_1102 ();
 FILLCELL_X2 FILLER_35_1110 ();
 FILLCELL_X2 FILLER_35_1125 ();
 FILLCELL_X1 FILLER_35_1127 ();
 FILLCELL_X16 FILLER_35_1160 ();
 FILLCELL_X2 FILLER_35_1176 ();
 FILLCELL_X32 FILLER_35_1198 ();
 FILLCELL_X32 FILLER_35_1230 ();
 FILLCELL_X1 FILLER_35_1262 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X2 FILLER_35_1315 ();
 FILLCELL_X1 FILLER_35_1317 ();
 FILLCELL_X8 FILLER_35_1321 ();
 FILLCELL_X1 FILLER_35_1329 ();
 FILLCELL_X2 FILLER_35_1344 ();
 FILLCELL_X1 FILLER_35_1346 ();
 FILLCELL_X1 FILLER_35_1351 ();
 FILLCELL_X1 FILLER_35_1356 ();
 FILLCELL_X1 FILLER_35_1362 ();
 FILLCELL_X1 FILLER_35_1387 ();
 FILLCELL_X4 FILLER_35_1392 ();
 FILLCELL_X1 FILLER_35_1406 ();
 FILLCELL_X1 FILLER_35_1410 ();
 FILLCELL_X2 FILLER_35_1420 ();
 FILLCELL_X1 FILLER_35_1422 ();
 FILLCELL_X4 FILLER_35_1429 ();
 FILLCELL_X2 FILLER_35_1440 ();
 FILLCELL_X1 FILLER_35_1442 ();
 FILLCELL_X32 FILLER_35_1461 ();
 FILLCELL_X32 FILLER_35_1493 ();
 FILLCELL_X32 FILLER_35_1525 ();
 FILLCELL_X32 FILLER_35_1557 ();
 FILLCELL_X32 FILLER_35_1589 ();
 FILLCELL_X16 FILLER_35_1621 ();
 FILLCELL_X8 FILLER_35_1637 ();
 FILLCELL_X4 FILLER_35_1645 ();
 FILLCELL_X2 FILLER_35_1649 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X8 FILLER_36_225 ();
 FILLCELL_X16 FILLER_36_237 ();
 FILLCELL_X8 FILLER_36_253 ();
 FILLCELL_X4 FILLER_36_261 ();
 FILLCELL_X1 FILLER_36_265 ();
 FILLCELL_X2 FILLER_36_305 ();
 FILLCELL_X1 FILLER_36_307 ();
 FILLCELL_X1 FILLER_36_312 ();
 FILLCELL_X4 FILLER_36_324 ();
 FILLCELL_X1 FILLER_36_328 ();
 FILLCELL_X4 FILLER_36_336 ();
 FILLCELL_X1 FILLER_36_345 ();
 FILLCELL_X1 FILLER_36_350 ();
 FILLCELL_X2 FILLER_36_355 ();
 FILLCELL_X1 FILLER_36_357 ();
 FILLCELL_X8 FILLER_36_363 ();
 FILLCELL_X2 FILLER_36_371 ();
 FILLCELL_X1 FILLER_36_373 ();
 FILLCELL_X4 FILLER_36_385 ();
 FILLCELL_X8 FILLER_36_408 ();
 FILLCELL_X4 FILLER_36_416 ();
 FILLCELL_X1 FILLER_36_420 ();
 FILLCELL_X2 FILLER_36_467 ();
 FILLCELL_X4 FILLER_36_472 ();
 FILLCELL_X4 FILLER_36_480 ();
 FILLCELL_X1 FILLER_36_484 ();
 FILLCELL_X2 FILLER_36_487 ();
 FILLCELL_X1 FILLER_36_489 ();
 FILLCELL_X4 FILLER_36_515 ();
 FILLCELL_X1 FILLER_36_519 ();
 FILLCELL_X2 FILLER_36_523 ();
 FILLCELL_X1 FILLER_36_525 ();
 FILLCELL_X4 FILLER_36_548 ();
 FILLCELL_X4 FILLER_36_561 ();
 FILLCELL_X2 FILLER_36_565 ();
 FILLCELL_X1 FILLER_36_567 ();
 FILLCELL_X2 FILLER_36_581 ();
 FILLCELL_X1 FILLER_36_583 ();
 FILLCELL_X4 FILLER_36_587 ();
 FILLCELL_X1 FILLER_36_591 ();
 FILLCELL_X4 FILLER_36_610 ();
 FILLCELL_X2 FILLER_36_623 ();
 FILLCELL_X1 FILLER_36_625 ();
 FILLCELL_X1 FILLER_36_632 ();
 FILLCELL_X2 FILLER_36_642 ();
 FILLCELL_X4 FILLER_36_662 ();
 FILLCELL_X8 FILLER_36_683 ();
 FILLCELL_X4 FILLER_36_691 ();
 FILLCELL_X4 FILLER_36_708 ();
 FILLCELL_X2 FILLER_36_712 ();
 FILLCELL_X1 FILLER_36_714 ();
 FILLCELL_X16 FILLER_36_722 ();
 FILLCELL_X1 FILLER_36_738 ();
 FILLCELL_X4 FILLER_36_750 ();
 FILLCELL_X2 FILLER_36_754 ();
 FILLCELL_X1 FILLER_36_756 ();
 FILLCELL_X4 FILLER_36_769 ();
 FILLCELL_X1 FILLER_36_773 ();
 FILLCELL_X1 FILLER_36_794 ();
 FILLCELL_X4 FILLER_36_806 ();
 FILLCELL_X2 FILLER_36_810 ();
 FILLCELL_X8 FILLER_36_830 ();
 FILLCELL_X8 FILLER_36_849 ();
 FILLCELL_X2 FILLER_36_857 ();
 FILLCELL_X32 FILLER_36_868 ();
 FILLCELL_X4 FILLER_36_900 ();
 FILLCELL_X1 FILLER_36_904 ();
 FILLCELL_X16 FILLER_36_923 ();
 FILLCELL_X8 FILLER_36_939 ();
 FILLCELL_X1 FILLER_36_947 ();
 FILLCELL_X1 FILLER_36_966 ();
 FILLCELL_X1 FILLER_36_973 ();
 FILLCELL_X2 FILLER_36_997 ();
 FILLCELL_X2 FILLER_36_1005 ();
 FILLCELL_X4 FILLER_36_1031 ();
 FILLCELL_X1 FILLER_36_1035 ();
 FILLCELL_X4 FILLER_36_1042 ();
 FILLCELL_X1 FILLER_36_1046 ();
 FILLCELL_X4 FILLER_36_1060 ();
 FILLCELL_X2 FILLER_36_1064 ();
 FILLCELL_X8 FILLER_36_1078 ();
 FILLCELL_X4 FILLER_36_1108 ();
 FILLCELL_X8 FILLER_36_1141 ();
 FILLCELL_X4 FILLER_36_1194 ();
 FILLCELL_X2 FILLER_36_1198 ();
 FILLCELL_X1 FILLER_36_1200 ();
 FILLCELL_X4 FILLER_36_1208 ();
 FILLCELL_X2 FILLER_36_1212 ();
 FILLCELL_X1 FILLER_36_1214 ();
 FILLCELL_X16 FILLER_36_1240 ();
 FILLCELL_X8 FILLER_36_1256 ();
 FILLCELL_X4 FILLER_36_1264 ();
 FILLCELL_X2 FILLER_36_1268 ();
 FILLCELL_X1 FILLER_36_1270 ();
 FILLCELL_X8 FILLER_36_1289 ();
 FILLCELL_X1 FILLER_36_1297 ();
 FILLCELL_X4 FILLER_36_1307 ();
 FILLCELL_X2 FILLER_36_1311 ();
 FILLCELL_X1 FILLER_36_1313 ();
 FILLCELL_X2 FILLER_36_1320 ();
 FILLCELL_X2 FILLER_36_1325 ();
 FILLCELL_X1 FILLER_36_1327 ();
 FILLCELL_X4 FILLER_36_1331 ();
 FILLCELL_X2 FILLER_36_1335 ();
 FILLCELL_X4 FILLER_36_1348 ();
 FILLCELL_X2 FILLER_36_1364 ();
 FILLCELL_X4 FILLER_36_1383 ();
 FILLCELL_X1 FILLER_36_1387 ();
 FILLCELL_X1 FILLER_36_1438 ();
 FILLCELL_X1 FILLER_36_1444 ();
 FILLCELL_X1 FILLER_36_1450 ();
 FILLCELL_X1 FILLER_36_1460 ();
 FILLCELL_X32 FILLER_36_1477 ();
 FILLCELL_X32 FILLER_36_1509 ();
 FILLCELL_X32 FILLER_36_1541 ();
 FILLCELL_X32 FILLER_36_1573 ();
 FILLCELL_X32 FILLER_36_1605 ();
 FILLCELL_X8 FILLER_36_1637 ();
 FILLCELL_X4 FILLER_36_1645 ();
 FILLCELL_X2 FILLER_36_1649 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X16 FILLER_37_193 ();
 FILLCELL_X8 FILLER_37_209 ();
 FILLCELL_X4 FILLER_37_217 ();
 FILLCELL_X16 FILLER_37_248 ();
 FILLCELL_X1 FILLER_37_264 ();
 FILLCELL_X8 FILLER_37_274 ();
 FILLCELL_X4 FILLER_37_282 ();
 FILLCELL_X8 FILLER_37_326 ();
 FILLCELL_X2 FILLER_37_334 ();
 FILLCELL_X1 FILLER_37_357 ();
 FILLCELL_X2 FILLER_37_368 ();
 FILLCELL_X1 FILLER_37_408 ();
 FILLCELL_X4 FILLER_37_429 ();
 FILLCELL_X1 FILLER_37_433 ();
 FILLCELL_X4 FILLER_37_463 ();
 FILLCELL_X2 FILLER_37_467 ();
 FILLCELL_X1 FILLER_37_484 ();
 FILLCELL_X2 FILLER_37_488 ();
 FILLCELL_X1 FILLER_37_490 ();
 FILLCELL_X1 FILLER_37_494 ();
 FILLCELL_X2 FILLER_37_499 ();
 FILLCELL_X2 FILLER_37_505 ();
 FILLCELL_X16 FILLER_37_511 ();
 FILLCELL_X2 FILLER_37_527 ();
 FILLCELL_X1 FILLER_37_529 ();
 FILLCELL_X1 FILLER_37_548 ();
 FILLCELL_X8 FILLER_37_563 ();
 FILLCELL_X2 FILLER_37_571 ();
 FILLCELL_X16 FILLER_37_593 ();
 FILLCELL_X2 FILLER_37_663 ();
 FILLCELL_X2 FILLER_37_676 ();
 FILLCELL_X1 FILLER_37_678 ();
 FILLCELL_X4 FILLER_37_698 ();
 FILLCELL_X1 FILLER_37_702 ();
 FILLCELL_X8 FILLER_37_708 ();
 FILLCELL_X4 FILLER_37_723 ();
 FILLCELL_X2 FILLER_37_727 ();
 FILLCELL_X8 FILLER_37_733 ();
 FILLCELL_X32 FILLER_37_754 ();
 FILLCELL_X1 FILLER_37_786 ();
 FILLCELL_X8 FILLER_37_816 ();
 FILLCELL_X4 FILLER_37_869 ();
 FILLCELL_X1 FILLER_37_873 ();
 FILLCELL_X8 FILLER_37_898 ();
 FILLCELL_X4 FILLER_37_906 ();
 FILLCELL_X1 FILLER_37_910 ();
 FILLCELL_X16 FILLER_37_918 ();
 FILLCELL_X1 FILLER_37_934 ();
 FILLCELL_X4 FILLER_37_960 ();
 FILLCELL_X1 FILLER_37_964 ();
 FILLCELL_X8 FILLER_37_968 ();
 FILLCELL_X2 FILLER_37_976 ();
 FILLCELL_X1 FILLER_37_978 ();
 FILLCELL_X4 FILLER_37_1002 ();
 FILLCELL_X4 FILLER_37_1011 ();
 FILLCELL_X1 FILLER_37_1015 ();
 FILLCELL_X1 FILLER_37_1031 ();
 FILLCELL_X8 FILLER_37_1054 ();
 FILLCELL_X4 FILLER_37_1062 ();
 FILLCELL_X8 FILLER_37_1093 ();
 FILLCELL_X2 FILLER_37_1101 ();
 FILLCELL_X1 FILLER_37_1103 ();
 FILLCELL_X4 FILLER_37_1109 ();
 FILLCELL_X8 FILLER_37_1119 ();
 FILLCELL_X2 FILLER_37_1127 ();
 FILLCELL_X4 FILLER_37_1133 ();
 FILLCELL_X1 FILLER_37_1137 ();
 FILLCELL_X8 FILLER_37_1144 ();
 FILLCELL_X2 FILLER_37_1152 ();
 FILLCELL_X1 FILLER_37_1154 ();
 FILLCELL_X4 FILLER_37_1161 ();
 FILLCELL_X2 FILLER_37_1165 ();
 FILLCELL_X1 FILLER_37_1173 ();
 FILLCELL_X1 FILLER_37_1181 ();
 FILLCELL_X16 FILLER_37_1214 ();
 FILLCELL_X2 FILLER_37_1230 ();
 FILLCELL_X1 FILLER_37_1232 ();
 FILLCELL_X2 FILLER_37_1260 ();
 FILLCELL_X1 FILLER_37_1262 ();
 FILLCELL_X16 FILLER_37_1264 ();
 FILLCELL_X4 FILLER_37_1280 ();
 FILLCELL_X2 FILLER_37_1284 ();
 FILLCELL_X1 FILLER_37_1286 ();
 FILLCELL_X8 FILLER_37_1321 ();
 FILLCELL_X2 FILLER_37_1333 ();
 FILLCELL_X1 FILLER_37_1335 ();
 FILLCELL_X1 FILLER_37_1343 ();
 FILLCELL_X1 FILLER_37_1354 ();
 FILLCELL_X4 FILLER_37_1383 ();
 FILLCELL_X2 FILLER_37_1387 ();
 FILLCELL_X1 FILLER_37_1393 ();
 FILLCELL_X1 FILLER_37_1405 ();
 FILLCELL_X1 FILLER_37_1411 ();
 FILLCELL_X4 FILLER_37_1426 ();
 FILLCELL_X1 FILLER_37_1448 ();
 FILLCELL_X8 FILLER_37_1467 ();
 FILLCELL_X1 FILLER_37_1475 ();
 FILLCELL_X32 FILLER_37_1483 ();
 FILLCELL_X32 FILLER_37_1515 ();
 FILLCELL_X32 FILLER_37_1547 ();
 FILLCELL_X32 FILLER_37_1579 ();
 FILLCELL_X32 FILLER_37_1611 ();
 FILLCELL_X8 FILLER_37_1643 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X16 FILLER_38_193 ();
 FILLCELL_X8 FILLER_38_209 ();
 FILLCELL_X1 FILLER_38_217 ();
 FILLCELL_X1 FILLER_38_236 ();
 FILLCELL_X8 FILLER_38_248 ();
 FILLCELL_X2 FILLER_38_256 ();
 FILLCELL_X1 FILLER_38_258 ();
 FILLCELL_X16 FILLER_38_271 ();
 FILLCELL_X8 FILLER_38_287 ();
 FILLCELL_X1 FILLER_38_304 ();
 FILLCELL_X2 FILLER_38_321 ();
 FILLCELL_X2 FILLER_38_344 ();
 FILLCELL_X1 FILLER_38_418 ();
 FILLCELL_X4 FILLER_38_428 ();
 FILLCELL_X4 FILLER_38_434 ();
 FILLCELL_X1 FILLER_38_438 ();
 FILLCELL_X8 FILLER_38_456 ();
 FILLCELL_X2 FILLER_38_464 ();
 FILLCELL_X4 FILLER_38_486 ();
 FILLCELL_X16 FILLER_38_509 ();
 FILLCELL_X4 FILLER_38_555 ();
 FILLCELL_X1 FILLER_38_559 ();
 FILLCELL_X32 FILLER_38_580 ();
 FILLCELL_X4 FILLER_38_612 ();
 FILLCELL_X2 FILLER_38_616 ();
 FILLCELL_X8 FILLER_38_620 ();
 FILLCELL_X2 FILLER_38_628 ();
 FILLCELL_X1 FILLER_38_630 ();
 FILLCELL_X4 FILLER_38_637 ();
 FILLCELL_X2 FILLER_38_641 ();
 FILLCELL_X16 FILLER_38_652 ();
 FILLCELL_X8 FILLER_38_671 ();
 FILLCELL_X8 FILLER_38_683 ();
 FILLCELL_X4 FILLER_38_691 ();
 FILLCELL_X2 FILLER_38_695 ();
 FILLCELL_X1 FILLER_38_697 ();
 FILLCELL_X4 FILLER_38_734 ();
 FILLCELL_X1 FILLER_38_755 ();
 FILLCELL_X8 FILLER_38_781 ();
 FILLCELL_X8 FILLER_38_806 ();
 FILLCELL_X1 FILLER_38_814 ();
 FILLCELL_X2 FILLER_38_824 ();
 FILLCELL_X8 FILLER_38_833 ();
 FILLCELL_X4 FILLER_38_841 ();
 FILLCELL_X2 FILLER_38_845 ();
 FILLCELL_X1 FILLER_38_847 ();
 FILLCELL_X2 FILLER_38_866 ();
 FILLCELL_X1 FILLER_38_868 ();
 FILLCELL_X2 FILLER_38_887 ();
 FILLCELL_X1 FILLER_38_889 ();
 FILLCELL_X2 FILLER_38_908 ();
 FILLCELL_X4 FILLER_38_917 ();
 FILLCELL_X1 FILLER_38_921 ();
 FILLCELL_X4 FILLER_38_953 ();
 FILLCELL_X2 FILLER_38_957 ();
 FILLCELL_X4 FILLER_38_967 ();
 FILLCELL_X2 FILLER_38_971 ();
 FILLCELL_X8 FILLER_38_976 ();
 FILLCELL_X1 FILLER_38_984 ();
 FILLCELL_X4 FILLER_38_988 ();
 FILLCELL_X1 FILLER_38_992 ();
 FILLCELL_X8 FILLER_38_998 ();
 FILLCELL_X4 FILLER_38_1006 ();
 FILLCELL_X2 FILLER_38_1010 ();
 FILLCELL_X1 FILLER_38_1012 ();
 FILLCELL_X4 FILLER_38_1016 ();
 FILLCELL_X4 FILLER_38_1029 ();
 FILLCELL_X1 FILLER_38_1033 ();
 FILLCELL_X2 FILLER_38_1054 ();
 FILLCELL_X4 FILLER_38_1061 ();
 FILLCELL_X1 FILLER_38_1065 ();
 FILLCELL_X16 FILLER_38_1075 ();
 FILLCELL_X1 FILLER_38_1091 ();
 FILLCELL_X16 FILLER_38_1109 ();
 FILLCELL_X8 FILLER_38_1125 ();
 FILLCELL_X2 FILLER_38_1133 ();
 FILLCELL_X8 FILLER_38_1183 ();
 FILLCELL_X2 FILLER_38_1198 ();
 FILLCELL_X1 FILLER_38_1200 ();
 FILLCELL_X1 FILLER_38_1206 ();
 FILLCELL_X16 FILLER_38_1261 ();
 FILLCELL_X8 FILLER_38_1277 ();
 FILLCELL_X2 FILLER_38_1285 ();
 FILLCELL_X1 FILLER_38_1287 ();
 FILLCELL_X8 FILLER_38_1300 ();
 FILLCELL_X2 FILLER_38_1308 ();
 FILLCELL_X2 FILLER_38_1320 ();
 FILLCELL_X2 FILLER_38_1329 ();
 FILLCELL_X1 FILLER_38_1335 ();
 FILLCELL_X2 FILLER_38_1353 ();
 FILLCELL_X2 FILLER_38_1368 ();
 FILLCELL_X1 FILLER_38_1370 ();
 FILLCELL_X2 FILLER_38_1387 ();
 FILLCELL_X1 FILLER_38_1394 ();
 FILLCELL_X1 FILLER_38_1412 ();
 FILLCELL_X4 FILLER_38_1443 ();
 FILLCELL_X2 FILLER_38_1447 ();
 FILLCELL_X32 FILLER_38_1456 ();
 FILLCELL_X32 FILLER_38_1488 ();
 FILLCELL_X32 FILLER_38_1520 ();
 FILLCELL_X32 FILLER_38_1552 ();
 FILLCELL_X32 FILLER_38_1584 ();
 FILLCELL_X32 FILLER_38_1616 ();
 FILLCELL_X2 FILLER_38_1648 ();
 FILLCELL_X1 FILLER_38_1650 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X16 FILLER_39_193 ();
 FILLCELL_X8 FILLER_39_209 ();
 FILLCELL_X4 FILLER_39_217 ();
 FILLCELL_X1 FILLER_39_221 ();
 FILLCELL_X4 FILLER_39_256 ();
 FILLCELL_X2 FILLER_39_260 ();
 FILLCELL_X1 FILLER_39_268 ();
 FILLCELL_X8 FILLER_39_272 ();
 FILLCELL_X2 FILLER_39_300 ();
 FILLCELL_X16 FILLER_39_321 ();
 FILLCELL_X8 FILLER_39_337 ();
 FILLCELL_X2 FILLER_39_345 ();
 FILLCELL_X1 FILLER_39_347 ();
 FILLCELL_X2 FILLER_39_368 ();
 FILLCELL_X8 FILLER_39_376 ();
 FILLCELL_X1 FILLER_39_384 ();
 FILLCELL_X1 FILLER_39_392 ();
 FILLCELL_X2 FILLER_39_397 ();
 FILLCELL_X2 FILLER_39_406 ();
 FILLCELL_X2 FILLER_39_414 ();
 FILLCELL_X4 FILLER_39_420 ();
 FILLCELL_X4 FILLER_39_463 ();
 FILLCELL_X1 FILLER_39_467 ();
 FILLCELL_X1 FILLER_39_471 ();
 FILLCELL_X1 FILLER_39_483 ();
 FILLCELL_X2 FILLER_39_488 ();
 FILLCELL_X1 FILLER_39_500 ();
 FILLCELL_X2 FILLER_39_508 ();
 FILLCELL_X1 FILLER_39_510 ();
 FILLCELL_X8 FILLER_39_515 ();
 FILLCELL_X4 FILLER_39_523 ();
 FILLCELL_X1 FILLER_39_527 ();
 FILLCELL_X2 FILLER_39_535 ();
 FILLCELL_X16 FILLER_39_549 ();
 FILLCELL_X1 FILLER_39_570 ();
 FILLCELL_X4 FILLER_39_573 ();
 FILLCELL_X1 FILLER_39_577 ();
 FILLCELL_X4 FILLER_39_582 ();
 FILLCELL_X1 FILLER_39_586 ();
 FILLCELL_X4 FILLER_39_597 ();
 FILLCELL_X2 FILLER_39_601 ();
 FILLCELL_X1 FILLER_39_603 ();
 FILLCELL_X8 FILLER_39_635 ();
 FILLCELL_X1 FILLER_39_643 ();
 FILLCELL_X8 FILLER_39_666 ();
 FILLCELL_X2 FILLER_39_674 ();
 FILLCELL_X8 FILLER_39_703 ();
 FILLCELL_X4 FILLER_39_711 ();
 FILLCELL_X2 FILLER_39_715 ();
 FILLCELL_X1 FILLER_39_717 ();
 FILLCELL_X1 FILLER_39_727 ();
 FILLCELL_X4 FILLER_39_767 ();
 FILLCELL_X2 FILLER_39_771 ();
 FILLCELL_X1 FILLER_39_773 ();
 FILLCELL_X8 FILLER_39_796 ();
 FILLCELL_X2 FILLER_39_804 ();
 FILLCELL_X1 FILLER_39_806 ();
 FILLCELL_X4 FILLER_39_821 ();
 FILLCELL_X2 FILLER_39_825 ();
 FILLCELL_X4 FILLER_39_833 ();
 FILLCELL_X2 FILLER_39_837 ();
 FILLCELL_X1 FILLER_39_839 ();
 FILLCELL_X1 FILLER_39_864 ();
 FILLCELL_X2 FILLER_39_878 ();
 FILLCELL_X4 FILLER_39_893 ();
 FILLCELL_X1 FILLER_39_897 ();
 FILLCELL_X16 FILLER_39_910 ();
 FILLCELL_X2 FILLER_39_926 ();
 FILLCELL_X16 FILLER_39_941 ();
 FILLCELL_X8 FILLER_39_957 ();
 FILLCELL_X4 FILLER_39_965 ();
 FILLCELL_X1 FILLER_39_969 ();
 FILLCELL_X4 FILLER_39_982 ();
 FILLCELL_X1 FILLER_39_1001 ();
 FILLCELL_X4 FILLER_39_1007 ();
 FILLCELL_X2 FILLER_39_1016 ();
 FILLCELL_X8 FILLER_39_1027 ();
 FILLCELL_X4 FILLER_39_1045 ();
 FILLCELL_X1 FILLER_39_1049 ();
 FILLCELL_X2 FILLER_39_1055 ();
 FILLCELL_X2 FILLER_39_1062 ();
 FILLCELL_X1 FILLER_39_1064 ();
 FILLCELL_X1 FILLER_39_1067 ();
 FILLCELL_X2 FILLER_39_1105 ();
 FILLCELL_X2 FILLER_39_1156 ();
 FILLCELL_X8 FILLER_39_1174 ();
 FILLCELL_X2 FILLER_39_1209 ();
 FILLCELL_X8 FILLER_39_1218 ();
 FILLCELL_X4 FILLER_39_1226 ();
 FILLCELL_X2 FILLER_39_1230 ();
 FILLCELL_X16 FILLER_39_1246 ();
 FILLCELL_X1 FILLER_39_1262 ();
 FILLCELL_X8 FILLER_39_1284 ();
 FILLCELL_X2 FILLER_39_1292 ();
 FILLCELL_X1 FILLER_39_1294 ();
 FILLCELL_X4 FILLER_39_1313 ();
 FILLCELL_X2 FILLER_39_1317 ();
 FILLCELL_X1 FILLER_39_1322 ();
 FILLCELL_X1 FILLER_39_1327 ();
 FILLCELL_X1 FILLER_39_1344 ();
 FILLCELL_X4 FILLER_39_1354 ();
 FILLCELL_X1 FILLER_39_1358 ();
 FILLCELL_X8 FILLER_39_1377 ();
 FILLCELL_X4 FILLER_39_1385 ();
 FILLCELL_X2 FILLER_39_1389 ();
 FILLCELL_X2 FILLER_39_1409 ();
 FILLCELL_X1 FILLER_39_1425 ();
 FILLCELL_X4 FILLER_39_1429 ();
 FILLCELL_X1 FILLER_39_1433 ();
 FILLCELL_X2 FILLER_39_1443 ();
 FILLCELL_X1 FILLER_39_1445 ();
 FILLCELL_X1 FILLER_39_1450 ();
 FILLCELL_X32 FILLER_39_1458 ();
 FILLCELL_X32 FILLER_39_1490 ();
 FILLCELL_X32 FILLER_39_1522 ();
 FILLCELL_X32 FILLER_39_1554 ();
 FILLCELL_X32 FILLER_39_1586 ();
 FILLCELL_X32 FILLER_39_1618 ();
 FILLCELL_X1 FILLER_39_1650 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X16 FILLER_40_193 ();
 FILLCELL_X8 FILLER_40_209 ();
 FILLCELL_X1 FILLER_40_217 ();
 FILLCELL_X1 FILLER_40_225 ();
 FILLCELL_X8 FILLER_40_241 ();
 FILLCELL_X2 FILLER_40_249 ();
 FILLCELL_X1 FILLER_40_251 ();
 FILLCELL_X4 FILLER_40_279 ();
 FILLCELL_X2 FILLER_40_283 ();
 FILLCELL_X1 FILLER_40_285 ();
 FILLCELL_X4 FILLER_40_291 ();
 FILLCELL_X1 FILLER_40_295 ();
 FILLCELL_X1 FILLER_40_300 ();
 FILLCELL_X2 FILLER_40_308 ();
 FILLCELL_X1 FILLER_40_314 ();
 FILLCELL_X1 FILLER_40_318 ();
 FILLCELL_X4 FILLER_40_338 ();
 FILLCELL_X2 FILLER_40_342 ();
 FILLCELL_X1 FILLER_40_344 ();
 FILLCELL_X4 FILLER_40_355 ();
 FILLCELL_X2 FILLER_40_359 ();
 FILLCELL_X8 FILLER_40_365 ();
 FILLCELL_X4 FILLER_40_373 ();
 FILLCELL_X1 FILLER_40_377 ();
 FILLCELL_X1 FILLER_40_381 ();
 FILLCELL_X8 FILLER_40_396 ();
 FILLCELL_X4 FILLER_40_404 ();
 FILLCELL_X2 FILLER_40_408 ();
 FILLCELL_X1 FILLER_40_410 ();
 FILLCELL_X2 FILLER_40_418 ();
 FILLCELL_X4 FILLER_40_424 ();
 FILLCELL_X1 FILLER_40_428 ();
 FILLCELL_X1 FILLER_40_431 ();
 FILLCELL_X1 FILLER_40_437 ();
 FILLCELL_X1 FILLER_40_448 ();
 FILLCELL_X4 FILLER_40_461 ();
 FILLCELL_X2 FILLER_40_465 ();
 FILLCELL_X1 FILLER_40_467 ();
 FILLCELL_X2 FILLER_40_484 ();
 FILLCELL_X1 FILLER_40_498 ();
 FILLCELL_X4 FILLER_40_503 ();
 FILLCELL_X2 FILLER_40_507 ();
 FILLCELL_X1 FILLER_40_509 ();
 FILLCELL_X4 FILLER_40_517 ();
 FILLCELL_X1 FILLER_40_521 ();
 FILLCELL_X4 FILLER_40_528 ();
 FILLCELL_X1 FILLER_40_532 ();
 FILLCELL_X8 FILLER_40_539 ();
 FILLCELL_X4 FILLER_40_547 ();
 FILLCELL_X2 FILLER_40_551 ();
 FILLCELL_X2 FILLER_40_557 ();
 FILLCELL_X1 FILLER_40_559 ();
 FILLCELL_X4 FILLER_40_586 ();
 FILLCELL_X1 FILLER_40_590 ();
 FILLCELL_X4 FILLER_40_615 ();
 FILLCELL_X1 FILLER_40_619 ();
 FILLCELL_X4 FILLER_40_627 ();
 FILLCELL_X4 FILLER_40_632 ();
 FILLCELL_X2 FILLER_40_636 ();
 FILLCELL_X2 FILLER_40_658 ();
 FILLCELL_X1 FILLER_40_660 ();
 FILLCELL_X16 FILLER_40_685 ();
 FILLCELL_X2 FILLER_40_701 ();
 FILLCELL_X1 FILLER_40_703 ();
 FILLCELL_X4 FILLER_40_733 ();
 FILLCELL_X2 FILLER_40_740 ();
 FILLCELL_X1 FILLER_40_755 ();
 FILLCELL_X1 FILLER_40_762 ();
 FILLCELL_X1 FILLER_40_767 ();
 FILLCELL_X16 FILLER_40_777 ();
 FILLCELL_X2 FILLER_40_793 ();
 FILLCELL_X8 FILLER_40_798 ();
 FILLCELL_X4 FILLER_40_806 ();
 FILLCELL_X1 FILLER_40_810 ();
 FILLCELL_X4 FILLER_40_831 ();
 FILLCELL_X1 FILLER_40_842 ();
 FILLCELL_X4 FILLER_40_874 ();
 FILLCELL_X1 FILLER_40_896 ();
 FILLCELL_X16 FILLER_40_915 ();
 FILLCELL_X8 FILLER_40_931 ();
 FILLCELL_X4 FILLER_40_939 ();
 FILLCELL_X2 FILLER_40_943 ();
 FILLCELL_X1 FILLER_40_945 ();
 FILLCELL_X2 FILLER_40_953 ();
 FILLCELL_X8 FILLER_40_975 ();
 FILLCELL_X16 FILLER_40_995 ();
 FILLCELL_X8 FILLER_40_1011 ();
 FILLCELL_X2 FILLER_40_1035 ();
 FILLCELL_X1 FILLER_40_1037 ();
 FILLCELL_X4 FILLER_40_1045 ();
 FILLCELL_X2 FILLER_40_1049 ();
 FILLCELL_X1 FILLER_40_1084 ();
 FILLCELL_X2 FILLER_40_1089 ();
 FILLCELL_X1 FILLER_40_1107 ();
 FILLCELL_X1 FILLER_40_1114 ();
 FILLCELL_X1 FILLER_40_1124 ();
 FILLCELL_X2 FILLER_40_1135 ();
 FILLCELL_X2 FILLER_40_1143 ();
 FILLCELL_X1 FILLER_40_1145 ();
 FILLCELL_X4 FILLER_40_1159 ();
 FILLCELL_X1 FILLER_40_1167 ();
 FILLCELL_X2 FILLER_40_1188 ();
 FILLCELL_X8 FILLER_40_1194 ();
 FILLCELL_X2 FILLER_40_1202 ();
 FILLCELL_X2 FILLER_40_1211 ();
 FILLCELL_X1 FILLER_40_1213 ();
 FILLCELL_X2 FILLER_40_1239 ();
 FILLCELL_X1 FILLER_40_1241 ();
 FILLCELL_X32 FILLER_40_1269 ();
 FILLCELL_X16 FILLER_40_1301 ();
 FILLCELL_X4 FILLER_40_1317 ();
 FILLCELL_X2 FILLER_40_1332 ();
 FILLCELL_X1 FILLER_40_1334 ();
 FILLCELL_X1 FILLER_40_1345 ();
 FILLCELL_X2 FILLER_40_1350 ();
 FILLCELL_X1 FILLER_40_1357 ();
 FILLCELL_X4 FILLER_40_1363 ();
 FILLCELL_X1 FILLER_40_1367 ();
 FILLCELL_X1 FILLER_40_1377 ();
 FILLCELL_X4 FILLER_40_1390 ();
 FILLCELL_X1 FILLER_40_1394 ();
 FILLCELL_X1 FILLER_40_1399 ();
 FILLCELL_X1 FILLER_40_1404 ();
 FILLCELL_X1 FILLER_40_1414 ();
 FILLCELL_X4 FILLER_40_1431 ();
 FILLCELL_X2 FILLER_40_1442 ();
 FILLCELL_X1 FILLER_40_1453 ();
 FILLCELL_X32 FILLER_40_1468 ();
 FILLCELL_X32 FILLER_40_1500 ();
 FILLCELL_X32 FILLER_40_1532 ();
 FILLCELL_X32 FILLER_40_1564 ();
 FILLCELL_X32 FILLER_40_1596 ();
 FILLCELL_X16 FILLER_40_1628 ();
 FILLCELL_X4 FILLER_40_1644 ();
 FILLCELL_X2 FILLER_40_1648 ();
 FILLCELL_X1 FILLER_40_1650 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X8 FILLER_41_193 ();
 FILLCELL_X4 FILLER_41_201 ();
 FILLCELL_X8 FILLER_41_239 ();
 FILLCELL_X1 FILLER_41_247 ();
 FILLCELL_X1 FILLER_41_285 ();
 FILLCELL_X2 FILLER_41_289 ();
 FILLCELL_X1 FILLER_41_311 ();
 FILLCELL_X2 FILLER_41_315 ();
 FILLCELL_X2 FILLER_41_320 ();
 FILLCELL_X1 FILLER_41_327 ();
 FILLCELL_X1 FILLER_41_333 ();
 FILLCELL_X4 FILLER_41_393 ();
 FILLCELL_X2 FILLER_41_397 ();
 FILLCELL_X1 FILLER_41_399 ();
 FILLCELL_X2 FILLER_41_423 ();
 FILLCELL_X1 FILLER_41_425 ();
 FILLCELL_X16 FILLER_41_447 ();
 FILLCELL_X8 FILLER_41_463 ();
 FILLCELL_X4 FILLER_41_471 ();
 FILLCELL_X2 FILLER_41_475 ();
 FILLCELL_X8 FILLER_41_480 ();
 FILLCELL_X1 FILLER_41_488 ();
 FILLCELL_X4 FILLER_41_507 ();
 FILLCELL_X4 FILLER_41_516 ();
 FILLCELL_X1 FILLER_41_520 ();
 FILLCELL_X4 FILLER_41_587 ();
 FILLCELL_X1 FILLER_41_591 ();
 FILLCELL_X8 FILLER_41_599 ();
 FILLCELL_X1 FILLER_41_607 ();
 FILLCELL_X4 FILLER_41_615 ();
 FILLCELL_X2 FILLER_41_619 ();
 FILLCELL_X1 FILLER_41_642 ();
 FILLCELL_X4 FILLER_41_650 ();
 FILLCELL_X2 FILLER_41_654 ();
 FILLCELL_X1 FILLER_41_656 ();
 FILLCELL_X8 FILLER_41_661 ();
 FILLCELL_X2 FILLER_41_669 ();
 FILLCELL_X1 FILLER_41_671 ();
 FILLCELL_X1 FILLER_41_677 ();
 FILLCELL_X32 FILLER_41_710 ();
 FILLCELL_X4 FILLER_41_742 ();
 FILLCELL_X2 FILLER_41_755 ();
 FILLCELL_X2 FILLER_41_760 ();
 FILLCELL_X1 FILLER_41_762 ();
 FILLCELL_X4 FILLER_41_768 ();
 FILLCELL_X1 FILLER_41_772 ();
 FILLCELL_X1 FILLER_41_787 ();
 FILLCELL_X4 FILLER_41_799 ();
 FILLCELL_X1 FILLER_41_803 ();
 FILLCELL_X8 FILLER_41_829 ();
 FILLCELL_X2 FILLER_41_837 ();
 FILLCELL_X1 FILLER_41_839 ();
 FILLCELL_X2 FILLER_41_871 ();
 FILLCELL_X1 FILLER_41_873 ();
 FILLCELL_X2 FILLER_41_921 ();
 FILLCELL_X1 FILLER_41_923 ();
 FILLCELL_X4 FILLER_41_965 ();
 FILLCELL_X2 FILLER_41_969 ();
 FILLCELL_X1 FILLER_41_971 ();
 FILLCELL_X4 FILLER_41_992 ();
 FILLCELL_X2 FILLER_41_996 ();
 FILLCELL_X1 FILLER_41_998 ();
 FILLCELL_X16 FILLER_41_1050 ();
 FILLCELL_X8 FILLER_41_1066 ();
 FILLCELL_X4 FILLER_41_1074 ();
 FILLCELL_X1 FILLER_41_1078 ();
 FILLCELL_X2 FILLER_41_1096 ();
 FILLCELL_X1 FILLER_41_1098 ();
 FILLCELL_X2 FILLER_41_1123 ();
 FILLCELL_X1 FILLER_41_1125 ();
 FILLCELL_X8 FILLER_41_1153 ();
 FILLCELL_X2 FILLER_41_1161 ();
 FILLCELL_X1 FILLER_41_1169 ();
 FILLCELL_X8 FILLER_41_1178 ();
 FILLCELL_X4 FILLER_41_1186 ();
 FILLCELL_X2 FILLER_41_1190 ();
 FILLCELL_X4 FILLER_41_1259 ();
 FILLCELL_X16 FILLER_41_1291 ();
 FILLCELL_X8 FILLER_41_1307 ();
 FILLCELL_X4 FILLER_41_1315 ();
 FILLCELL_X4 FILLER_41_1328 ();
 FILLCELL_X1 FILLER_41_1332 ();
 FILLCELL_X1 FILLER_41_1338 ();
 FILLCELL_X4 FILLER_41_1353 ();
 FILLCELL_X1 FILLER_41_1357 ();
 FILLCELL_X1 FILLER_41_1361 ();
 FILLCELL_X2 FILLER_41_1392 ();
 FILLCELL_X1 FILLER_41_1394 ();
 FILLCELL_X1 FILLER_41_1406 ();
 FILLCELL_X1 FILLER_41_1418 ();
 FILLCELL_X4 FILLER_41_1428 ();
 FILLCELL_X2 FILLER_41_1432 ();
 FILLCELL_X32 FILLER_41_1441 ();
 FILLCELL_X32 FILLER_41_1473 ();
 FILLCELL_X32 FILLER_41_1505 ();
 FILLCELL_X32 FILLER_41_1537 ();
 FILLCELL_X32 FILLER_41_1569 ();
 FILLCELL_X32 FILLER_41_1601 ();
 FILLCELL_X16 FILLER_41_1633 ();
 FILLCELL_X2 FILLER_41_1649 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X4 FILLER_42_225 ();
 FILLCELL_X2 FILLER_42_229 ();
 FILLCELL_X2 FILLER_42_262 ();
 FILLCELL_X16 FILLER_42_288 ();
 FILLCELL_X8 FILLER_42_304 ();
 FILLCELL_X2 FILLER_42_312 ();
 FILLCELL_X4 FILLER_42_330 ();
 FILLCELL_X2 FILLER_42_334 ();
 FILLCELL_X1 FILLER_42_336 ();
 FILLCELL_X4 FILLER_42_344 ();
 FILLCELL_X2 FILLER_42_348 ();
 FILLCELL_X1 FILLER_42_350 ();
 FILLCELL_X2 FILLER_42_354 ();
 FILLCELL_X1 FILLER_42_356 ();
 FILLCELL_X16 FILLER_42_389 ();
 FILLCELL_X1 FILLER_42_408 ();
 FILLCELL_X1 FILLER_42_426 ();
 FILLCELL_X1 FILLER_42_436 ();
 FILLCELL_X1 FILLER_42_441 ();
 FILLCELL_X16 FILLER_42_455 ();
 FILLCELL_X4 FILLER_42_475 ();
 FILLCELL_X4 FILLER_42_488 ();
 FILLCELL_X2 FILLER_42_492 ();
 FILLCELL_X8 FILLER_42_499 ();
 FILLCELL_X4 FILLER_42_507 ();
 FILLCELL_X2 FILLER_42_511 ();
 FILLCELL_X1 FILLER_42_513 ();
 FILLCELL_X4 FILLER_42_527 ();
 FILLCELL_X8 FILLER_42_538 ();
 FILLCELL_X2 FILLER_42_546 ();
 FILLCELL_X4 FILLER_42_586 ();
 FILLCELL_X2 FILLER_42_590 ();
 FILLCELL_X1 FILLER_42_592 ();
 FILLCELL_X8 FILLER_42_607 ();
 FILLCELL_X4 FILLER_42_615 ();
 FILLCELL_X4 FILLER_42_626 ();
 FILLCELL_X1 FILLER_42_630 ();
 FILLCELL_X8 FILLER_42_632 ();
 FILLCELL_X1 FILLER_42_640 ();
 FILLCELL_X4 FILLER_42_662 ();
 FILLCELL_X2 FILLER_42_714 ();
 FILLCELL_X1 FILLER_42_716 ();
 FILLCELL_X1 FILLER_42_721 ();
 FILLCELL_X8 FILLER_42_742 ();
 FILLCELL_X1 FILLER_42_750 ();
 FILLCELL_X4 FILLER_42_772 ();
 FILLCELL_X16 FILLER_42_814 ();
 FILLCELL_X8 FILLER_42_830 ();
 FILLCELL_X2 FILLER_42_843 ();
 FILLCELL_X1 FILLER_42_845 ();
 FILLCELL_X4 FILLER_42_852 ();
 FILLCELL_X1 FILLER_42_856 ();
 FILLCELL_X1 FILLER_42_926 ();
 FILLCELL_X8 FILLER_42_932 ();
 FILLCELL_X1 FILLER_42_940 ();
 FILLCELL_X2 FILLER_42_951 ();
 FILLCELL_X1 FILLER_42_961 ();
 FILLCELL_X2 FILLER_42_964 ();
 FILLCELL_X2 FILLER_42_1007 ();
 FILLCELL_X2 FILLER_42_1014 ();
 FILLCELL_X1 FILLER_42_1016 ();
 FILLCELL_X2 FILLER_42_1030 ();
 FILLCELL_X2 FILLER_42_1035 ();
 FILLCELL_X2 FILLER_42_1093 ();
 FILLCELL_X1 FILLER_42_1095 ();
 FILLCELL_X1 FILLER_42_1108 ();
 FILLCELL_X4 FILLER_42_1113 ();
 FILLCELL_X2 FILLER_42_1117 ();
 FILLCELL_X2 FILLER_42_1137 ();
 FILLCELL_X1 FILLER_42_1161 ();
 FILLCELL_X1 FILLER_42_1184 ();
 FILLCELL_X1 FILLER_42_1190 ();
 FILLCELL_X16 FILLER_42_1223 ();
 FILLCELL_X8 FILLER_42_1239 ();
 FILLCELL_X2 FILLER_42_1247 ();
 FILLCELL_X1 FILLER_42_1249 ();
 FILLCELL_X4 FILLER_42_1257 ();
 FILLCELL_X2 FILLER_42_1261 ();
 FILLCELL_X1 FILLER_42_1271 ();
 FILLCELL_X16 FILLER_42_1312 ();
 FILLCELL_X8 FILLER_42_1328 ();
 FILLCELL_X1 FILLER_42_1336 ();
 FILLCELL_X1 FILLER_42_1372 ();
 FILLCELL_X2 FILLER_42_1377 ();
 FILLCELL_X1 FILLER_42_1379 ();
 FILLCELL_X1 FILLER_42_1389 ();
 FILLCELL_X1 FILLER_42_1397 ();
 FILLCELL_X2 FILLER_42_1407 ();
 FILLCELL_X2 FILLER_42_1431 ();
 FILLCELL_X1 FILLER_42_1433 ();
 FILLCELL_X32 FILLER_42_1450 ();
 FILLCELL_X8 FILLER_42_1482 ();
 FILLCELL_X4 FILLER_42_1490 ();
 FILLCELL_X1 FILLER_42_1494 ();
 FILLCELL_X32 FILLER_42_1502 ();
 FILLCELL_X32 FILLER_42_1534 ();
 FILLCELL_X32 FILLER_42_1566 ();
 FILLCELL_X32 FILLER_42_1598 ();
 FILLCELL_X16 FILLER_42_1630 ();
 FILLCELL_X4 FILLER_42_1646 ();
 FILLCELL_X1 FILLER_42_1650 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X8 FILLER_43_193 ();
 FILLCELL_X2 FILLER_43_201 ();
 FILLCELL_X8 FILLER_43_226 ();
 FILLCELL_X4 FILLER_43_234 ();
 FILLCELL_X2 FILLER_43_238 ();
 FILLCELL_X1 FILLER_43_240 ();
 FILLCELL_X16 FILLER_43_248 ();
 FILLCELL_X4 FILLER_43_264 ();
 FILLCELL_X2 FILLER_43_268 ();
 FILLCELL_X4 FILLER_43_274 ();
 FILLCELL_X2 FILLER_43_278 ();
 FILLCELL_X1 FILLER_43_280 ();
 FILLCELL_X2 FILLER_43_305 ();
 FILLCELL_X1 FILLER_43_307 ();
 FILLCELL_X4 FILLER_43_324 ();
 FILLCELL_X2 FILLER_43_362 ();
 FILLCELL_X1 FILLER_43_364 ();
 FILLCELL_X2 FILLER_43_394 ();
 FILLCELL_X1 FILLER_43_396 ();
 FILLCELL_X4 FILLER_43_434 ();
 FILLCELL_X8 FILLER_43_458 ();
 FILLCELL_X1 FILLER_43_466 ();
 FILLCELL_X1 FILLER_43_471 ();
 FILLCELL_X1 FILLER_43_474 ();
 FILLCELL_X1 FILLER_43_490 ();
 FILLCELL_X2 FILLER_43_510 ();
 FILLCELL_X1 FILLER_43_519 ();
 FILLCELL_X1 FILLER_43_526 ();
 FILLCELL_X1 FILLER_43_534 ();
 FILLCELL_X2 FILLER_43_540 ();
 FILLCELL_X1 FILLER_43_542 ();
 FILLCELL_X4 FILLER_43_559 ();
 FILLCELL_X8 FILLER_43_568 ();
 FILLCELL_X4 FILLER_43_582 ();
 FILLCELL_X2 FILLER_43_586 ();
 FILLCELL_X1 FILLER_43_588 ();
 FILLCELL_X8 FILLER_43_596 ();
 FILLCELL_X1 FILLER_43_604 ();
 FILLCELL_X8 FILLER_43_625 ();
 FILLCELL_X2 FILLER_43_633 ();
 FILLCELL_X4 FILLER_43_697 ();
 FILLCELL_X1 FILLER_43_701 ();
 FILLCELL_X16 FILLER_43_757 ();
 FILLCELL_X1 FILLER_43_795 ();
 FILLCELL_X1 FILLER_43_809 ();
 FILLCELL_X4 FILLER_43_813 ();
 FILLCELL_X1 FILLER_43_817 ();
 FILLCELL_X4 FILLER_43_825 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X4 FILLER_43_879 ();
 FILLCELL_X8 FILLER_43_901 ();
 FILLCELL_X2 FILLER_43_909 ();
 FILLCELL_X1 FILLER_43_911 ();
 FILLCELL_X4 FILLER_43_917 ();
 FILLCELL_X2 FILLER_43_921 ();
 FILLCELL_X4 FILLER_43_930 ();
 FILLCELL_X2 FILLER_43_934 ();
 FILLCELL_X8 FILLER_43_975 ();
 FILLCELL_X2 FILLER_43_1003 ();
 FILLCELL_X1 FILLER_43_1052 ();
 FILLCELL_X1 FILLER_43_1064 ();
 FILLCELL_X1 FILLER_43_1080 ();
 FILLCELL_X4 FILLER_43_1094 ();
 FILLCELL_X2 FILLER_43_1098 ();
 FILLCELL_X1 FILLER_43_1100 ();
 FILLCELL_X8 FILLER_43_1112 ();
 FILLCELL_X4 FILLER_43_1124 ();
 FILLCELL_X2 FILLER_43_1128 ();
 FILLCELL_X1 FILLER_43_1130 ();
 FILLCELL_X2 FILLER_43_1160 ();
 FILLCELL_X2 FILLER_43_1168 ();
 FILLCELL_X1 FILLER_43_1170 ();
 FILLCELL_X2 FILLER_43_1175 ();
 FILLCELL_X1 FILLER_43_1177 ();
 FILLCELL_X4 FILLER_43_1198 ();
 FILLCELL_X2 FILLER_43_1208 ();
 FILLCELL_X16 FILLER_43_1214 ();
 FILLCELL_X8 FILLER_43_1230 ();
 FILLCELL_X4 FILLER_43_1238 ();
 FILLCELL_X1 FILLER_43_1242 ();
 FILLCELL_X2 FILLER_43_1271 ();
 FILLCELL_X8 FILLER_43_1300 ();
 FILLCELL_X2 FILLER_43_1308 ();
 FILLCELL_X1 FILLER_43_1310 ();
 FILLCELL_X16 FILLER_43_1318 ();
 FILLCELL_X2 FILLER_43_1334 ();
 FILLCELL_X4 FILLER_43_1367 ();
 FILLCELL_X2 FILLER_43_1375 ();
 FILLCELL_X2 FILLER_43_1400 ();
 FILLCELL_X2 FILLER_43_1427 ();
 FILLCELL_X16 FILLER_43_1438 ();
 FILLCELL_X8 FILLER_43_1454 ();
 FILLCELL_X2 FILLER_43_1462 ();
 FILLCELL_X4 FILLER_43_1478 ();
 FILLCELL_X2 FILLER_43_1482 ();
 FILLCELL_X1 FILLER_43_1484 ();
 FILLCELL_X1 FILLER_43_1503 ();
 FILLCELL_X2 FILLER_43_1525 ();
 FILLCELL_X4 FILLER_43_1544 ();
 FILLCELL_X2 FILLER_43_1548 ();
 FILLCELL_X8 FILLER_43_1557 ();
 FILLCELL_X32 FILLER_43_1569 ();
 FILLCELL_X32 FILLER_43_1601 ();
 FILLCELL_X16 FILLER_43_1633 ();
 FILLCELL_X2 FILLER_43_1649 ();
 FILLCELL_X16 FILLER_44_1 ();
 FILLCELL_X4 FILLER_44_17 ();
 FILLCELL_X1 FILLER_44_21 ();
 FILLCELL_X32 FILLER_44_26 ();
 FILLCELL_X32 FILLER_44_58 ();
 FILLCELL_X32 FILLER_44_90 ();
 FILLCELL_X32 FILLER_44_122 ();
 FILLCELL_X32 FILLER_44_154 ();
 FILLCELL_X16 FILLER_44_186 ();
 FILLCELL_X8 FILLER_44_202 ();
 FILLCELL_X4 FILLER_44_210 ();
 FILLCELL_X2 FILLER_44_214 ();
 FILLCELL_X4 FILLER_44_242 ();
 FILLCELL_X2 FILLER_44_277 ();
 FILLCELL_X1 FILLER_44_279 ();
 FILLCELL_X1 FILLER_44_286 ();
 FILLCELL_X4 FILLER_44_294 ();
 FILLCELL_X2 FILLER_44_298 ();
 FILLCELL_X2 FILLER_44_361 ();
 FILLCELL_X2 FILLER_44_367 ();
 FILLCELL_X4 FILLER_44_375 ();
 FILLCELL_X1 FILLER_44_386 ();
 FILLCELL_X2 FILLER_44_405 ();
 FILLCELL_X1 FILLER_44_407 ();
 FILLCELL_X16 FILLER_44_418 ();
 FILLCELL_X2 FILLER_44_434 ();
 FILLCELL_X1 FILLER_44_436 ();
 FILLCELL_X2 FILLER_44_444 ();
 FILLCELL_X1 FILLER_44_446 ();
 FILLCELL_X2 FILLER_44_452 ();
 FILLCELL_X1 FILLER_44_454 ();
 FILLCELL_X8 FILLER_44_465 ();
 FILLCELL_X2 FILLER_44_473 ();
 FILLCELL_X1 FILLER_44_475 ();
 FILLCELL_X1 FILLER_44_480 ();
 FILLCELL_X4 FILLER_44_488 ();
 FILLCELL_X1 FILLER_44_492 ();
 FILLCELL_X4 FILLER_44_497 ();
 FILLCELL_X2 FILLER_44_501 ();
 FILLCELL_X2 FILLER_44_563 ();
 FILLCELL_X1 FILLER_44_565 ();
 FILLCELL_X8 FILLER_44_576 ();
 FILLCELL_X4 FILLER_44_584 ();
 FILLCELL_X1 FILLER_44_588 ();
 FILLCELL_X1 FILLER_44_616 ();
 FILLCELL_X2 FILLER_44_663 ();
 FILLCELL_X1 FILLER_44_665 ();
 FILLCELL_X2 FILLER_44_691 ();
 FILLCELL_X4 FILLER_44_695 ();
 FILLCELL_X2 FILLER_44_699 ();
 FILLCELL_X1 FILLER_44_701 ();
 FILLCELL_X2 FILLER_44_716 ();
 FILLCELL_X8 FILLER_44_729 ();
 FILLCELL_X1 FILLER_44_775 ();
 FILLCELL_X4 FILLER_44_797 ();
 FILLCELL_X4 FILLER_44_808 ();
 FILLCELL_X1 FILLER_44_812 ();
 FILLCELL_X4 FILLER_44_838 ();
 FILLCELL_X8 FILLER_44_862 ();
 FILLCELL_X8 FILLER_44_877 ();
 FILLCELL_X8 FILLER_44_891 ();
 FILLCELL_X2 FILLER_44_915 ();
 FILLCELL_X1 FILLER_44_934 ();
 FILLCELL_X2 FILLER_44_976 ();
 FILLCELL_X1 FILLER_44_978 ();
 FILLCELL_X1 FILLER_44_997 ();
 FILLCELL_X1 FILLER_44_1003 ();
 FILLCELL_X1 FILLER_44_1010 ();
 FILLCELL_X16 FILLER_44_1013 ();
 FILLCELL_X1 FILLER_44_1031 ();
 FILLCELL_X8 FILLER_44_1035 ();
 FILLCELL_X8 FILLER_44_1067 ();
 FILLCELL_X4 FILLER_44_1075 ();
 FILLCELL_X2 FILLER_44_1079 ();
 FILLCELL_X2 FILLER_44_1109 ();
 FILLCELL_X4 FILLER_44_1113 ();
 FILLCELL_X2 FILLER_44_1117 ();
 FILLCELL_X1 FILLER_44_1119 ();
 FILLCELL_X1 FILLER_44_1144 ();
 FILLCELL_X4 FILLER_44_1149 ();
 FILLCELL_X2 FILLER_44_1153 ();
 FILLCELL_X1 FILLER_44_1155 ();
 FILLCELL_X1 FILLER_44_1164 ();
 FILLCELL_X1 FILLER_44_1169 ();
 FILLCELL_X16 FILLER_44_1172 ();
 FILLCELL_X8 FILLER_44_1188 ();
 FILLCELL_X2 FILLER_44_1196 ();
 FILLCELL_X2 FILLER_44_1202 ();
 FILLCELL_X1 FILLER_44_1204 ();
 FILLCELL_X8 FILLER_44_1230 ();
 FILLCELL_X4 FILLER_44_1279 ();
 FILLCELL_X1 FILLER_44_1283 ();
 FILLCELL_X1 FILLER_44_1298 ();
 FILLCELL_X16 FILLER_44_1319 ();
 FILLCELL_X2 FILLER_44_1335 ();
 FILLCELL_X8 FILLER_44_1360 ();
 FILLCELL_X4 FILLER_44_1368 ();
 FILLCELL_X8 FILLER_44_1404 ();
 FILLCELL_X1 FILLER_44_1412 ();
 FILLCELL_X16 FILLER_44_1427 ();
 FILLCELL_X4 FILLER_44_1443 ();
 FILLCELL_X8 FILLER_44_1456 ();
 FILLCELL_X1 FILLER_44_1464 ();
 FILLCELL_X8 FILLER_44_1474 ();
 FILLCELL_X1 FILLER_44_1482 ();
 FILLCELL_X4 FILLER_44_1490 ();
 FILLCELL_X2 FILLER_44_1494 ();
 FILLCELL_X4 FILLER_44_1498 ();
 FILLCELL_X2 FILLER_44_1502 ();
 FILLCELL_X1 FILLER_44_1504 ();
 FILLCELL_X32 FILLER_44_1509 ();
 FILLCELL_X2 FILLER_44_1541 ();
 FILLCELL_X1 FILLER_44_1543 ();
 FILLCELL_X2 FILLER_44_1570 ();
 FILLCELL_X1 FILLER_44_1575 ();
 FILLCELL_X8 FILLER_44_1583 ();
 FILLCELL_X32 FILLER_44_1598 ();
 FILLCELL_X16 FILLER_44_1630 ();
 FILLCELL_X4 FILLER_44_1646 ();
 FILLCELL_X1 FILLER_44_1650 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X1 FILLER_45_193 ();
 FILLCELL_X1 FILLER_45_223 ();
 FILLCELL_X4 FILLER_45_231 ();
 FILLCELL_X1 FILLER_45_235 ();
 FILLCELL_X2 FILLER_45_243 ();
 FILLCELL_X1 FILLER_45_245 ();
 FILLCELL_X2 FILLER_45_258 ();
 FILLCELL_X2 FILLER_45_263 ();
 FILLCELL_X4 FILLER_45_281 ();
 FILLCELL_X1 FILLER_45_285 ();
 FILLCELL_X1 FILLER_45_320 ();
 FILLCELL_X16 FILLER_45_339 ();
 FILLCELL_X4 FILLER_45_355 ();
 FILLCELL_X1 FILLER_45_359 ();
 FILLCELL_X8 FILLER_45_363 ();
 FILLCELL_X4 FILLER_45_371 ();
 FILLCELL_X2 FILLER_45_375 ();
 FILLCELL_X1 FILLER_45_377 ();
 FILLCELL_X2 FILLER_45_382 ();
 FILLCELL_X16 FILLER_45_390 ();
 FILLCELL_X1 FILLER_45_406 ();
 FILLCELL_X4 FILLER_45_414 ();
 FILLCELL_X2 FILLER_45_418 ();
 FILLCELL_X2 FILLER_45_434 ();
 FILLCELL_X1 FILLER_45_445 ();
 FILLCELL_X1 FILLER_45_453 ();
 FILLCELL_X1 FILLER_45_498 ();
 FILLCELL_X1 FILLER_45_504 ();
 FILLCELL_X1 FILLER_45_515 ();
 FILLCELL_X2 FILLER_45_521 ();
 FILLCELL_X1 FILLER_45_523 ();
 FILLCELL_X2 FILLER_45_529 ();
 FILLCELL_X1 FILLER_45_571 ();
 FILLCELL_X1 FILLER_45_586 ();
 FILLCELL_X8 FILLER_45_593 ();
 FILLCELL_X2 FILLER_45_601 ();
 FILLCELL_X1 FILLER_45_603 ();
 FILLCELL_X1 FILLER_45_625 ();
 FILLCELL_X4 FILLER_45_644 ();
 FILLCELL_X2 FILLER_45_648 ();
 FILLCELL_X1 FILLER_45_650 ();
 FILLCELL_X4 FILLER_45_658 ();
 FILLCELL_X1 FILLER_45_662 ();
 FILLCELL_X4 FILLER_45_674 ();
 FILLCELL_X2 FILLER_45_678 ();
 FILLCELL_X1 FILLER_45_680 ();
 FILLCELL_X1 FILLER_45_691 ();
 FILLCELL_X4 FILLER_45_709 ();
 FILLCELL_X2 FILLER_45_713 ();
 FILLCELL_X8 FILLER_45_720 ();
 FILLCELL_X2 FILLER_45_738 ();
 FILLCELL_X1 FILLER_45_752 ();
 FILLCELL_X4 FILLER_45_756 ();
 FILLCELL_X1 FILLER_45_760 ();
 FILLCELL_X4 FILLER_45_771 ();
 FILLCELL_X1 FILLER_45_775 ();
 FILLCELL_X1 FILLER_45_786 ();
 FILLCELL_X1 FILLER_45_807 ();
 FILLCELL_X8 FILLER_45_813 ();
 FILLCELL_X1 FILLER_45_821 ();
 FILLCELL_X4 FILLER_45_853 ();
 FILLCELL_X2 FILLER_45_857 ();
 FILLCELL_X1 FILLER_45_868 ();
 FILLCELL_X16 FILLER_45_874 ();
 FILLCELL_X16 FILLER_45_894 ();
 FILLCELL_X2 FILLER_45_910 ();
 FILLCELL_X8 FILLER_45_915 ();
 FILLCELL_X1 FILLER_45_923 ();
 FILLCELL_X8 FILLER_45_930 ();
 FILLCELL_X4 FILLER_45_938 ();
 FILLCELL_X1 FILLER_45_942 ();
 FILLCELL_X4 FILLER_45_955 ();
 FILLCELL_X1 FILLER_45_959 ();
 FILLCELL_X4 FILLER_45_985 ();
 FILLCELL_X2 FILLER_45_989 ();
 FILLCELL_X4 FILLER_45_1011 ();
 FILLCELL_X1 FILLER_45_1015 ();
 FILLCELL_X2 FILLER_45_1023 ();
 FILLCELL_X1 FILLER_45_1025 ();
 FILLCELL_X4 FILLER_45_1044 ();
 FILLCELL_X2 FILLER_45_1048 ();
 FILLCELL_X8 FILLER_45_1072 ();
 FILLCELL_X1 FILLER_45_1080 ();
 FILLCELL_X1 FILLER_45_1129 ();
 FILLCELL_X4 FILLER_45_1137 ();
 FILLCELL_X2 FILLER_45_1150 ();
 FILLCELL_X1 FILLER_45_1152 ();
 FILLCELL_X2 FILLER_45_1181 ();
 FILLCELL_X1 FILLER_45_1203 ();
 FILLCELL_X8 FILLER_45_1208 ();
 FILLCELL_X2 FILLER_45_1216 ();
 FILLCELL_X4 FILLER_45_1258 ();
 FILLCELL_X1 FILLER_45_1262 ();
 FILLCELL_X8 FILLER_45_1264 ();
 FILLCELL_X2 FILLER_45_1272 ();
 FILLCELL_X2 FILLER_45_1306 ();
 FILLCELL_X32 FILLER_45_1315 ();
 FILLCELL_X2 FILLER_45_1347 ();
 FILLCELL_X2 FILLER_45_1356 ();
 FILLCELL_X1 FILLER_45_1358 ();
 FILLCELL_X32 FILLER_45_1406 ();
 FILLCELL_X8 FILLER_45_1438 ();
 FILLCELL_X2 FILLER_45_1446 ();
 FILLCELL_X2 FILLER_45_1471 ();
 FILLCELL_X4 FILLER_45_1489 ();
 FILLCELL_X4 FILLER_45_1514 ();
 FILLCELL_X2 FILLER_45_1518 ();
 FILLCELL_X2 FILLER_45_1528 ();
 FILLCELL_X1 FILLER_45_1530 ();
 FILLCELL_X2 FILLER_45_1547 ();
 FILLCELL_X8 FILLER_45_1562 ();
 FILLCELL_X2 FILLER_45_1570 ();
 FILLCELL_X1 FILLER_45_1572 ();
 FILLCELL_X4 FILLER_45_1577 ();
 FILLCELL_X1 FILLER_45_1585 ();
 FILLCELL_X8 FILLER_45_1589 ();
 FILLCELL_X8 FILLER_45_1601 ();
 FILLCELL_X4 FILLER_45_1609 ();
 FILLCELL_X1 FILLER_45_1613 ();
 FILLCELL_X16 FILLER_45_1621 ();
 FILLCELL_X8 FILLER_45_1637 ();
 FILLCELL_X4 FILLER_45_1645 ();
 FILLCELL_X2 FILLER_45_1649 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X16 FILLER_46_161 ();
 FILLCELL_X8 FILLER_46_177 ();
 FILLCELL_X4 FILLER_46_185 ();
 FILLCELL_X2 FILLER_46_189 ();
 FILLCELL_X1 FILLER_46_191 ();
 FILLCELL_X4 FILLER_46_253 ();
 FILLCELL_X2 FILLER_46_257 ();
 FILLCELL_X8 FILLER_46_263 ();
 FILLCELL_X8 FILLER_46_346 ();
 FILLCELL_X4 FILLER_46_354 ();
 FILLCELL_X1 FILLER_46_358 ();
 FILLCELL_X2 FILLER_46_379 ();
 FILLCELL_X1 FILLER_46_381 ();
 FILLCELL_X2 FILLER_46_443 ();
 FILLCELL_X16 FILLER_46_465 ();
 FILLCELL_X2 FILLER_46_481 ();
 FILLCELL_X1 FILLER_46_488 ();
 FILLCELL_X1 FILLER_46_492 ();
 FILLCELL_X16 FILLER_46_505 ();
 FILLCELL_X2 FILLER_46_535 ();
 FILLCELL_X1 FILLER_46_537 ();
 FILLCELL_X4 FILLER_46_560 ();
 FILLCELL_X2 FILLER_46_564 ();
 FILLCELL_X1 FILLER_46_570 ();
 FILLCELL_X1 FILLER_46_585 ();
 FILLCELL_X4 FILLER_46_595 ();
 FILLCELL_X2 FILLER_46_599 ();
 FILLCELL_X4 FILLER_46_610 ();
 FILLCELL_X1 FILLER_46_614 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X2 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_641 ();
 FILLCELL_X4 FILLER_46_673 ();
 FILLCELL_X2 FILLER_46_677 ();
 FILLCELL_X2 FILLER_46_685 ();
 FILLCELL_X1 FILLER_46_687 ();
 FILLCELL_X2 FILLER_46_708 ();
 FILLCELL_X1 FILLER_46_710 ();
 FILLCELL_X1 FILLER_46_715 ();
 FILLCELL_X2 FILLER_46_723 ();
 FILLCELL_X1 FILLER_46_727 ();
 FILLCELL_X2 FILLER_46_731 ();
 FILLCELL_X16 FILLER_46_753 ();
 FILLCELL_X4 FILLER_46_769 ();
 FILLCELL_X1 FILLER_46_773 ();
 FILLCELL_X1 FILLER_46_797 ();
 FILLCELL_X1 FILLER_46_834 ();
 FILLCELL_X2 FILLER_46_840 ();
 FILLCELL_X32 FILLER_46_850 ();
 FILLCELL_X8 FILLER_46_882 ();
 FILLCELL_X2 FILLER_46_890 ();
 FILLCELL_X4 FILLER_46_899 ();
 FILLCELL_X2 FILLER_46_903 ();
 FILLCELL_X1 FILLER_46_905 ();
 FILLCELL_X4 FILLER_46_921 ();
 FILLCELL_X1 FILLER_46_925 ();
 FILLCELL_X1 FILLER_46_942 ();
 FILLCELL_X2 FILLER_46_958 ();
 FILLCELL_X2 FILLER_46_965 ();
 FILLCELL_X1 FILLER_46_967 ();
 FILLCELL_X8 FILLER_46_977 ();
 FILLCELL_X1 FILLER_46_985 ();
 FILLCELL_X4 FILLER_46_996 ();
 FILLCELL_X2 FILLER_46_1000 ();
 FILLCELL_X4 FILLER_46_1053 ();
 FILLCELL_X8 FILLER_46_1073 ();
 FILLCELL_X1 FILLER_46_1081 ();
 FILLCELL_X1 FILLER_46_1091 ();
 FILLCELL_X8 FILLER_46_1106 ();
 FILLCELL_X2 FILLER_46_1114 ();
 FILLCELL_X1 FILLER_46_1130 ();
 FILLCELL_X2 FILLER_46_1137 ();
 FILLCELL_X1 FILLER_46_1139 ();
 FILLCELL_X2 FILLER_46_1146 ();
 FILLCELL_X1 FILLER_46_1148 ();
 FILLCELL_X8 FILLER_46_1163 ();
 FILLCELL_X1 FILLER_46_1173 ();
 FILLCELL_X2 FILLER_46_1178 ();
 FILLCELL_X1 FILLER_46_1180 ();
 FILLCELL_X2 FILLER_46_1197 ();
 FILLCELL_X2 FILLER_46_1209 ();
 FILLCELL_X8 FILLER_46_1225 ();
 FILLCELL_X2 FILLER_46_1260 ();
 FILLCELL_X1 FILLER_46_1292 ();
 FILLCELL_X4 FILLER_46_1306 ();
 FILLCELL_X2 FILLER_46_1343 ();
 FILLCELL_X4 FILLER_46_1365 ();
 FILLCELL_X1 FILLER_46_1369 ();
 FILLCELL_X2 FILLER_46_1377 ();
 FILLCELL_X1 FILLER_46_1388 ();
 FILLCELL_X2 FILLER_46_1398 ();
 FILLCELL_X1 FILLER_46_1400 ();
 FILLCELL_X1 FILLER_46_1422 ();
 FILLCELL_X4 FILLER_46_1437 ();
 FILLCELL_X4 FILLER_46_1450 ();
 FILLCELL_X2 FILLER_46_1470 ();
 FILLCELL_X1 FILLER_46_1472 ();
 FILLCELL_X1 FILLER_46_1477 ();
 FILLCELL_X8 FILLER_46_1506 ();
 FILLCELL_X1 FILLER_46_1514 ();
 FILLCELL_X16 FILLER_46_1527 ();
 FILLCELL_X2 FILLER_46_1543 ();
 FILLCELL_X1 FILLER_46_1545 ();
 FILLCELL_X4 FILLER_46_1559 ();
 FILLCELL_X8 FILLER_46_1568 ();
 FILLCELL_X4 FILLER_46_1583 ();
 FILLCELL_X4 FILLER_46_1591 ();
 FILLCELL_X1 FILLER_46_1595 ();
 FILLCELL_X32 FILLER_46_1607 ();
 FILLCELL_X8 FILLER_46_1639 ();
 FILLCELL_X4 FILLER_46_1647 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X2 FILLER_47_193 ();
 FILLCELL_X2 FILLER_47_208 ();
 FILLCELL_X16 FILLER_47_219 ();
 FILLCELL_X1 FILLER_47_235 ();
 FILLCELL_X4 FILLER_47_243 ();
 FILLCELL_X2 FILLER_47_251 ();
 FILLCELL_X1 FILLER_47_253 ();
 FILLCELL_X1 FILLER_47_263 ();
 FILLCELL_X2 FILLER_47_266 ();
 FILLCELL_X1 FILLER_47_268 ();
 FILLCELL_X2 FILLER_47_273 ();
 FILLCELL_X8 FILLER_47_278 ();
 FILLCELL_X2 FILLER_47_286 ();
 FILLCELL_X1 FILLER_47_295 ();
 FILLCELL_X8 FILLER_47_303 ();
 FILLCELL_X4 FILLER_47_311 ();
 FILLCELL_X2 FILLER_47_315 ();
 FILLCELL_X1 FILLER_47_317 ();
 FILLCELL_X16 FILLER_47_345 ();
 FILLCELL_X4 FILLER_47_361 ();
 FILLCELL_X2 FILLER_47_365 ();
 FILLCELL_X1 FILLER_47_371 ();
 FILLCELL_X1 FILLER_47_375 ();
 FILLCELL_X4 FILLER_47_408 ();
 FILLCELL_X8 FILLER_47_417 ();
 FILLCELL_X2 FILLER_47_425 ();
 FILLCELL_X1 FILLER_47_427 ();
 FILLCELL_X4 FILLER_47_433 ();
 FILLCELL_X2 FILLER_47_437 ();
 FILLCELL_X2 FILLER_47_446 ();
 FILLCELL_X1 FILLER_47_448 ();
 FILLCELL_X4 FILLER_47_453 ();
 FILLCELL_X4 FILLER_47_470 ();
 FILLCELL_X2 FILLER_47_496 ();
 FILLCELL_X4 FILLER_47_502 ();
 FILLCELL_X2 FILLER_47_506 ();
 FILLCELL_X1 FILLER_47_508 ();
 FILLCELL_X4 FILLER_47_532 ();
 FILLCELL_X8 FILLER_47_543 ();
 FILLCELL_X2 FILLER_47_551 ();
 FILLCELL_X4 FILLER_47_587 ();
 FILLCELL_X4 FILLER_47_611 ();
 FILLCELL_X1 FILLER_47_615 ();
 FILLCELL_X1 FILLER_47_623 ();
 FILLCELL_X4 FILLER_47_655 ();
 FILLCELL_X2 FILLER_47_659 ();
 FILLCELL_X1 FILLER_47_661 ();
 FILLCELL_X4 FILLER_47_685 ();
 FILLCELL_X4 FILLER_47_700 ();
 FILLCELL_X1 FILLER_47_704 ();
 FILLCELL_X2 FILLER_47_749 ();
 FILLCELL_X4 FILLER_47_772 ();
 FILLCELL_X1 FILLER_47_776 ();
 FILLCELL_X4 FILLER_47_784 ();
 FILLCELL_X16 FILLER_47_792 ();
 FILLCELL_X1 FILLER_47_808 ();
 FILLCELL_X8 FILLER_47_825 ();
 FILLCELL_X8 FILLER_47_842 ();
 FILLCELL_X4 FILLER_47_850 ();
 FILLCELL_X1 FILLER_47_879 ();
 FILLCELL_X1 FILLER_47_890 ();
 FILLCELL_X1 FILLER_47_916 ();
 FILLCELL_X2 FILLER_47_930 ();
 FILLCELL_X1 FILLER_47_932 ();
 FILLCELL_X1 FILLER_47_946 ();
 FILLCELL_X4 FILLER_47_1002 ();
 FILLCELL_X4 FILLER_47_1009 ();
 FILLCELL_X1 FILLER_47_1013 ();
 FILLCELL_X1 FILLER_47_1023 ();
 FILLCELL_X1 FILLER_47_1045 ();
 FILLCELL_X1 FILLER_47_1058 ();
 FILLCELL_X1 FILLER_47_1069 ();
 FILLCELL_X16 FILLER_47_1103 ();
 FILLCELL_X2 FILLER_47_1119 ();
 FILLCELL_X1 FILLER_47_1121 ();
 FILLCELL_X1 FILLER_47_1128 ();
 FILLCELL_X4 FILLER_47_1132 ();
 FILLCELL_X1 FILLER_47_1136 ();
 FILLCELL_X1 FILLER_47_1147 ();
 FILLCELL_X1 FILLER_47_1154 ();
 FILLCELL_X8 FILLER_47_1161 ();
 FILLCELL_X1 FILLER_47_1169 ();
 FILLCELL_X2 FILLER_47_1194 ();
 FILLCELL_X1 FILLER_47_1202 ();
 FILLCELL_X2 FILLER_47_1209 ();
 FILLCELL_X1 FILLER_47_1211 ();
 FILLCELL_X4 FILLER_47_1246 ();
 FILLCELL_X2 FILLER_47_1250 ();
 FILLCELL_X1 FILLER_47_1252 ();
 FILLCELL_X2 FILLER_47_1260 ();
 FILLCELL_X1 FILLER_47_1262 ();
 FILLCELL_X2 FILLER_47_1311 ();
 FILLCELL_X1 FILLER_47_1313 ();
 FILLCELL_X8 FILLER_47_1334 ();
 FILLCELL_X4 FILLER_47_1342 ();
 FILLCELL_X2 FILLER_47_1346 ();
 FILLCELL_X1 FILLER_47_1348 ();
 FILLCELL_X1 FILLER_47_1354 ();
 FILLCELL_X8 FILLER_47_1362 ();
 FILLCELL_X2 FILLER_47_1370 ();
 FILLCELL_X1 FILLER_47_1372 ();
 FILLCELL_X1 FILLER_47_1378 ();
 FILLCELL_X2 FILLER_47_1386 ();
 FILLCELL_X2 FILLER_47_1397 ();
 FILLCELL_X1 FILLER_47_1399 ();
 FILLCELL_X4 FILLER_47_1411 ();
 FILLCELL_X2 FILLER_47_1415 ();
 FILLCELL_X1 FILLER_47_1417 ();
 FILLCELL_X8 FILLER_47_1434 ();
 FILLCELL_X2 FILLER_47_1442 ();
 FILLCELL_X1 FILLER_47_1444 ();
 FILLCELL_X8 FILLER_47_1482 ();
 FILLCELL_X1 FILLER_47_1490 ();
 FILLCELL_X4 FILLER_47_1495 ();
 FILLCELL_X2 FILLER_47_1499 ();
 FILLCELL_X8 FILLER_47_1510 ();
 FILLCELL_X2 FILLER_47_1518 ();
 FILLCELL_X1 FILLER_47_1520 ();
 FILLCELL_X2 FILLER_47_1525 ();
 FILLCELL_X1 FILLER_47_1527 ();
 FILLCELL_X1 FILLER_47_1533 ();
 FILLCELL_X4 FILLER_47_1541 ();
 FILLCELL_X2 FILLER_47_1545 ();
 FILLCELL_X1 FILLER_47_1547 ();
 FILLCELL_X2 FILLER_47_1559 ();
 FILLCELL_X4 FILLER_47_1565 ();
 FILLCELL_X2 FILLER_47_1569 ();
 FILLCELL_X1 FILLER_47_1571 ();
 FILLCELL_X4 FILLER_47_1583 ();
 FILLCELL_X8 FILLER_47_1598 ();
 FILLCELL_X2 FILLER_47_1610 ();
 FILLCELL_X2 FILLER_47_1620 ();
 FILLCELL_X16 FILLER_47_1629 ();
 FILLCELL_X4 FILLER_47_1645 ();
 FILLCELL_X2 FILLER_47_1649 ();
 FILLCELL_X4 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_8 ();
 FILLCELL_X32 FILLER_48_40 ();
 FILLCELL_X32 FILLER_48_72 ();
 FILLCELL_X32 FILLER_48_104 ();
 FILLCELL_X32 FILLER_48_136 ();
 FILLCELL_X16 FILLER_48_168 ();
 FILLCELL_X8 FILLER_48_184 ();
 FILLCELL_X4 FILLER_48_192 ();
 FILLCELL_X1 FILLER_48_204 ();
 FILLCELL_X8 FILLER_48_215 ();
 FILLCELL_X4 FILLER_48_223 ();
 FILLCELL_X1 FILLER_48_227 ();
 FILLCELL_X1 FILLER_48_260 ();
 FILLCELL_X1 FILLER_48_265 ();
 FILLCELL_X1 FILLER_48_273 ();
 FILLCELL_X4 FILLER_48_285 ();
 FILLCELL_X2 FILLER_48_314 ();
 FILLCELL_X2 FILLER_48_322 ();
 FILLCELL_X4 FILLER_48_331 ();
 FILLCELL_X1 FILLER_48_335 ();
 FILLCELL_X4 FILLER_48_340 ();
 FILLCELL_X2 FILLER_48_348 ();
 FILLCELL_X1 FILLER_48_350 ();
 FILLCELL_X8 FILLER_48_373 ();
 FILLCELL_X2 FILLER_48_381 ();
 FILLCELL_X4 FILLER_48_403 ();
 FILLCELL_X2 FILLER_48_407 ();
 FILLCELL_X1 FILLER_48_409 ();
 FILLCELL_X4 FILLER_48_417 ();
 FILLCELL_X1 FILLER_48_421 ();
 FILLCELL_X2 FILLER_48_426 ();
 FILLCELL_X1 FILLER_48_428 ();
 FILLCELL_X4 FILLER_48_451 ();
 FILLCELL_X2 FILLER_48_455 ();
 FILLCELL_X2 FILLER_48_501 ();
 FILLCELL_X8 FILLER_48_545 ();
 FILLCELL_X4 FILLER_48_553 ();
 FILLCELL_X2 FILLER_48_557 ();
 FILLCELL_X2 FILLER_48_563 ();
 FILLCELL_X8 FILLER_48_575 ();
 FILLCELL_X4 FILLER_48_583 ();
 FILLCELL_X1 FILLER_48_587 ();
 FILLCELL_X1 FILLER_48_598 ();
 FILLCELL_X4 FILLER_48_610 ();
 FILLCELL_X1 FILLER_48_614 ();
 FILLCELL_X4 FILLER_48_619 ();
 FILLCELL_X1 FILLER_48_623 ();
 FILLCELL_X1 FILLER_48_632 ();
 FILLCELL_X8 FILLER_48_640 ();
 FILLCELL_X4 FILLER_48_662 ();
 FILLCELL_X2 FILLER_48_666 ();
 FILLCELL_X16 FILLER_48_687 ();
 FILLCELL_X4 FILLER_48_703 ();
 FILLCELL_X1 FILLER_48_707 ();
 FILLCELL_X4 FILLER_48_729 ();
 FILLCELL_X2 FILLER_48_733 ();
 FILLCELL_X4 FILLER_48_763 ();
 FILLCELL_X1 FILLER_48_767 ();
 FILLCELL_X8 FILLER_48_777 ();
 FILLCELL_X1 FILLER_48_785 ();
 FILLCELL_X8 FILLER_48_799 ();
 FILLCELL_X8 FILLER_48_848 ();
 FILLCELL_X2 FILLER_48_856 ();
 FILLCELL_X1 FILLER_48_858 ();
 FILLCELL_X4 FILLER_48_891 ();
 FILLCELL_X1 FILLER_48_895 ();
 FILLCELL_X4 FILLER_48_901 ();
 FILLCELL_X4 FILLER_48_922 ();
 FILLCELL_X2 FILLER_48_926 ();
 FILLCELL_X1 FILLER_48_928 ();
 FILLCELL_X4 FILLER_48_941 ();
 FILLCELL_X2 FILLER_48_945 ();
 FILLCELL_X4 FILLER_48_956 ();
 FILLCELL_X1 FILLER_48_960 ();
 FILLCELL_X4 FILLER_48_968 ();
 FILLCELL_X1 FILLER_48_972 ();
 FILLCELL_X1 FILLER_48_979 ();
 FILLCELL_X4 FILLER_48_991 ();
 FILLCELL_X1 FILLER_48_995 ();
 FILLCELL_X2 FILLER_48_1003 ();
 FILLCELL_X8 FILLER_48_1018 ();
 FILLCELL_X2 FILLER_48_1026 ();
 FILLCELL_X4 FILLER_48_1040 ();
 FILLCELL_X2 FILLER_48_1044 ();
 FILLCELL_X8 FILLER_48_1055 ();
 FILLCELL_X4 FILLER_48_1094 ();
 FILLCELL_X8 FILLER_48_1104 ();
 FILLCELL_X2 FILLER_48_1112 ();
 FILLCELL_X1 FILLER_48_1114 ();
 FILLCELL_X1 FILLER_48_1120 ();
 FILLCELL_X2 FILLER_48_1123 ();
 FILLCELL_X1 FILLER_48_1139 ();
 FILLCELL_X1 FILLER_48_1152 ();
 FILLCELL_X4 FILLER_48_1190 ();
 FILLCELL_X1 FILLER_48_1194 ();
 FILLCELL_X8 FILLER_48_1207 ();
 FILLCELL_X2 FILLER_48_1215 ();
 FILLCELL_X1 FILLER_48_1277 ();
 FILLCELL_X1 FILLER_48_1328 ();
 FILLCELL_X4 FILLER_48_1349 ();
 FILLCELL_X8 FILLER_48_1366 ();
 FILLCELL_X1 FILLER_48_1387 ();
 FILLCELL_X4 FILLER_48_1404 ();
 FILLCELL_X2 FILLER_48_1408 ();
 FILLCELL_X2 FILLER_48_1423 ();
 FILLCELL_X1 FILLER_48_1432 ();
 FILLCELL_X16 FILLER_48_1440 ();
 FILLCELL_X2 FILLER_48_1456 ();
 FILLCELL_X2 FILLER_48_1467 ();
 FILLCELL_X4 FILLER_48_1484 ();
 FILLCELL_X1 FILLER_48_1488 ();
 FILLCELL_X1 FILLER_48_1492 ();
 FILLCELL_X4 FILLER_48_1500 ();
 FILLCELL_X2 FILLER_48_1508 ();
 FILLCELL_X1 FILLER_48_1510 ();
 FILLCELL_X32 FILLER_48_1525 ();
 FILLCELL_X2 FILLER_48_1557 ();
 FILLCELL_X1 FILLER_48_1579 ();
 FILLCELL_X16 FILLER_48_1589 ();
 FILLCELL_X2 FILLER_48_1605 ();
 FILLCELL_X1 FILLER_48_1620 ();
 FILLCELL_X2 FILLER_48_1624 ();
 FILLCELL_X1 FILLER_48_1626 ();
 FILLCELL_X16 FILLER_48_1631 ();
 FILLCELL_X4 FILLER_48_1647 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X16 FILLER_49_161 ();
 FILLCELL_X2 FILLER_49_177 ();
 FILLCELL_X2 FILLER_49_207 ();
 FILLCELL_X8 FILLER_49_215 ();
 FILLCELL_X2 FILLER_49_223 ();
 FILLCELL_X1 FILLER_49_225 ();
 FILLCELL_X4 FILLER_49_239 ();
 FILLCELL_X1 FILLER_49_272 ();
 FILLCELL_X2 FILLER_49_281 ();
 FILLCELL_X8 FILLER_49_307 ();
 FILLCELL_X4 FILLER_49_315 ();
 FILLCELL_X1 FILLER_49_319 ();
 FILLCELL_X16 FILLER_49_353 ();
 FILLCELL_X4 FILLER_49_369 ();
 FILLCELL_X2 FILLER_49_393 ();
 FILLCELL_X1 FILLER_49_395 ();
 FILLCELL_X4 FILLER_49_438 ();
 FILLCELL_X4 FILLER_49_448 ();
 FILLCELL_X2 FILLER_49_452 ();
 FILLCELL_X1 FILLER_49_454 ();
 FILLCELL_X8 FILLER_49_466 ();
 FILLCELL_X8 FILLER_49_481 ();
 FILLCELL_X4 FILLER_49_489 ();
 FILLCELL_X2 FILLER_49_493 ();
 FILLCELL_X1 FILLER_49_495 ();
 FILLCELL_X8 FILLER_49_503 ();
 FILLCELL_X4 FILLER_49_518 ();
 FILLCELL_X1 FILLER_49_522 ();
 FILLCELL_X1 FILLER_49_530 ();
 FILLCELL_X16 FILLER_49_566 ();
 FILLCELL_X1 FILLER_49_582 ();
 FILLCELL_X1 FILLER_49_595 ();
 FILLCELL_X1 FILLER_49_604 ();
 FILLCELL_X1 FILLER_49_609 ();
 FILLCELL_X1 FILLER_49_630 ();
 FILLCELL_X1 FILLER_49_651 ();
 FILLCELL_X2 FILLER_49_672 ();
 FILLCELL_X2 FILLER_49_694 ();
 FILLCELL_X2 FILLER_49_702 ();
 FILLCELL_X1 FILLER_49_704 ();
 FILLCELL_X1 FILLER_49_711 ();
 FILLCELL_X2 FILLER_49_716 ();
 FILLCELL_X1 FILLER_49_718 ();
 FILLCELL_X8 FILLER_49_735 ();
 FILLCELL_X2 FILLER_49_743 ();
 FILLCELL_X1 FILLER_49_745 ();
 FILLCELL_X4 FILLER_49_769 ();
 FILLCELL_X4 FILLER_49_833 ();
 FILLCELL_X1 FILLER_49_837 ();
 FILLCELL_X2 FILLER_49_856 ();
 FILLCELL_X1 FILLER_49_858 ();
 FILLCELL_X2 FILLER_49_864 ();
 FILLCELL_X1 FILLER_49_866 ();
 FILLCELL_X2 FILLER_49_871 ();
 FILLCELL_X2 FILLER_49_880 ();
 FILLCELL_X2 FILLER_49_892 ();
 FILLCELL_X4 FILLER_49_936 ();
 FILLCELL_X2 FILLER_49_967 ();
 FILLCELL_X1 FILLER_49_969 ();
 FILLCELL_X2 FILLER_49_975 ();
 FILLCELL_X4 FILLER_49_982 ();
 FILLCELL_X8 FILLER_49_1003 ();
 FILLCELL_X2 FILLER_49_1011 ();
 FILLCELL_X8 FILLER_49_1035 ();
 FILLCELL_X1 FILLER_49_1043 ();
 FILLCELL_X1 FILLER_49_1072 ();
 FILLCELL_X4 FILLER_49_1085 ();
 FILLCELL_X1 FILLER_49_1111 ();
 FILLCELL_X8 FILLER_49_1137 ();
 FILLCELL_X1 FILLER_49_1145 ();
 FILLCELL_X2 FILLER_49_1148 ();
 FILLCELL_X1 FILLER_49_1150 ();
 FILLCELL_X4 FILLER_49_1158 ();
 FILLCELL_X2 FILLER_49_1162 ();
 FILLCELL_X1 FILLER_49_1170 ();
 FILLCELL_X1 FILLER_49_1187 ();
 FILLCELL_X8 FILLER_49_1206 ();
 FILLCELL_X1 FILLER_49_1214 ();
 FILLCELL_X2 FILLER_49_1222 ();
 FILLCELL_X4 FILLER_49_1237 ();
 FILLCELL_X4 FILLER_49_1248 ();
 FILLCELL_X1 FILLER_49_1252 ();
 FILLCELL_X2 FILLER_49_1278 ();
 FILLCELL_X4 FILLER_49_1293 ();
 FILLCELL_X4 FILLER_49_1300 ();
 FILLCELL_X1 FILLER_49_1304 ();
 FILLCELL_X16 FILLER_49_1332 ();
 FILLCELL_X4 FILLER_49_1348 ();
 FILLCELL_X1 FILLER_49_1352 ();
 FILLCELL_X32 FILLER_49_1373 ();
 FILLCELL_X8 FILLER_49_1405 ();
 FILLCELL_X4 FILLER_49_1413 ();
 FILLCELL_X1 FILLER_49_1417 ();
 FILLCELL_X16 FILLER_49_1422 ();
 FILLCELL_X8 FILLER_49_1438 ();
 FILLCELL_X4 FILLER_49_1446 ();
 FILLCELL_X2 FILLER_49_1465 ();
 FILLCELL_X1 FILLER_49_1471 ();
 FILLCELL_X1 FILLER_49_1479 ();
 FILLCELL_X1 FILLER_49_1488 ();
 FILLCELL_X2 FILLER_49_1496 ();
 FILLCELL_X1 FILLER_49_1498 ();
 FILLCELL_X4 FILLER_49_1510 ();
 FILLCELL_X2 FILLER_49_1514 ();
 FILLCELL_X2 FILLER_49_1533 ();
 FILLCELL_X2 FILLER_49_1557 ();
 FILLCELL_X1 FILLER_49_1563 ();
 FILLCELL_X2 FILLER_49_1568 ();
 FILLCELL_X2 FILLER_49_1575 ();
 FILLCELL_X2 FILLER_49_1581 ();
 FILLCELL_X2 FILLER_49_1587 ();
 FILLCELL_X4 FILLER_49_1593 ();
 FILLCELL_X2 FILLER_49_1622 ();
 FILLCELL_X16 FILLER_49_1628 ();
 FILLCELL_X4 FILLER_49_1644 ();
 FILLCELL_X2 FILLER_49_1648 ();
 FILLCELL_X1 FILLER_49_1650 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X16 FILLER_50_161 ();
 FILLCELL_X1 FILLER_50_177 ();
 FILLCELL_X8 FILLER_50_221 ();
 FILLCELL_X4 FILLER_50_242 ();
 FILLCELL_X2 FILLER_50_246 ();
 FILLCELL_X1 FILLER_50_248 ();
 FILLCELL_X2 FILLER_50_252 ();
 FILLCELL_X1 FILLER_50_254 ();
 FILLCELL_X1 FILLER_50_267 ();
 FILLCELL_X1 FILLER_50_270 ();
 FILLCELL_X16 FILLER_50_282 ();
 FILLCELL_X1 FILLER_50_298 ();
 FILLCELL_X2 FILLER_50_306 ();
 FILLCELL_X4 FILLER_50_317 ();
 FILLCELL_X4 FILLER_50_328 ();
 FILLCELL_X1 FILLER_50_332 ();
 FILLCELL_X4 FILLER_50_360 ();
 FILLCELL_X2 FILLER_50_364 ();
 FILLCELL_X1 FILLER_50_387 ();
 FILLCELL_X8 FILLER_50_415 ();
 FILLCELL_X2 FILLER_50_423 ();
 FILLCELL_X4 FILLER_50_428 ();
 FILLCELL_X8 FILLER_50_442 ();
 FILLCELL_X2 FILLER_50_450 ();
 FILLCELL_X2 FILLER_50_459 ();
 FILLCELL_X2 FILLER_50_468 ();
 FILLCELL_X1 FILLER_50_470 ();
 FILLCELL_X1 FILLER_50_478 ();
 FILLCELL_X2 FILLER_50_492 ();
 FILLCELL_X1 FILLER_50_494 ();
 FILLCELL_X2 FILLER_50_522 ();
 FILLCELL_X4 FILLER_50_583 ();
 FILLCELL_X2 FILLER_50_613 ();
 FILLCELL_X8 FILLER_50_622 ();
 FILLCELL_X1 FILLER_50_630 ();
 FILLCELL_X4 FILLER_50_632 ();
 FILLCELL_X1 FILLER_50_636 ();
 FILLCELL_X4 FILLER_50_644 ();
 FILLCELL_X1 FILLER_50_648 ();
 FILLCELL_X1 FILLER_50_701 ();
 FILLCELL_X4 FILLER_50_714 ();
 FILLCELL_X2 FILLER_50_718 ();
 FILLCELL_X4 FILLER_50_741 ();
 FILLCELL_X1 FILLER_50_752 ();
 FILLCELL_X2 FILLER_50_760 ();
 FILLCELL_X1 FILLER_50_762 ();
 FILLCELL_X1 FILLER_50_770 ();
 FILLCELL_X4 FILLER_50_784 ();
 FILLCELL_X8 FILLER_50_795 ();
 FILLCELL_X32 FILLER_50_823 ();
 FILLCELL_X8 FILLER_50_855 ();
 FILLCELL_X4 FILLER_50_863 ();
 FILLCELL_X2 FILLER_50_867 ();
 FILLCELL_X1 FILLER_50_869 ();
 FILLCELL_X1 FILLER_50_874 ();
 FILLCELL_X1 FILLER_50_879 ();
 FILLCELL_X1 FILLER_50_890 ();
 FILLCELL_X2 FILLER_50_922 ();
 FILLCELL_X1 FILLER_50_924 ();
 FILLCELL_X8 FILLER_50_930 ();
 FILLCELL_X4 FILLER_50_938 ();
 FILLCELL_X2 FILLER_50_942 ();
 FILLCELL_X1 FILLER_50_944 ();
 FILLCELL_X1 FILLER_50_979 ();
 FILLCELL_X1 FILLER_50_1000 ();
 FILLCELL_X1 FILLER_50_1023 ();
 FILLCELL_X4 FILLER_50_1031 ();
 FILLCELL_X2 FILLER_50_1035 ();
 FILLCELL_X1 FILLER_50_1037 ();
 FILLCELL_X1 FILLER_50_1050 ();
 FILLCELL_X1 FILLER_50_1070 ();
 FILLCELL_X8 FILLER_50_1074 ();
 FILLCELL_X4 FILLER_50_1094 ();
 FILLCELL_X2 FILLER_50_1098 ();
 FILLCELL_X2 FILLER_50_1106 ();
 FILLCELL_X1 FILLER_50_1108 ();
 FILLCELL_X2 FILLER_50_1111 ();
 FILLCELL_X1 FILLER_50_1113 ();
 FILLCELL_X2 FILLER_50_1123 ();
 FILLCELL_X8 FILLER_50_1141 ();
 FILLCELL_X2 FILLER_50_1149 ();
 FILLCELL_X1 FILLER_50_1151 ();
 FILLCELL_X1 FILLER_50_1158 ();
 FILLCELL_X8 FILLER_50_1168 ();
 FILLCELL_X2 FILLER_50_1176 ();
 FILLCELL_X1 FILLER_50_1178 ();
 FILLCELL_X4 FILLER_50_1185 ();
 FILLCELL_X2 FILLER_50_1189 ();
 FILLCELL_X8 FILLER_50_1197 ();
 FILLCELL_X4 FILLER_50_1205 ();
 FILLCELL_X1 FILLER_50_1209 ();
 FILLCELL_X2 FILLER_50_1224 ();
 FILLCELL_X1 FILLER_50_1226 ();
 FILLCELL_X8 FILLER_50_1230 ();
 FILLCELL_X1 FILLER_50_1238 ();
 FILLCELL_X4 FILLER_50_1259 ();
 FILLCELL_X1 FILLER_50_1263 ();
 FILLCELL_X2 FILLER_50_1271 ();
 FILLCELL_X4 FILLER_50_1280 ();
 FILLCELL_X1 FILLER_50_1284 ();
 FILLCELL_X8 FILLER_50_1288 ();
 FILLCELL_X2 FILLER_50_1303 ();
 FILLCELL_X8 FILLER_50_1340 ();
 FILLCELL_X4 FILLER_50_1348 ();
 FILLCELL_X2 FILLER_50_1352 ();
 FILLCELL_X32 FILLER_50_1374 ();
 FILLCELL_X4 FILLER_50_1406 ();
 FILLCELL_X8 FILLER_50_1428 ();
 FILLCELL_X1 FILLER_50_1436 ();
 FILLCELL_X8 FILLER_50_1464 ();
 FILLCELL_X4 FILLER_50_1472 ();
 FILLCELL_X8 FILLER_50_1507 ();
 FILLCELL_X2 FILLER_50_1515 ();
 FILLCELL_X1 FILLER_50_1517 ();
 FILLCELL_X4 FILLER_50_1528 ();
 FILLCELL_X1 FILLER_50_1541 ();
 FILLCELL_X8 FILLER_50_1573 ();
 FILLCELL_X2 FILLER_50_1581 ();
 FILLCELL_X1 FILLER_50_1592 ();
 FILLCELL_X16 FILLER_50_1632 ();
 FILLCELL_X2 FILLER_50_1648 ();
 FILLCELL_X1 FILLER_50_1650 ();
 FILLCELL_X8 FILLER_51_1 ();
 FILLCELL_X2 FILLER_51_9 ();
 FILLCELL_X1 FILLER_51_11 ();
 FILLCELL_X32 FILLER_51_15 ();
 FILLCELL_X32 FILLER_51_47 ();
 FILLCELL_X32 FILLER_51_79 ();
 FILLCELL_X32 FILLER_51_111 ();
 FILLCELL_X32 FILLER_51_143 ();
 FILLCELL_X16 FILLER_51_175 ();
 FILLCELL_X1 FILLER_51_252 ();
 FILLCELL_X1 FILLER_51_257 ();
 FILLCELL_X2 FILLER_51_262 ();
 FILLCELL_X2 FILLER_51_268 ();
 FILLCELL_X4 FILLER_51_279 ();
 FILLCELL_X2 FILLER_51_285 ();
 FILLCELL_X2 FILLER_51_297 ();
 FILLCELL_X1 FILLER_51_299 ();
 FILLCELL_X4 FILLER_51_305 ();
 FILLCELL_X1 FILLER_51_309 ();
 FILLCELL_X2 FILLER_51_317 ();
 FILLCELL_X4 FILLER_51_329 ();
 FILLCELL_X2 FILLER_51_333 ();
 FILLCELL_X1 FILLER_51_344 ();
 FILLCELL_X2 FILLER_51_357 ();
 FILLCELL_X1 FILLER_51_359 ();
 FILLCELL_X2 FILLER_51_380 ();
 FILLCELL_X2 FILLER_51_395 ();
 FILLCELL_X2 FILLER_51_403 ();
 FILLCELL_X1 FILLER_51_405 ();
 FILLCELL_X4 FILLER_51_433 ();
 FILLCELL_X1 FILLER_51_437 ();
 FILLCELL_X1 FILLER_51_488 ();
 FILLCELL_X8 FILLER_51_509 ();
 FILLCELL_X8 FILLER_51_542 ();
 FILLCELL_X2 FILLER_51_550 ();
 FILLCELL_X1 FILLER_51_552 ();
 FILLCELL_X16 FILLER_51_556 ();
 FILLCELL_X8 FILLER_51_572 ();
 FILLCELL_X4 FILLER_51_580 ();
 FILLCELL_X8 FILLER_51_616 ();
 FILLCELL_X1 FILLER_51_624 ();
 FILLCELL_X4 FILLER_51_645 ();
 FILLCELL_X2 FILLER_51_656 ();
 FILLCELL_X2 FILLER_51_665 ();
 FILLCELL_X1 FILLER_51_667 ();
 FILLCELL_X2 FILLER_51_672 ();
 FILLCELL_X4 FILLER_51_685 ();
 FILLCELL_X2 FILLER_51_701 ();
 FILLCELL_X2 FILLER_51_709 ();
 FILLCELL_X1 FILLER_51_711 ();
 FILLCELL_X1 FILLER_51_715 ();
 FILLCELL_X4 FILLER_51_725 ();
 FILLCELL_X4 FILLER_51_732 ();
 FILLCELL_X1 FILLER_51_736 ();
 FILLCELL_X2 FILLER_51_757 ();
 FILLCELL_X1 FILLER_51_770 ();
 FILLCELL_X2 FILLER_51_809 ();
 FILLCELL_X8 FILLER_51_831 ();
 FILLCELL_X1 FILLER_51_839 ();
 FILLCELL_X4 FILLER_51_869 ();
 FILLCELL_X8 FILLER_51_879 ();
 FILLCELL_X1 FILLER_51_887 ();
 FILLCELL_X8 FILLER_51_892 ();
 FILLCELL_X4 FILLER_51_900 ();
 FILLCELL_X2 FILLER_51_904 ();
 FILLCELL_X2 FILLER_51_926 ();
 FILLCELL_X2 FILLER_51_930 ();
 FILLCELL_X4 FILLER_51_937 ();
 FILLCELL_X2 FILLER_51_952 ();
 FILLCELL_X2 FILLER_51_959 ();
 FILLCELL_X1 FILLER_51_961 ();
 FILLCELL_X2 FILLER_51_967 ();
 FILLCELL_X1 FILLER_51_969 ();
 FILLCELL_X16 FILLER_51_978 ();
 FILLCELL_X2 FILLER_51_994 ();
 FILLCELL_X1 FILLER_51_996 ();
 FILLCELL_X1 FILLER_51_999 ();
 FILLCELL_X8 FILLER_51_1007 ();
 FILLCELL_X1 FILLER_51_1015 ();
 FILLCELL_X2 FILLER_51_1023 ();
 FILLCELL_X1 FILLER_51_1025 ();
 FILLCELL_X4 FILLER_51_1039 ();
 FILLCELL_X2 FILLER_51_1043 ();
 FILLCELL_X4 FILLER_51_1067 ();
 FILLCELL_X2 FILLER_51_1071 ();
 FILLCELL_X1 FILLER_51_1089 ();
 FILLCELL_X2 FILLER_51_1101 ();
 FILLCELL_X2 FILLER_51_1120 ();
 FILLCELL_X2 FILLER_51_1150 ();
 FILLCELL_X1 FILLER_51_1152 ();
 FILLCELL_X4 FILLER_51_1165 ();
 FILLCELL_X2 FILLER_51_1169 ();
 FILLCELL_X2 FILLER_51_1187 ();
 FILLCELL_X1 FILLER_51_1189 ();
 FILLCELL_X8 FILLER_51_1200 ();
 FILLCELL_X1 FILLER_51_1208 ();
 FILLCELL_X4 FILLER_51_1216 ();
 FILLCELL_X4 FILLER_51_1236 ();
 FILLCELL_X2 FILLER_51_1260 ();
 FILLCELL_X1 FILLER_51_1262 ();
 FILLCELL_X4 FILLER_51_1264 ();
 FILLCELL_X8 FILLER_51_1295 ();
 FILLCELL_X2 FILLER_51_1303 ();
 FILLCELL_X1 FILLER_51_1305 ();
 FILLCELL_X2 FILLER_51_1333 ();
 FILLCELL_X1 FILLER_51_1335 ();
 FILLCELL_X4 FILLER_51_1350 ();
 FILLCELL_X8 FILLER_51_1376 ();
 FILLCELL_X4 FILLER_51_1384 ();
 FILLCELL_X2 FILLER_51_1388 ();
 FILLCELL_X1 FILLER_51_1390 ();
 FILLCELL_X2 FILLER_51_1418 ();
 FILLCELL_X2 FILLER_51_1434 ();
 FILLCELL_X4 FILLER_51_1443 ();
 FILLCELL_X4 FILLER_51_1450 ();
 FILLCELL_X8 FILLER_51_1477 ();
 FILLCELL_X1 FILLER_51_1485 ();
 FILLCELL_X4 FILLER_51_1493 ();
 FILLCELL_X2 FILLER_51_1497 ();
 FILLCELL_X8 FILLER_51_1505 ();
 FILLCELL_X1 FILLER_51_1513 ();
 FILLCELL_X2 FILLER_51_1520 ();
 FILLCELL_X1 FILLER_51_1531 ();
 FILLCELL_X2 FILLER_51_1544 ();
 FILLCELL_X1 FILLER_51_1546 ();
 FILLCELL_X8 FILLER_51_1550 ();
 FILLCELL_X2 FILLER_51_1558 ();
 FILLCELL_X1 FILLER_51_1560 ();
 FILLCELL_X8 FILLER_51_1564 ();
 FILLCELL_X4 FILLER_51_1572 ();
 FILLCELL_X1 FILLER_51_1593 ();
 FILLCELL_X1 FILLER_51_1598 ();
 FILLCELL_X1 FILLER_51_1620 ();
 FILLCELL_X8 FILLER_51_1636 ();
 FILLCELL_X4 FILLER_51_1644 ();
 FILLCELL_X2 FILLER_51_1648 ();
 FILLCELL_X1 FILLER_51_1650 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X8 FILLER_52_161 ();
 FILLCELL_X2 FILLER_52_169 ();
 FILLCELL_X1 FILLER_52_171 ();
 FILLCELL_X16 FILLER_52_192 ();
 FILLCELL_X4 FILLER_52_208 ();
 FILLCELL_X2 FILLER_52_212 ();
 FILLCELL_X1 FILLER_52_214 ();
 FILLCELL_X2 FILLER_52_226 ();
 FILLCELL_X1 FILLER_52_228 ();
 FILLCELL_X2 FILLER_52_240 ();
 FILLCELL_X1 FILLER_52_242 ();
 FILLCELL_X16 FILLER_52_247 ();
 FILLCELL_X2 FILLER_52_263 ();
 FILLCELL_X2 FILLER_52_272 ();
 FILLCELL_X4 FILLER_52_306 ();
 FILLCELL_X2 FILLER_52_310 ();
 FILLCELL_X1 FILLER_52_312 ();
 FILLCELL_X2 FILLER_52_318 ();
 FILLCELL_X1 FILLER_52_320 ();
 FILLCELL_X1 FILLER_52_326 ();
 FILLCELL_X1 FILLER_52_354 ();
 FILLCELL_X2 FILLER_52_375 ();
 FILLCELL_X2 FILLER_52_384 ();
 FILLCELL_X4 FILLER_52_406 ();
 FILLCELL_X2 FILLER_52_419 ();
 FILLCELL_X8 FILLER_52_448 ();
 FILLCELL_X2 FILLER_52_456 ();
 FILLCELL_X1 FILLER_52_458 ();
 FILLCELL_X1 FILLER_52_471 ();
 FILLCELL_X2 FILLER_52_479 ();
 FILLCELL_X8 FILLER_52_487 ();
 FILLCELL_X1 FILLER_52_495 ();
 FILLCELL_X1 FILLER_52_510 ();
 FILLCELL_X8 FILLER_52_515 ();
 FILLCELL_X4 FILLER_52_523 ();
 FILLCELL_X1 FILLER_52_527 ();
 FILLCELL_X16 FILLER_52_535 ();
 FILLCELL_X4 FILLER_52_551 ();
 FILLCELL_X1 FILLER_52_555 ();
 FILLCELL_X4 FILLER_52_560 ();
 FILLCELL_X2 FILLER_52_564 ();
 FILLCELL_X1 FILLER_52_566 ();
 FILLCELL_X1 FILLER_52_617 ();
 FILLCELL_X8 FILLER_52_622 ();
 FILLCELL_X1 FILLER_52_630 ();
 FILLCELL_X1 FILLER_52_632 ();
 FILLCELL_X1 FILLER_52_647 ();
 FILLCELL_X4 FILLER_52_690 ();
 FILLCELL_X1 FILLER_52_714 ();
 FILLCELL_X2 FILLER_52_723 ();
 FILLCELL_X2 FILLER_52_733 ();
 FILLCELL_X8 FILLER_52_742 ();
 FILLCELL_X1 FILLER_52_750 ();
 FILLCELL_X4 FILLER_52_754 ();
 FILLCELL_X2 FILLER_52_758 ();
 FILLCELL_X8 FILLER_52_793 ();
 FILLCELL_X32 FILLER_52_820 ();
 FILLCELL_X4 FILLER_52_852 ();
 FILLCELL_X2 FILLER_52_856 ();
 FILLCELL_X8 FILLER_52_897 ();
 FILLCELL_X2 FILLER_52_908 ();
 FILLCELL_X2 FILLER_52_933 ();
 FILLCELL_X2 FILLER_52_946 ();
 FILLCELL_X1 FILLER_52_948 ();
 FILLCELL_X1 FILLER_52_995 ();
 FILLCELL_X1 FILLER_52_1001 ();
 FILLCELL_X4 FILLER_52_1007 ();
 FILLCELL_X4 FILLER_52_1014 ();
 FILLCELL_X2 FILLER_52_1029 ();
 FILLCELL_X1 FILLER_52_1031 ();
 FILLCELL_X4 FILLER_52_1038 ();
 FILLCELL_X2 FILLER_52_1042 ();
 FILLCELL_X1 FILLER_52_1056 ();
 FILLCELL_X4 FILLER_52_1064 ();
 FILLCELL_X2 FILLER_52_1075 ();
 FILLCELL_X8 FILLER_52_1080 ();
 FILLCELL_X4 FILLER_52_1088 ();
 FILLCELL_X1 FILLER_52_1110 ();
 FILLCELL_X1 FILLER_52_1134 ();
 FILLCELL_X4 FILLER_52_1142 ();
 FILLCELL_X4 FILLER_52_1151 ();
 FILLCELL_X8 FILLER_52_1173 ();
 FILLCELL_X1 FILLER_52_1181 ();
 FILLCELL_X2 FILLER_52_1207 ();
 FILLCELL_X1 FILLER_52_1209 ();
 FILLCELL_X8 FILLER_52_1216 ();
 FILLCELL_X4 FILLER_52_1224 ();
 FILLCELL_X2 FILLER_52_1228 ();
 FILLCELL_X1 FILLER_52_1230 ();
 FILLCELL_X2 FILLER_52_1245 ();
 FILLCELL_X4 FILLER_52_1252 ();
 FILLCELL_X1 FILLER_52_1256 ();
 FILLCELL_X1 FILLER_52_1264 ();
 FILLCELL_X1 FILLER_52_1272 ();
 FILLCELL_X4 FILLER_52_1305 ();
 FILLCELL_X8 FILLER_52_1323 ();
 FILLCELL_X1 FILLER_52_1331 ();
 FILLCELL_X1 FILLER_52_1346 ();
 FILLCELL_X2 FILLER_52_1372 ();
 FILLCELL_X1 FILLER_52_1374 ();
 FILLCELL_X8 FILLER_52_1382 ();
 FILLCELL_X4 FILLER_52_1390 ();
 FILLCELL_X1 FILLER_52_1394 ();
 FILLCELL_X4 FILLER_52_1409 ();
 FILLCELL_X2 FILLER_52_1413 ();
 FILLCELL_X2 FILLER_52_1427 ();
 FILLCELL_X1 FILLER_52_1434 ();
 FILLCELL_X2 FILLER_52_1463 ();
 FILLCELL_X4 FILLER_52_1470 ();
 FILLCELL_X4 FILLER_52_1483 ();
 FILLCELL_X1 FILLER_52_1516 ();
 FILLCELL_X8 FILLER_52_1525 ();
 FILLCELL_X1 FILLER_52_1533 ();
 FILLCELL_X4 FILLER_52_1539 ();
 FILLCELL_X1 FILLER_52_1543 ();
 FILLCELL_X4 FILLER_52_1548 ();
 FILLCELL_X1 FILLER_52_1552 ();
 FILLCELL_X4 FILLER_52_1566 ();
 FILLCELL_X2 FILLER_52_1570 ();
 FILLCELL_X1 FILLER_52_1591 ();
 FILLCELL_X1 FILLER_52_1601 ();
 FILLCELL_X2 FILLER_52_1607 ();
 FILLCELL_X2 FILLER_52_1613 ();
 FILLCELL_X1 FILLER_52_1619 ();
 FILLCELL_X16 FILLER_52_1629 ();
 FILLCELL_X4 FILLER_52_1645 ();
 FILLCELL_X2 FILLER_52_1649 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X16 FILLER_53_129 ();
 FILLCELL_X4 FILLER_53_145 ();
 FILLCELL_X2 FILLER_53_149 ();
 FILLCELL_X4 FILLER_53_205 ();
 FILLCELL_X2 FILLER_53_212 ();
 FILLCELL_X8 FILLER_53_245 ();
 FILLCELL_X4 FILLER_53_253 ();
 FILLCELL_X4 FILLER_53_271 ();
 FILLCELL_X4 FILLER_53_305 ();
 FILLCELL_X2 FILLER_53_309 ();
 FILLCELL_X1 FILLER_53_311 ();
 FILLCELL_X4 FILLER_53_332 ();
 FILLCELL_X2 FILLER_53_340 ();
 FILLCELL_X1 FILLER_53_342 ();
 FILLCELL_X2 FILLER_53_345 ();
 FILLCELL_X1 FILLER_53_347 ();
 FILLCELL_X16 FILLER_53_351 ();
 FILLCELL_X1 FILLER_53_367 ();
 FILLCELL_X8 FILLER_53_373 ();
 FILLCELL_X4 FILLER_53_381 ();
 FILLCELL_X2 FILLER_53_392 ();
 FILLCELL_X4 FILLER_53_405 ();
 FILLCELL_X2 FILLER_53_409 ();
 FILLCELL_X1 FILLER_53_411 ();
 FILLCELL_X4 FILLER_53_431 ();
 FILLCELL_X8 FILLER_53_445 ();
 FILLCELL_X2 FILLER_53_453 ();
 FILLCELL_X4 FILLER_53_482 ();
 FILLCELL_X2 FILLER_53_499 ();
 FILLCELL_X4 FILLER_53_511 ();
 FILLCELL_X1 FILLER_53_515 ();
 FILLCELL_X2 FILLER_53_538 ();
 FILLCELL_X1 FILLER_53_540 ();
 FILLCELL_X2 FILLER_53_561 ();
 FILLCELL_X2 FILLER_53_570 ();
 FILLCELL_X1 FILLER_53_572 ();
 FILLCELL_X4 FILLER_53_580 ();
 FILLCELL_X1 FILLER_53_584 ();
 FILLCELL_X4 FILLER_53_621 ();
 FILLCELL_X1 FILLER_53_625 ();
 FILLCELL_X1 FILLER_53_666 ();
 FILLCELL_X16 FILLER_53_674 ();
 FILLCELL_X1 FILLER_53_694 ();
 FILLCELL_X1 FILLER_53_722 ();
 FILLCELL_X8 FILLER_53_766 ();
 FILLCELL_X4 FILLER_53_774 ();
 FILLCELL_X1 FILLER_53_778 ();
 FILLCELL_X4 FILLER_53_803 ();
 FILLCELL_X2 FILLER_53_807 ();
 FILLCELL_X2 FILLER_53_816 ();
 FILLCELL_X1 FILLER_53_818 ();
 FILLCELL_X2 FILLER_53_851 ();
 FILLCELL_X1 FILLER_53_853 ();
 FILLCELL_X4 FILLER_53_859 ();
 FILLCELL_X1 FILLER_53_863 ();
 FILLCELL_X2 FILLER_53_896 ();
 FILLCELL_X1 FILLER_53_917 ();
 FILLCELL_X1 FILLER_53_922 ();
 FILLCELL_X2 FILLER_53_930 ();
 FILLCELL_X2 FILLER_53_936 ();
 FILLCELL_X16 FILLER_53_962 ();
 FILLCELL_X8 FILLER_53_978 ();
 FILLCELL_X4 FILLER_53_986 ();
 FILLCELL_X2 FILLER_53_990 ();
 FILLCELL_X1 FILLER_53_992 ();
 FILLCELL_X2 FILLER_53_1004 ();
 FILLCELL_X1 FILLER_53_1035 ();
 FILLCELL_X8 FILLER_53_1039 ();
 FILLCELL_X4 FILLER_53_1047 ();
 FILLCELL_X8 FILLER_53_1068 ();
 FILLCELL_X2 FILLER_53_1076 ();
 FILLCELL_X1 FILLER_53_1080 ();
 FILLCELL_X2 FILLER_53_1087 ();
 FILLCELL_X8 FILLER_53_1095 ();
 FILLCELL_X4 FILLER_53_1103 ();
 FILLCELL_X8 FILLER_53_1114 ();
 FILLCELL_X2 FILLER_53_1157 ();
 FILLCELL_X1 FILLER_53_1159 ();
 FILLCELL_X2 FILLER_53_1166 ();
 FILLCELL_X2 FILLER_53_1186 ();
 FILLCELL_X1 FILLER_53_1188 ();
 FILLCELL_X8 FILLER_53_1195 ();
 FILLCELL_X8 FILLER_53_1209 ();
 FILLCELL_X4 FILLER_53_1217 ();
 FILLCELL_X2 FILLER_53_1221 ();
 FILLCELL_X1 FILLER_53_1223 ();
 FILLCELL_X2 FILLER_53_1251 ();
 FILLCELL_X1 FILLER_53_1253 ();
 FILLCELL_X2 FILLER_53_1261 ();
 FILLCELL_X4 FILLER_53_1284 ();
 FILLCELL_X8 FILLER_53_1295 ();
 FILLCELL_X1 FILLER_53_1303 ();
 FILLCELL_X4 FILLER_53_1338 ();
 FILLCELL_X2 FILLER_53_1342 ();
 FILLCELL_X4 FILLER_53_1364 ();
 FILLCELL_X8 FILLER_53_1382 ();
 FILLCELL_X4 FILLER_53_1412 ();
 FILLCELL_X1 FILLER_53_1416 ();
 FILLCELL_X16 FILLER_53_1433 ();
 FILLCELL_X4 FILLER_53_1449 ();
 FILLCELL_X2 FILLER_53_1453 ();
 FILLCELL_X1 FILLER_53_1467 ();
 FILLCELL_X1 FILLER_53_1472 ();
 FILLCELL_X2 FILLER_53_1483 ();
 FILLCELL_X2 FILLER_53_1494 ();
 FILLCELL_X1 FILLER_53_1496 ();
 FILLCELL_X4 FILLER_53_1510 ();
 FILLCELL_X2 FILLER_53_1514 ();
 FILLCELL_X4 FILLER_53_1529 ();
 FILLCELL_X1 FILLER_53_1533 ();
 FILLCELL_X1 FILLER_53_1550 ();
 FILLCELL_X2 FILLER_53_1555 ();
 FILLCELL_X1 FILLER_53_1557 ();
 FILLCELL_X4 FILLER_53_1563 ();
 FILLCELL_X1 FILLER_53_1567 ();
 FILLCELL_X2 FILLER_53_1572 ();
 FILLCELL_X2 FILLER_53_1592 ();
 FILLCELL_X1 FILLER_53_1594 ();
 FILLCELL_X2 FILLER_53_1609 ();
 FILLCELL_X4 FILLER_53_1615 ();
 FILLCELL_X2 FILLER_53_1619 ();
 FILLCELL_X16 FILLER_53_1628 ();
 FILLCELL_X4 FILLER_53_1644 ();
 FILLCELL_X2 FILLER_53_1648 ();
 FILLCELL_X1 FILLER_53_1650 ();
 FILLCELL_X4 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_8 ();
 FILLCELL_X32 FILLER_54_40 ();
 FILLCELL_X32 FILLER_54_72 ();
 FILLCELL_X16 FILLER_54_104 ();
 FILLCELL_X8 FILLER_54_120 ();
 FILLCELL_X4 FILLER_54_128 ();
 FILLCELL_X1 FILLER_54_132 ();
 FILLCELL_X16 FILLER_54_189 ();
 FILLCELL_X8 FILLER_54_205 ();
 FILLCELL_X4 FILLER_54_213 ();
 FILLCELL_X8 FILLER_54_230 ();
 FILLCELL_X4 FILLER_54_238 ();
 FILLCELL_X1 FILLER_54_242 ();
 FILLCELL_X1 FILLER_54_257 ();
 FILLCELL_X1 FILLER_54_265 ();
 FILLCELL_X2 FILLER_54_273 ();
 FILLCELL_X4 FILLER_54_281 ();
 FILLCELL_X4 FILLER_54_289 ();
 FILLCELL_X2 FILLER_54_293 ();
 FILLCELL_X1 FILLER_54_295 ();
 FILLCELL_X1 FILLER_54_310 ();
 FILLCELL_X1 FILLER_54_335 ();
 FILLCELL_X8 FILLER_54_347 ();
 FILLCELL_X4 FILLER_54_355 ();
 FILLCELL_X8 FILLER_54_390 ();
 FILLCELL_X4 FILLER_54_398 ();
 FILLCELL_X2 FILLER_54_402 ();
 FILLCELL_X2 FILLER_54_408 ();
 FILLCELL_X1 FILLER_54_410 ();
 FILLCELL_X4 FILLER_54_438 ();
 FILLCELL_X8 FILLER_54_469 ();
 FILLCELL_X8 FILLER_54_480 ();
 FILLCELL_X4 FILLER_54_528 ();
 FILLCELL_X1 FILLER_54_532 ();
 FILLCELL_X4 FILLER_54_538 ();
 FILLCELL_X2 FILLER_54_569 ();
 FILLCELL_X2 FILLER_54_591 ();
 FILLCELL_X1 FILLER_54_593 ();
 FILLCELL_X2 FILLER_54_600 ();
 FILLCELL_X1 FILLER_54_602 ();
 FILLCELL_X2 FILLER_54_610 ();
 FILLCELL_X1 FILLER_54_612 ();
 FILLCELL_X8 FILLER_54_623 ();
 FILLCELL_X4 FILLER_54_659 ();
 FILLCELL_X1 FILLER_54_663 ();
 FILLCELL_X1 FILLER_54_696 ();
 FILLCELL_X4 FILLER_54_701 ();
 FILLCELL_X1 FILLER_54_705 ();
 FILLCELL_X1 FILLER_54_716 ();
 FILLCELL_X1 FILLER_54_721 ();
 FILLCELL_X1 FILLER_54_725 ();
 FILLCELL_X2 FILLER_54_736 ();
 FILLCELL_X4 FILLER_54_745 ();
 FILLCELL_X2 FILLER_54_749 ();
 FILLCELL_X2 FILLER_54_779 ();
 FILLCELL_X4 FILLER_54_788 ();
 FILLCELL_X2 FILLER_54_792 ();
 FILLCELL_X1 FILLER_54_807 ();
 FILLCELL_X16 FILLER_54_828 ();
 FILLCELL_X2 FILLER_54_844 ();
 FILLCELL_X1 FILLER_54_846 ();
 FILLCELL_X1 FILLER_54_871 ();
 FILLCELL_X2 FILLER_54_877 ();
 FILLCELL_X16 FILLER_54_886 ();
 FILLCELL_X4 FILLER_54_902 ();
 FILLCELL_X4 FILLER_54_928 ();
 FILLCELL_X1 FILLER_54_943 ();
 FILLCELL_X1 FILLER_54_959 ();
 FILLCELL_X2 FILLER_54_978 ();
 FILLCELL_X1 FILLER_54_980 ();
 FILLCELL_X4 FILLER_54_1015 ();
 FILLCELL_X1 FILLER_54_1019 ();
 FILLCELL_X4 FILLER_54_1024 ();
 FILLCELL_X2 FILLER_54_1028 ();
 FILLCELL_X1 FILLER_54_1030 ();
 FILLCELL_X8 FILLER_54_1037 ();
 FILLCELL_X4 FILLER_54_1049 ();
 FILLCELL_X8 FILLER_54_1063 ();
 FILLCELL_X4 FILLER_54_1071 ();
 FILLCELL_X2 FILLER_54_1097 ();
 FILLCELL_X2 FILLER_54_1108 ();
 FILLCELL_X1 FILLER_54_1110 ();
 FILLCELL_X8 FILLER_54_1130 ();
 FILLCELL_X4 FILLER_54_1146 ();
 FILLCELL_X2 FILLER_54_1161 ();
 FILLCELL_X1 FILLER_54_1163 ();
 FILLCELL_X4 FILLER_54_1167 ();
 FILLCELL_X1 FILLER_54_1171 ();
 FILLCELL_X8 FILLER_54_1179 ();
 FILLCELL_X4 FILLER_54_1187 ();
 FILLCELL_X2 FILLER_54_1191 ();
 FILLCELL_X8 FILLER_54_1224 ();
 FILLCELL_X2 FILLER_54_1232 ();
 FILLCELL_X1 FILLER_54_1234 ();
 FILLCELL_X4 FILLER_54_1255 ();
 FILLCELL_X2 FILLER_54_1259 ();
 FILLCELL_X1 FILLER_54_1261 ();
 FILLCELL_X4 FILLER_54_1299 ();
 FILLCELL_X2 FILLER_54_1303 ();
 FILLCELL_X1 FILLER_54_1305 ();
 FILLCELL_X4 FILLER_54_1326 ();
 FILLCELL_X2 FILLER_54_1330 ();
 FILLCELL_X8 FILLER_54_1339 ();
 FILLCELL_X4 FILLER_54_1354 ();
 FILLCELL_X1 FILLER_54_1358 ();
 FILLCELL_X8 FILLER_54_1386 ();
 FILLCELL_X2 FILLER_54_1394 ();
 FILLCELL_X1 FILLER_54_1396 ();
 FILLCELL_X4 FILLER_54_1417 ();
 FILLCELL_X2 FILLER_54_1421 ();
 FILLCELL_X1 FILLER_54_1443 ();
 FILLCELL_X2 FILLER_54_1451 ();
 FILLCELL_X1 FILLER_54_1453 ();
 FILLCELL_X1 FILLER_54_1468 ();
 FILLCELL_X2 FILLER_54_1476 ();
 FILLCELL_X2 FILLER_54_1483 ();
 FILLCELL_X2 FILLER_54_1488 ();
 FILLCELL_X4 FILLER_54_1498 ();
 FILLCELL_X1 FILLER_54_1502 ();
 FILLCELL_X1 FILLER_54_1510 ();
 FILLCELL_X1 FILLER_54_1515 ();
 FILLCELL_X1 FILLER_54_1520 ();
 FILLCELL_X2 FILLER_54_1532 ();
 FILLCELL_X4 FILLER_54_1543 ();
 FILLCELL_X2 FILLER_54_1557 ();
 FILLCELL_X1 FILLER_54_1585 ();
 FILLCELL_X1 FILLER_54_1589 ();
 FILLCELL_X2 FILLER_54_1593 ();
 FILLCELL_X1 FILLER_54_1599 ();
 FILLCELL_X2 FILLER_54_1604 ();
 FILLCELL_X4 FILLER_54_1610 ();
 FILLCELL_X2 FILLER_54_1614 ();
 FILLCELL_X1 FILLER_54_1619 ();
 FILLCELL_X16 FILLER_54_1631 ();
 FILLCELL_X4 FILLER_54_1647 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X8 FILLER_55_129 ();
 FILLCELL_X2 FILLER_55_137 ();
 FILLCELL_X1 FILLER_55_139 ();
 FILLCELL_X2 FILLER_55_147 ();
 FILLCELL_X1 FILLER_55_149 ();
 FILLCELL_X8 FILLER_55_185 ();
 FILLCELL_X4 FILLER_55_193 ();
 FILLCELL_X2 FILLER_55_242 ();
 FILLCELL_X4 FILLER_55_251 ();
 FILLCELL_X2 FILLER_55_255 ();
 FILLCELL_X1 FILLER_55_284 ();
 FILLCELL_X4 FILLER_55_292 ();
 FILLCELL_X1 FILLER_55_296 ();
 FILLCELL_X2 FILLER_55_324 ();
 FILLCELL_X1 FILLER_55_326 ();
 FILLCELL_X2 FILLER_55_337 ();
 FILLCELL_X1 FILLER_55_339 ();
 FILLCELL_X8 FILLER_55_367 ();
 FILLCELL_X2 FILLER_55_375 ();
 FILLCELL_X4 FILLER_55_427 ();
 FILLCELL_X2 FILLER_55_431 ();
 FILLCELL_X8 FILLER_55_444 ();
 FILLCELL_X4 FILLER_55_452 ();
 FILLCELL_X2 FILLER_55_456 ();
 FILLCELL_X4 FILLER_55_465 ();
 FILLCELL_X4 FILLER_55_474 ();
 FILLCELL_X2 FILLER_55_478 ();
 FILLCELL_X1 FILLER_55_480 ();
 FILLCELL_X2 FILLER_55_491 ();
 FILLCELL_X1 FILLER_55_493 ();
 FILLCELL_X4 FILLER_55_499 ();
 FILLCELL_X2 FILLER_55_503 ();
 FILLCELL_X1 FILLER_55_505 ();
 FILLCELL_X4 FILLER_55_512 ();
 FILLCELL_X1 FILLER_55_516 ();
 FILLCELL_X1 FILLER_55_544 ();
 FILLCELL_X4 FILLER_55_570 ();
 FILLCELL_X8 FILLER_55_585 ();
 FILLCELL_X4 FILLER_55_593 ();
 FILLCELL_X2 FILLER_55_597 ();
 FILLCELL_X1 FILLER_55_604 ();
 FILLCELL_X2 FILLER_55_610 ();
 FILLCELL_X1 FILLER_55_612 ();
 FILLCELL_X16 FILLER_55_630 ();
 FILLCELL_X4 FILLER_55_646 ();
 FILLCELL_X16 FILLER_55_657 ();
 FILLCELL_X1 FILLER_55_673 ();
 FILLCELL_X16 FILLER_55_681 ();
 FILLCELL_X8 FILLER_55_697 ();
 FILLCELL_X1 FILLER_55_705 ();
 FILLCELL_X2 FILLER_55_728 ();
 FILLCELL_X8 FILLER_55_766 ();
 FILLCELL_X4 FILLER_55_774 ();
 FILLCELL_X2 FILLER_55_798 ();
 FILLCELL_X1 FILLER_55_800 ();
 FILLCELL_X16 FILLER_55_814 ();
 FILLCELL_X1 FILLER_55_830 ();
 FILLCELL_X1 FILLER_55_836 ();
 FILLCELL_X8 FILLER_55_846 ();
 FILLCELL_X4 FILLER_55_854 ();
 FILLCELL_X4 FILLER_55_882 ();
 FILLCELL_X2 FILLER_55_886 ();
 FILLCELL_X2 FILLER_55_893 ();
 FILLCELL_X4 FILLER_55_908 ();
 FILLCELL_X2 FILLER_55_912 ();
 FILLCELL_X2 FILLER_55_931 ();
 FILLCELL_X1 FILLER_55_933 ();
 FILLCELL_X4 FILLER_55_936 ();
 FILLCELL_X1 FILLER_55_940 ();
 FILLCELL_X4 FILLER_55_945 ();
 FILLCELL_X2 FILLER_55_949 ();
 FILLCELL_X1 FILLER_55_984 ();
 FILLCELL_X2 FILLER_55_1011 ();
 FILLCELL_X1 FILLER_55_1026 ();
 FILLCELL_X2 FILLER_55_1045 ();
 FILLCELL_X1 FILLER_55_1060 ();
 FILLCELL_X1 FILLER_55_1085 ();
 FILLCELL_X1 FILLER_55_1097 ();
 FILLCELL_X1 FILLER_55_1129 ();
 FILLCELL_X8 FILLER_55_1144 ();
 FILLCELL_X8 FILLER_55_1176 ();
 FILLCELL_X4 FILLER_55_1184 ();
 FILLCELL_X32 FILLER_55_1191 ();
 FILLCELL_X4 FILLER_55_1237 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X4 FILLER_55_1271 ();
 FILLCELL_X2 FILLER_55_1275 ();
 FILLCELL_X1 FILLER_55_1277 ();
 FILLCELL_X1 FILLER_55_1281 ();
 FILLCELL_X1 FILLER_55_1292 ();
 FILLCELL_X4 FILLER_55_1345 ();
 FILLCELL_X1 FILLER_55_1349 ();
 FILLCELL_X2 FILLER_55_1360 ();
 FILLCELL_X1 FILLER_55_1362 ();
 FILLCELL_X8 FILLER_55_1366 ();
 FILLCELL_X2 FILLER_55_1374 ();
 FILLCELL_X16 FILLER_55_1383 ();
 FILLCELL_X4 FILLER_55_1399 ();
 FILLCELL_X2 FILLER_55_1403 ();
 FILLCELL_X1 FILLER_55_1405 ();
 FILLCELL_X1 FILLER_55_1418 ();
 FILLCELL_X8 FILLER_55_1430 ();
 FILLCELL_X4 FILLER_55_1447 ();
 FILLCELL_X1 FILLER_55_1451 ();
 FILLCELL_X8 FILLER_55_1457 ();
 FILLCELL_X4 FILLER_55_1465 ();
 FILLCELL_X1 FILLER_55_1469 ();
 FILLCELL_X1 FILLER_55_1495 ();
 FILLCELL_X1 FILLER_55_1501 ();
 FILLCELL_X1 FILLER_55_1517 ();
 FILLCELL_X8 FILLER_55_1522 ();
 FILLCELL_X4 FILLER_55_1530 ();
 FILLCELL_X16 FILLER_55_1538 ();
 FILLCELL_X4 FILLER_55_1554 ();
 FILLCELL_X4 FILLER_55_1576 ();
 FILLCELL_X1 FILLER_55_1580 ();
 FILLCELL_X2 FILLER_55_1586 ();
 FILLCELL_X1 FILLER_55_1588 ();
 FILLCELL_X4 FILLER_55_1593 ();
 FILLCELL_X2 FILLER_55_1597 ();
 FILLCELL_X8 FILLER_55_1603 ();
 FILLCELL_X4 FILLER_55_1611 ();
 FILLCELL_X1 FILLER_55_1615 ();
 FILLCELL_X1 FILLER_55_1620 ();
 FILLCELL_X16 FILLER_55_1625 ();
 FILLCELL_X8 FILLER_55_1641 ();
 FILLCELL_X2 FILLER_55_1649 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X8 FILLER_56_129 ();
 FILLCELL_X4 FILLER_56_137 ();
 FILLCELL_X4 FILLER_56_148 ();
 FILLCELL_X2 FILLER_56_152 ();
 FILLCELL_X1 FILLER_56_154 ();
 FILLCELL_X2 FILLER_56_162 ();
 FILLCELL_X1 FILLER_56_164 ();
 FILLCELL_X8 FILLER_56_185 ();
 FILLCELL_X2 FILLER_56_193 ();
 FILLCELL_X2 FILLER_56_215 ();
 FILLCELL_X1 FILLER_56_217 ();
 FILLCELL_X1 FILLER_56_235 ();
 FILLCELL_X16 FILLER_56_245 ();
 FILLCELL_X1 FILLER_56_261 ();
 FILLCELL_X4 FILLER_56_293 ();
 FILLCELL_X1 FILLER_56_297 ();
 FILLCELL_X8 FILLER_56_301 ();
 FILLCELL_X1 FILLER_56_309 ();
 FILLCELL_X2 FILLER_56_329 ();
 FILLCELL_X1 FILLER_56_331 ();
 FILLCELL_X8 FILLER_56_348 ();
 FILLCELL_X4 FILLER_56_356 ();
 FILLCELL_X1 FILLER_56_360 ();
 FILLCELL_X4 FILLER_56_367 ();
 FILLCELL_X8 FILLER_56_381 ();
 FILLCELL_X1 FILLER_56_389 ();
 FILLCELL_X4 FILLER_56_420 ();
 FILLCELL_X1 FILLER_56_424 ();
 FILLCELL_X2 FILLER_56_472 ();
 FILLCELL_X2 FILLER_56_478 ();
 FILLCELL_X1 FILLER_56_480 ();
 FILLCELL_X1 FILLER_56_490 ();
 FILLCELL_X1 FILLER_56_495 ();
 FILLCELL_X1 FILLER_56_500 ();
 FILLCELL_X1 FILLER_56_504 ();
 FILLCELL_X8 FILLER_56_511 ();
 FILLCELL_X2 FILLER_56_519 ();
 FILLCELL_X1 FILLER_56_521 ();
 FILLCELL_X2 FILLER_56_544 ();
 FILLCELL_X1 FILLER_56_551 ();
 FILLCELL_X1 FILLER_56_569 ();
 FILLCELL_X8 FILLER_56_580 ();
 FILLCELL_X4 FILLER_56_588 ();
 FILLCELL_X2 FILLER_56_592 ();
 FILLCELL_X4 FILLER_56_605 ();
 FILLCELL_X8 FILLER_56_619 ();
 FILLCELL_X1 FILLER_56_627 ();
 FILLCELL_X2 FILLER_56_632 ();
 FILLCELL_X2 FILLER_56_640 ();
 FILLCELL_X1 FILLER_56_642 ();
 FILLCELL_X4 FILLER_56_648 ();
 FILLCELL_X1 FILLER_56_652 ();
 FILLCELL_X8 FILLER_56_690 ();
 FILLCELL_X4 FILLER_56_702 ();
 FILLCELL_X2 FILLER_56_706 ();
 FILLCELL_X8 FILLER_56_714 ();
 FILLCELL_X2 FILLER_56_722 ();
 FILLCELL_X8 FILLER_56_735 ();
 FILLCELL_X2 FILLER_56_743 ();
 FILLCELL_X4 FILLER_56_749 ();
 FILLCELL_X2 FILLER_56_753 ();
 FILLCELL_X1 FILLER_56_755 ();
 FILLCELL_X2 FILLER_56_760 ();
 FILLCELL_X8 FILLER_56_767 ();
 FILLCELL_X4 FILLER_56_775 ();
 FILLCELL_X2 FILLER_56_779 ();
 FILLCELL_X1 FILLER_56_799 ();
 FILLCELL_X1 FILLER_56_816 ();
 FILLCELL_X8 FILLER_56_852 ();
 FILLCELL_X4 FILLER_56_864 ();
 FILLCELL_X1 FILLER_56_868 ();
 FILLCELL_X1 FILLER_56_887 ();
 FILLCELL_X2 FILLER_56_905 ();
 FILLCELL_X1 FILLER_56_907 ();
 FILLCELL_X4 FILLER_56_938 ();
 FILLCELL_X1 FILLER_56_942 ();
 FILLCELL_X4 FILLER_56_951 ();
 FILLCELL_X2 FILLER_56_984 ();
 FILLCELL_X8 FILLER_56_989 ();
 FILLCELL_X1 FILLER_56_997 ();
 FILLCELL_X2 FILLER_56_1028 ();
 FILLCELL_X1 FILLER_56_1030 ();
 FILLCELL_X4 FILLER_56_1037 ();
 FILLCELL_X1 FILLER_56_1041 ();
 FILLCELL_X4 FILLER_56_1045 ();
 FILLCELL_X1 FILLER_56_1049 ();
 FILLCELL_X1 FILLER_56_1059 ();
 FILLCELL_X4 FILLER_56_1063 ();
 FILLCELL_X1 FILLER_56_1067 ();
 FILLCELL_X4 FILLER_56_1084 ();
 FILLCELL_X1 FILLER_56_1088 ();
 FILLCELL_X1 FILLER_56_1092 ();
 FILLCELL_X2 FILLER_56_1100 ();
 FILLCELL_X4 FILLER_56_1108 ();
 FILLCELL_X4 FILLER_56_1118 ();
 FILLCELL_X2 FILLER_56_1122 ();
 FILLCELL_X1 FILLER_56_1124 ();
 FILLCELL_X1 FILLER_56_1166 ();
 FILLCELL_X1 FILLER_56_1187 ();
 FILLCELL_X8 FILLER_56_1198 ();
 FILLCELL_X4 FILLER_56_1206 ();
 FILLCELL_X1 FILLER_56_1210 ();
 FILLCELL_X8 FILLER_56_1225 ();
 FILLCELL_X2 FILLER_56_1233 ();
 FILLCELL_X4 FILLER_56_1247 ();
 FILLCELL_X1 FILLER_56_1251 ();
 FILLCELL_X2 FILLER_56_1259 ();
 FILLCELL_X4 FILLER_56_1268 ();
 FILLCELL_X1 FILLER_56_1272 ();
 FILLCELL_X1 FILLER_56_1287 ();
 FILLCELL_X2 FILLER_56_1306 ();
 FILLCELL_X1 FILLER_56_1321 ();
 FILLCELL_X2 FILLER_56_1342 ();
 FILLCELL_X2 FILLER_56_1351 ();
 FILLCELL_X1 FILLER_56_1353 ();
 FILLCELL_X1 FILLER_56_1357 ();
 FILLCELL_X16 FILLER_56_1385 ();
 FILLCELL_X8 FILLER_56_1401 ();
 FILLCELL_X1 FILLER_56_1413 ();
 FILLCELL_X1 FILLER_56_1425 ();
 FILLCELL_X2 FILLER_56_1444 ();
 FILLCELL_X2 FILLER_56_1455 ();
 FILLCELL_X1 FILLER_56_1457 ();
 FILLCELL_X4 FILLER_56_1468 ();
 FILLCELL_X1 FILLER_56_1472 ();
 FILLCELL_X8 FILLER_56_1493 ();
 FILLCELL_X1 FILLER_56_1501 ();
 FILLCELL_X1 FILLER_56_1506 ();
 FILLCELL_X1 FILLER_56_1511 ();
 FILLCELL_X1 FILLER_56_1517 ();
 FILLCELL_X2 FILLER_56_1527 ();
 FILLCELL_X1 FILLER_56_1529 ();
 FILLCELL_X2 FILLER_56_1538 ();
 FILLCELL_X2 FILLER_56_1550 ();
 FILLCELL_X1 FILLER_56_1552 ();
 FILLCELL_X8 FILLER_56_1557 ();
 FILLCELL_X1 FILLER_56_1568 ();
 FILLCELL_X4 FILLER_56_1584 ();
 FILLCELL_X2 FILLER_56_1601 ();
 FILLCELL_X32 FILLER_56_1614 ();
 FILLCELL_X4 FILLER_56_1646 ();
 FILLCELL_X1 FILLER_56_1650 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X4 FILLER_57_129 ();
 FILLCELL_X1 FILLER_57_133 ();
 FILLCELL_X4 FILLER_57_154 ();
 FILLCELL_X2 FILLER_57_158 ();
 FILLCELL_X1 FILLER_57_160 ();
 FILLCELL_X8 FILLER_57_175 ();
 FILLCELL_X2 FILLER_57_183 ();
 FILLCELL_X2 FILLER_57_192 ();
 FILLCELL_X1 FILLER_57_220 ();
 FILLCELL_X2 FILLER_57_234 ();
 FILLCELL_X2 FILLER_57_253 ();
 FILLCELL_X2 FILLER_57_309 ();
 FILLCELL_X8 FILLER_57_315 ();
 FILLCELL_X2 FILLER_57_323 ();
 FILLCELL_X1 FILLER_57_325 ();
 FILLCELL_X2 FILLER_57_339 ();
 FILLCELL_X1 FILLER_57_341 ();
 FILLCELL_X4 FILLER_57_346 ();
 FILLCELL_X1 FILLER_57_350 ();
 FILLCELL_X8 FILLER_57_381 ();
 FILLCELL_X2 FILLER_57_389 ();
 FILLCELL_X2 FILLER_57_403 ();
 FILLCELL_X16 FILLER_57_412 ();
 FILLCELL_X2 FILLER_57_444 ();
 FILLCELL_X1 FILLER_57_446 ();
 FILLCELL_X2 FILLER_57_453 ();
 FILLCELL_X2 FILLER_57_465 ();
 FILLCELL_X8 FILLER_57_470 ();
 FILLCELL_X4 FILLER_57_495 ();
 FILLCELL_X2 FILLER_57_499 ();
 FILLCELL_X1 FILLER_57_511 ();
 FILLCELL_X4 FILLER_57_521 ();
 FILLCELL_X2 FILLER_57_525 ();
 FILLCELL_X1 FILLER_57_527 ();
 FILLCELL_X1 FILLER_57_548 ();
 FILLCELL_X2 FILLER_57_553 ();
 FILLCELL_X2 FILLER_57_627 ();
 FILLCELL_X2 FILLER_57_652 ();
 FILLCELL_X2 FILLER_57_657 ();
 FILLCELL_X2 FILLER_57_668 ();
 FILLCELL_X2 FILLER_57_673 ();
 FILLCELL_X1 FILLER_57_675 ();
 FILLCELL_X1 FILLER_57_680 ();
 FILLCELL_X1 FILLER_57_701 ();
 FILLCELL_X4 FILLER_57_715 ();
 FILLCELL_X1 FILLER_57_728 ();
 FILLCELL_X1 FILLER_57_735 ();
 FILLCELL_X4 FILLER_57_747 ();
 FILLCELL_X2 FILLER_57_751 ();
 FILLCELL_X1 FILLER_57_753 ();
 FILLCELL_X8 FILLER_57_763 ();
 FILLCELL_X4 FILLER_57_771 ();
 FILLCELL_X2 FILLER_57_775 ();
 FILLCELL_X1 FILLER_57_777 ();
 FILLCELL_X2 FILLER_57_824 ();
 FILLCELL_X1 FILLER_57_838 ();
 FILLCELL_X16 FILLER_57_845 ();
 FILLCELL_X4 FILLER_57_861 ();
 FILLCELL_X2 FILLER_57_882 ();
 FILLCELL_X8 FILLER_57_904 ();
 FILLCELL_X8 FILLER_57_919 ();
 FILLCELL_X4 FILLER_57_927 ();
 FILLCELL_X2 FILLER_57_931 ();
 FILLCELL_X1 FILLER_57_933 ();
 FILLCELL_X4 FILLER_57_959 ();
 FILLCELL_X16 FILLER_57_999 ();
 FILLCELL_X1 FILLER_57_1015 ();
 FILLCELL_X8 FILLER_57_1023 ();
 FILLCELL_X2 FILLER_57_1038 ();
 FILLCELL_X1 FILLER_57_1057 ();
 FILLCELL_X16 FILLER_57_1078 ();
 FILLCELL_X8 FILLER_57_1094 ();
 FILLCELL_X2 FILLER_57_1109 ();
 FILLCELL_X2 FILLER_57_1137 ();
 FILLCELL_X8 FILLER_57_1143 ();
 FILLCELL_X8 FILLER_57_1155 ();
 FILLCELL_X1 FILLER_57_1172 ();
 FILLCELL_X1 FILLER_57_1200 ();
 FILLCELL_X1 FILLER_57_1206 ();
 FILLCELL_X4 FILLER_57_1246 ();
 FILLCELL_X2 FILLER_57_1250 ();
 FILLCELL_X4 FILLER_57_1259 ();
 FILLCELL_X2 FILLER_57_1283 ();
 FILLCELL_X2 FILLER_57_1298 ();
 FILLCELL_X1 FILLER_57_1300 ();
 FILLCELL_X2 FILLER_57_1327 ();
 FILLCELL_X4 FILLER_57_1336 ();
 FILLCELL_X1 FILLER_57_1340 ();
 FILLCELL_X4 FILLER_57_1354 ();
 FILLCELL_X1 FILLER_57_1358 ();
 FILLCELL_X2 FILLER_57_1366 ();
 FILLCELL_X16 FILLER_57_1385 ();
 FILLCELL_X4 FILLER_57_1419 ();
 FILLCELL_X2 FILLER_57_1432 ();
 FILLCELL_X4 FILLER_57_1452 ();
 FILLCELL_X1 FILLER_57_1487 ();
 FILLCELL_X1 FILLER_57_1497 ();
 FILLCELL_X1 FILLER_57_1503 ();
 FILLCELL_X1 FILLER_57_1507 ();
 FILLCELL_X2 FILLER_57_1513 ();
 FILLCELL_X2 FILLER_57_1537 ();
 FILLCELL_X2 FILLER_57_1554 ();
 FILLCELL_X1 FILLER_57_1571 ();
 FILLCELL_X4 FILLER_57_1577 ();
 FILLCELL_X1 FILLER_57_1581 ();
 FILLCELL_X2 FILLER_57_1586 ();
 FILLCELL_X1 FILLER_57_1588 ();
 FILLCELL_X2 FILLER_57_1617 ();
 FILLCELL_X16 FILLER_57_1623 ();
 FILLCELL_X8 FILLER_57_1639 ();
 FILLCELL_X4 FILLER_57_1647 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X4 FILLER_58_129 ();
 FILLCELL_X2 FILLER_58_133 ();
 FILLCELL_X1 FILLER_58_135 ();
 FILLCELL_X2 FILLER_58_150 ();
 FILLCELL_X4 FILLER_58_179 ();
 FILLCELL_X2 FILLER_58_183 ();
 FILLCELL_X1 FILLER_58_185 ();
 FILLCELL_X16 FILLER_58_193 ();
 FILLCELL_X2 FILLER_58_268 ();
 FILLCELL_X4 FILLER_58_274 ();
 FILLCELL_X8 FILLER_58_285 ();
 FILLCELL_X1 FILLER_58_293 ();
 FILLCELL_X2 FILLER_58_341 ();
 FILLCELL_X4 FILLER_58_346 ();
 FILLCELL_X2 FILLER_58_350 ();
 FILLCELL_X1 FILLER_58_355 ();
 FILLCELL_X1 FILLER_58_360 ();
 FILLCELL_X2 FILLER_58_365 ();
 FILLCELL_X2 FILLER_58_370 ();
 FILLCELL_X8 FILLER_58_396 ();
 FILLCELL_X2 FILLER_58_404 ();
 FILLCELL_X1 FILLER_58_416 ();
 FILLCELL_X4 FILLER_58_430 ();
 FILLCELL_X1 FILLER_58_438 ();
 FILLCELL_X2 FILLER_58_445 ();
 FILLCELL_X2 FILLER_58_453 ();
 FILLCELL_X2 FILLER_58_462 ();
 FILLCELL_X1 FILLER_58_464 ();
 FILLCELL_X4 FILLER_58_479 ();
 FILLCELL_X2 FILLER_58_518 ();
 FILLCELL_X1 FILLER_58_520 ();
 FILLCELL_X2 FILLER_58_527 ();
 FILLCELL_X1 FILLER_58_529 ();
 FILLCELL_X2 FILLER_58_536 ();
 FILLCELL_X1 FILLER_58_538 ();
 FILLCELL_X8 FILLER_58_552 ();
 FILLCELL_X2 FILLER_58_560 ();
 FILLCELL_X1 FILLER_58_562 ();
 FILLCELL_X1 FILLER_58_567 ();
 FILLCELL_X1 FILLER_58_572 ();
 FILLCELL_X8 FILLER_58_587 ();
 FILLCELL_X1 FILLER_58_595 ();
 FILLCELL_X8 FILLER_58_602 ();
 FILLCELL_X4 FILLER_58_610 ();
 FILLCELL_X1 FILLER_58_614 ();
 FILLCELL_X8 FILLER_58_622 ();
 FILLCELL_X1 FILLER_58_630 ();
 FILLCELL_X2 FILLER_58_650 ();
 FILLCELL_X4 FILLER_58_701 ();
 FILLCELL_X1 FILLER_58_716 ();
 FILLCELL_X1 FILLER_58_720 ();
 FILLCELL_X1 FILLER_58_725 ();
 FILLCELL_X1 FILLER_58_735 ();
 FILLCELL_X1 FILLER_58_743 ();
 FILLCELL_X2 FILLER_58_797 ();
 FILLCELL_X1 FILLER_58_799 ();
 FILLCELL_X8 FILLER_58_802 ();
 FILLCELL_X1 FILLER_58_810 ();
 FILLCELL_X1 FILLER_58_824 ();
 FILLCELL_X1 FILLER_58_842 ();
 FILLCELL_X2 FILLER_58_850 ();
 FILLCELL_X4 FILLER_58_881 ();
 FILLCELL_X1 FILLER_58_885 ();
 FILLCELL_X2 FILLER_58_893 ();
 FILLCELL_X1 FILLER_58_895 ();
 FILLCELL_X2 FILLER_58_900 ();
 FILLCELL_X8 FILLER_58_906 ();
 FILLCELL_X4 FILLER_58_914 ();
 FILLCELL_X1 FILLER_58_918 ();
 FILLCELL_X2 FILLER_58_934 ();
 FILLCELL_X1 FILLER_58_936 ();
 FILLCELL_X2 FILLER_58_946 ();
 FILLCELL_X1 FILLER_58_948 ();
 FILLCELL_X4 FILLER_58_954 ();
 FILLCELL_X1 FILLER_58_958 ();
 FILLCELL_X4 FILLER_58_964 ();
 FILLCELL_X2 FILLER_58_968 ();
 FILLCELL_X4 FILLER_58_972 ();
 FILLCELL_X1 FILLER_58_976 ();
 FILLCELL_X2 FILLER_58_995 ();
 FILLCELL_X1 FILLER_58_997 ();
 FILLCELL_X4 FILLER_58_1000 ();
 FILLCELL_X2 FILLER_58_1004 ();
 FILLCELL_X1 FILLER_58_1006 ();
 FILLCELL_X8 FILLER_58_1014 ();
 FILLCELL_X4 FILLER_58_1022 ();
 FILLCELL_X1 FILLER_58_1026 ();
 FILLCELL_X4 FILLER_58_1046 ();
 FILLCELL_X4 FILLER_58_1056 ();
 FILLCELL_X4 FILLER_58_1067 ();
 FILLCELL_X1 FILLER_58_1077 ();
 FILLCELL_X1 FILLER_58_1087 ();
 FILLCELL_X1 FILLER_58_1098 ();
 FILLCELL_X1 FILLER_58_1105 ();
 FILLCELL_X1 FILLER_58_1112 ();
 FILLCELL_X2 FILLER_58_1126 ();
 FILLCELL_X1 FILLER_58_1130 ();
 FILLCELL_X16 FILLER_58_1135 ();
 FILLCELL_X8 FILLER_58_1165 ();
 FILLCELL_X2 FILLER_58_1173 ();
 FILLCELL_X1 FILLER_58_1175 ();
 FILLCELL_X4 FILLER_58_1201 ();
 FILLCELL_X4 FILLER_58_1210 ();
 FILLCELL_X2 FILLER_58_1214 ();
 FILLCELL_X1 FILLER_58_1216 ();
 FILLCELL_X2 FILLER_58_1242 ();
 FILLCELL_X1 FILLER_58_1244 ();
 FILLCELL_X4 FILLER_58_1279 ();
 FILLCELL_X4 FILLER_58_1362 ();
 FILLCELL_X2 FILLER_58_1366 ();
 FILLCELL_X16 FILLER_58_1388 ();
 FILLCELL_X4 FILLER_58_1404 ();
 FILLCELL_X2 FILLER_58_1408 ();
 FILLCELL_X1 FILLER_58_1410 ();
 FILLCELL_X1 FILLER_58_1420 ();
 FILLCELL_X1 FILLER_58_1430 ();
 FILLCELL_X2 FILLER_58_1444 ();
 FILLCELL_X1 FILLER_58_1446 ();
 FILLCELL_X1 FILLER_58_1456 ();
 FILLCELL_X4 FILLER_58_1466 ();
 FILLCELL_X1 FILLER_58_1470 ();
 FILLCELL_X4 FILLER_58_1475 ();
 FILLCELL_X4 FILLER_58_1488 ();
 FILLCELL_X1 FILLER_58_1492 ();
 FILLCELL_X4 FILLER_58_1514 ();
 FILLCELL_X1 FILLER_58_1518 ();
 FILLCELL_X8 FILLER_58_1533 ();
 FILLCELL_X1 FILLER_58_1541 ();
 FILLCELL_X8 FILLER_58_1554 ();
 FILLCELL_X1 FILLER_58_1562 ();
 FILLCELL_X16 FILLER_58_1581 ();
 FILLCELL_X4 FILLER_58_1597 ();
 FILLCELL_X1 FILLER_58_1617 ();
 FILLCELL_X8 FILLER_58_1642 ();
 FILLCELL_X1 FILLER_58_1650 ();
 FILLCELL_X16 FILLER_59_1 ();
 FILLCELL_X2 FILLER_59_17 ();
 FILLCELL_X32 FILLER_59_22 ();
 FILLCELL_X32 FILLER_59_54 ();
 FILLCELL_X32 FILLER_59_86 ();
 FILLCELL_X8 FILLER_59_118 ();
 FILLCELL_X4 FILLER_59_126 ();
 FILLCELL_X2 FILLER_59_130 ();
 FILLCELL_X4 FILLER_59_160 ();
 FILLCELL_X1 FILLER_59_164 ();
 FILLCELL_X8 FILLER_59_172 ();
 FILLCELL_X4 FILLER_59_180 ();
 FILLCELL_X2 FILLER_59_184 ();
 FILLCELL_X1 FILLER_59_186 ();
 FILLCELL_X4 FILLER_59_216 ();
 FILLCELL_X1 FILLER_59_220 ();
 FILLCELL_X2 FILLER_59_224 ();
 FILLCELL_X1 FILLER_59_231 ();
 FILLCELL_X1 FILLER_59_243 ();
 FILLCELL_X1 FILLER_59_257 ();
 FILLCELL_X16 FILLER_59_269 ();
 FILLCELL_X8 FILLER_59_285 ();
 FILLCELL_X4 FILLER_59_293 ();
 FILLCELL_X2 FILLER_59_297 ();
 FILLCELL_X1 FILLER_59_313 ();
 FILLCELL_X8 FILLER_59_319 ();
 FILLCELL_X1 FILLER_59_327 ();
 FILLCELL_X2 FILLER_59_337 ();
 FILLCELL_X1 FILLER_59_339 ();
 FILLCELL_X8 FILLER_59_344 ();
 FILLCELL_X4 FILLER_59_352 ();
 FILLCELL_X2 FILLER_59_359 ();
 FILLCELL_X2 FILLER_59_378 ();
 FILLCELL_X8 FILLER_59_409 ();
 FILLCELL_X1 FILLER_59_428 ();
 FILLCELL_X8 FILLER_59_452 ();
 FILLCELL_X16 FILLER_59_463 ();
 FILLCELL_X4 FILLER_59_479 ();
 FILLCELL_X4 FILLER_59_489 ();
 FILLCELL_X2 FILLER_59_493 ();
 FILLCELL_X1 FILLER_59_495 ();
 FILLCELL_X4 FILLER_59_499 ();
 FILLCELL_X2 FILLER_59_523 ();
 FILLCELL_X1 FILLER_59_525 ();
 FILLCELL_X16 FILLER_59_537 ();
 FILLCELL_X2 FILLER_59_553 ();
 FILLCELL_X4 FILLER_59_558 ();
 FILLCELL_X1 FILLER_59_562 ();
 FILLCELL_X8 FILLER_59_608 ();
 FILLCELL_X4 FILLER_59_616 ();
 FILLCELL_X2 FILLER_59_620 ();
 FILLCELL_X1 FILLER_59_635 ();
 FILLCELL_X2 FILLER_59_645 ();
 FILLCELL_X2 FILLER_59_665 ();
 FILLCELL_X2 FILLER_59_675 ();
 FILLCELL_X1 FILLER_59_681 ();
 FILLCELL_X1 FILLER_59_686 ();
 FILLCELL_X1 FILLER_59_692 ();
 FILLCELL_X1 FILLER_59_697 ();
 FILLCELL_X2 FILLER_59_719 ();
 FILLCELL_X1 FILLER_59_721 ();
 FILLCELL_X1 FILLER_59_729 ();
 FILLCELL_X2 FILLER_59_743 ();
 FILLCELL_X2 FILLER_59_764 ();
 FILLCELL_X1 FILLER_59_766 ();
 FILLCELL_X8 FILLER_59_783 ();
 FILLCELL_X4 FILLER_59_791 ();
 FILLCELL_X2 FILLER_59_795 ();
 FILLCELL_X4 FILLER_59_828 ();
 FILLCELL_X16 FILLER_59_850 ();
 FILLCELL_X4 FILLER_59_866 ();
 FILLCELL_X2 FILLER_59_881 ();
 FILLCELL_X1 FILLER_59_883 ();
 FILLCELL_X4 FILLER_59_910 ();
 FILLCELL_X8 FILLER_59_916 ();
 FILLCELL_X4 FILLER_59_936 ();
 FILLCELL_X2 FILLER_59_945 ();
 FILLCELL_X1 FILLER_59_947 ();
 FILLCELL_X4 FILLER_59_973 ();
 FILLCELL_X8 FILLER_59_1027 ();
 FILLCELL_X2 FILLER_59_1048 ();
 FILLCELL_X1 FILLER_59_1050 ();
 FILLCELL_X2 FILLER_59_1089 ();
 FILLCELL_X2 FILLER_59_1113 ();
 FILLCELL_X1 FILLER_59_1115 ();
 FILLCELL_X8 FILLER_59_1122 ();
 FILLCELL_X1 FILLER_59_1130 ();
 FILLCELL_X1 FILLER_59_1135 ();
 FILLCELL_X16 FILLER_59_1177 ();
 FILLCELL_X4 FILLER_59_1193 ();
 FILLCELL_X1 FILLER_59_1197 ();
 FILLCELL_X8 FILLER_59_1202 ();
 FILLCELL_X4 FILLER_59_1210 ();
 FILLCELL_X2 FILLER_59_1214 ();
 FILLCELL_X1 FILLER_59_1216 ();
 FILLCELL_X2 FILLER_59_1224 ();
 FILLCELL_X1 FILLER_59_1226 ();
 FILLCELL_X4 FILLER_59_1234 ();
 FILLCELL_X16 FILLER_59_1245 ();
 FILLCELL_X2 FILLER_59_1261 ();
 FILLCELL_X8 FILLER_59_1284 ();
 FILLCELL_X4 FILLER_59_1292 ();
 FILLCELL_X8 FILLER_59_1337 ();
 FILLCELL_X1 FILLER_59_1345 ();
 FILLCELL_X1 FILLER_59_1366 ();
 FILLCELL_X16 FILLER_59_1374 ();
 FILLCELL_X8 FILLER_59_1399 ();
 FILLCELL_X4 FILLER_59_1407 ();
 FILLCELL_X2 FILLER_59_1418 ();
 FILLCELL_X1 FILLER_59_1420 ();
 FILLCELL_X2 FILLER_59_1447 ();
 FILLCELL_X2 FILLER_59_1460 ();
 FILLCELL_X2 FILLER_59_1471 ();
 FILLCELL_X4 FILLER_59_1477 ();
 FILLCELL_X2 FILLER_59_1490 ();
 FILLCELL_X4 FILLER_59_1501 ();
 FILLCELL_X8 FILLER_59_1517 ();
 FILLCELL_X4 FILLER_59_1525 ();
 FILLCELL_X1 FILLER_59_1529 ();
 FILLCELL_X1 FILLER_59_1541 ();
 FILLCELL_X16 FILLER_59_1546 ();
 FILLCELL_X4 FILLER_59_1562 ();
 FILLCELL_X4 FILLER_59_1577 ();
 FILLCELL_X2 FILLER_59_1581 ();
 FILLCELL_X1 FILLER_59_1583 ();
 FILLCELL_X8 FILLER_59_1587 ();
 FILLCELL_X2 FILLER_59_1595 ();
 FILLCELL_X4 FILLER_59_1611 ();
 FILLCELL_X1 FILLER_59_1624 ();
 FILLCELL_X16 FILLER_59_1632 ();
 FILLCELL_X2 FILLER_59_1648 ();
 FILLCELL_X1 FILLER_59_1650 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X16 FILLER_60_97 ();
 FILLCELL_X8 FILLER_60_113 ();
 FILLCELL_X4 FILLER_60_121 ();
 FILLCELL_X2 FILLER_60_125 ();
 FILLCELL_X2 FILLER_60_154 ();
 FILLCELL_X2 FILLER_60_183 ();
 FILLCELL_X4 FILLER_60_222 ();
 FILLCELL_X2 FILLER_60_242 ();
 FILLCELL_X1 FILLER_60_244 ();
 FILLCELL_X4 FILLER_60_270 ();
 FILLCELL_X1 FILLER_60_274 ();
 FILLCELL_X8 FILLER_60_284 ();
 FILLCELL_X2 FILLER_60_297 ();
 FILLCELL_X1 FILLER_60_299 ();
 FILLCELL_X1 FILLER_60_305 ();
 FILLCELL_X1 FILLER_60_310 ();
 FILLCELL_X1 FILLER_60_324 ();
 FILLCELL_X2 FILLER_60_373 ();
 FILLCELL_X1 FILLER_60_375 ();
 FILLCELL_X16 FILLER_60_393 ();
 FILLCELL_X4 FILLER_60_409 ();
 FILLCELL_X2 FILLER_60_413 ();
 FILLCELL_X1 FILLER_60_415 ();
 FILLCELL_X1 FILLER_60_440 ();
 FILLCELL_X1 FILLER_60_447 ();
 FILLCELL_X4 FILLER_60_453 ();
 FILLCELL_X2 FILLER_60_457 ();
 FILLCELL_X4 FILLER_60_481 ();
 FILLCELL_X4 FILLER_60_501 ();
 FILLCELL_X1 FILLER_60_505 ();
 FILLCELL_X4 FILLER_60_511 ();
 FILLCELL_X2 FILLER_60_515 ();
 FILLCELL_X2 FILLER_60_524 ();
 FILLCELL_X8 FILLER_60_533 ();
 FILLCELL_X1 FILLER_60_541 ();
 FILLCELL_X32 FILLER_60_562 ();
 FILLCELL_X1 FILLER_60_594 ();
 FILLCELL_X2 FILLER_60_608 ();
 FILLCELL_X1 FILLER_60_610 ();
 FILLCELL_X1 FILLER_60_632 ();
 FILLCELL_X2 FILLER_60_643 ();
 FILLCELL_X2 FILLER_60_658 ();
 FILLCELL_X2 FILLER_60_664 ();
 FILLCELL_X1 FILLER_60_666 ();
 FILLCELL_X4 FILLER_60_674 ();
 FILLCELL_X1 FILLER_60_678 ();
 FILLCELL_X4 FILLER_60_700 ();
 FILLCELL_X2 FILLER_60_704 ();
 FILLCELL_X2 FILLER_60_722 ();
 FILLCELL_X1 FILLER_60_732 ();
 FILLCELL_X4 FILLER_60_780 ();
 FILLCELL_X2 FILLER_60_788 ();
 FILLCELL_X1 FILLER_60_790 ();
 FILLCELL_X8 FILLER_60_815 ();
 FILLCELL_X2 FILLER_60_840 ();
 FILLCELL_X2 FILLER_60_872 ();
 FILLCELL_X8 FILLER_60_880 ();
 FILLCELL_X1 FILLER_60_888 ();
 FILLCELL_X4 FILLER_60_894 ();
 FILLCELL_X2 FILLER_60_898 ();
 FILLCELL_X1 FILLER_60_900 ();
 FILLCELL_X4 FILLER_60_951 ();
 FILLCELL_X2 FILLER_60_967 ();
 FILLCELL_X1 FILLER_60_975 ();
 FILLCELL_X2 FILLER_60_978 ();
 FILLCELL_X1 FILLER_60_980 ();
 FILLCELL_X4 FILLER_60_996 ();
 FILLCELL_X1 FILLER_60_1000 ();
 FILLCELL_X1 FILLER_60_1020 ();
 FILLCELL_X2 FILLER_60_1044 ();
 FILLCELL_X2 FILLER_60_1058 ();
 FILLCELL_X1 FILLER_60_1060 ();
 FILLCELL_X2 FILLER_60_1066 ();
 FILLCELL_X2 FILLER_60_1084 ();
 FILLCELL_X4 FILLER_60_1092 ();
 FILLCELL_X2 FILLER_60_1096 ();
 FILLCELL_X2 FILLER_60_1110 ();
 FILLCELL_X1 FILLER_60_1112 ();
 FILLCELL_X1 FILLER_60_1115 ();
 FILLCELL_X1 FILLER_60_1123 ();
 FILLCELL_X1 FILLER_60_1128 ();
 FILLCELL_X4 FILLER_60_1135 ();
 FILLCELL_X8 FILLER_60_1167 ();
 FILLCELL_X4 FILLER_60_1175 ();
 FILLCELL_X2 FILLER_60_1179 ();
 FILLCELL_X1 FILLER_60_1201 ();
 FILLCELL_X2 FILLER_60_1229 ();
 FILLCELL_X1 FILLER_60_1231 ();
 FILLCELL_X8 FILLER_60_1239 ();
 FILLCELL_X2 FILLER_60_1247 ();
 FILLCELL_X16 FILLER_60_1269 ();
 FILLCELL_X2 FILLER_60_1285 ();
 FILLCELL_X1 FILLER_60_1290 ();
 FILLCELL_X2 FILLER_60_1303 ();
 FILLCELL_X1 FILLER_60_1305 ();
 FILLCELL_X4 FILLER_60_1313 ();
 FILLCELL_X1 FILLER_60_1317 ();
 FILLCELL_X2 FILLER_60_1325 ();
 FILLCELL_X2 FILLER_60_1334 ();
 FILLCELL_X1 FILLER_60_1336 ();
 FILLCELL_X2 FILLER_60_1357 ();
 FILLCELL_X1 FILLER_60_1359 ();
 FILLCELL_X16 FILLER_60_1377 ();
 FILLCELL_X1 FILLER_60_1429 ();
 FILLCELL_X4 FILLER_60_1442 ();
 FILLCELL_X1 FILLER_60_1446 ();
 FILLCELL_X4 FILLER_60_1451 ();
 FILLCELL_X4 FILLER_60_1459 ();
 FILLCELL_X1 FILLER_60_1463 ();
 FILLCELL_X8 FILLER_60_1492 ();
 FILLCELL_X1 FILLER_60_1505 ();
 FILLCELL_X1 FILLER_60_1509 ();
 FILLCELL_X2 FILLER_60_1513 ();
 FILLCELL_X2 FILLER_60_1522 ();
 FILLCELL_X2 FILLER_60_1528 ();
 FILLCELL_X2 FILLER_60_1538 ();
 FILLCELL_X2 FILLER_60_1544 ();
 FILLCELL_X4 FILLER_60_1562 ();
 FILLCELL_X4 FILLER_60_1569 ();
 FILLCELL_X2 FILLER_60_1573 ();
 FILLCELL_X1 FILLER_60_1575 ();
 FILLCELL_X4 FILLER_60_1579 ();
 FILLCELL_X2 FILLER_60_1583 ();
 FILLCELL_X1 FILLER_60_1585 ();
 FILLCELL_X8 FILLER_60_1591 ();
 FILLCELL_X2 FILLER_60_1599 ();
 FILLCELL_X1 FILLER_60_1601 ();
 FILLCELL_X2 FILLER_60_1606 ();
 FILLCELL_X4 FILLER_60_1626 ();
 FILLCELL_X2 FILLER_60_1630 ();
 FILLCELL_X16 FILLER_60_1635 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X4 FILLER_61_129 ();
 FILLCELL_X2 FILLER_61_133 ();
 FILLCELL_X1 FILLER_61_135 ();
 FILLCELL_X32 FILLER_61_143 ();
 FILLCELL_X4 FILLER_61_175 ();
 FILLCELL_X2 FILLER_61_213 ();
 FILLCELL_X1 FILLER_61_215 ();
 FILLCELL_X1 FILLER_61_223 ();
 FILLCELL_X1 FILLER_61_228 ();
 FILLCELL_X1 FILLER_61_249 ();
 FILLCELL_X1 FILLER_61_254 ();
 FILLCELL_X1 FILLER_61_258 ();
 FILLCELL_X1 FILLER_61_263 ();
 FILLCELL_X1 FILLER_61_284 ();
 FILLCELL_X8 FILLER_61_320 ();
 FILLCELL_X2 FILLER_61_328 ();
 FILLCELL_X1 FILLER_61_330 ();
 FILLCELL_X1 FILLER_61_333 ();
 FILLCELL_X1 FILLER_61_345 ();
 FILLCELL_X16 FILLER_61_361 ();
 FILLCELL_X1 FILLER_61_377 ();
 FILLCELL_X1 FILLER_61_385 ();
 FILLCELL_X2 FILLER_61_395 ();
 FILLCELL_X2 FILLER_61_404 ();
 FILLCELL_X4 FILLER_61_430 ();
 FILLCELL_X1 FILLER_61_434 ();
 FILLCELL_X16 FILLER_61_444 ();
 FILLCELL_X4 FILLER_61_460 ();
 FILLCELL_X2 FILLER_61_464 ();
 FILLCELL_X1 FILLER_61_466 ();
 FILLCELL_X1 FILLER_61_501 ();
 FILLCELL_X8 FILLER_61_547 ();
 FILLCELL_X4 FILLER_61_555 ();
 FILLCELL_X2 FILLER_61_559 ();
 FILLCELL_X1 FILLER_61_561 ();
 FILLCELL_X8 FILLER_61_570 ();
 FILLCELL_X2 FILLER_61_578 ();
 FILLCELL_X1 FILLER_61_580 ();
 FILLCELL_X8 FILLER_61_584 ();
 FILLCELL_X4 FILLER_61_592 ();
 FILLCELL_X1 FILLER_61_596 ();
 FILLCELL_X2 FILLER_61_604 ();
 FILLCELL_X1 FILLER_61_606 ();
 FILLCELL_X1 FILLER_61_618 ();
 FILLCELL_X4 FILLER_61_624 ();
 FILLCELL_X2 FILLER_61_628 ();
 FILLCELL_X1 FILLER_61_630 ();
 FILLCELL_X2 FILLER_61_642 ();
 FILLCELL_X8 FILLER_61_649 ();
 FILLCELL_X2 FILLER_61_657 ();
 FILLCELL_X1 FILLER_61_659 ();
 FILLCELL_X4 FILLER_61_681 ();
 FILLCELL_X1 FILLER_61_685 ();
 FILLCELL_X2 FILLER_61_696 ();
 FILLCELL_X1 FILLER_61_698 ();
 FILLCELL_X4 FILLER_61_706 ();
 FILLCELL_X2 FILLER_61_710 ();
 FILLCELL_X4 FILLER_61_715 ();
 FILLCELL_X1 FILLER_61_719 ();
 FILLCELL_X4 FILLER_61_736 ();
 FILLCELL_X2 FILLER_61_740 ();
 FILLCELL_X1 FILLER_61_742 ();
 FILLCELL_X4 FILLER_61_748 ();
 FILLCELL_X8 FILLER_61_759 ();
 FILLCELL_X2 FILLER_61_767 ();
 FILLCELL_X1 FILLER_61_769 ();
 FILLCELL_X2 FILLER_61_781 ();
 FILLCELL_X2 FILLER_61_809 ();
 FILLCELL_X16 FILLER_61_820 ();
 FILLCELL_X8 FILLER_61_836 ();
 FILLCELL_X1 FILLER_61_844 ();
 FILLCELL_X4 FILLER_61_850 ();
 FILLCELL_X1 FILLER_61_854 ();
 FILLCELL_X1 FILLER_61_892 ();
 FILLCELL_X16 FILLER_61_918 ();
 FILLCELL_X4 FILLER_61_934 ();
 FILLCELL_X2 FILLER_61_938 ();
 FILLCELL_X1 FILLER_61_940 ();
 FILLCELL_X4 FILLER_61_947 ();
 FILLCELL_X2 FILLER_61_958 ();
 FILLCELL_X1 FILLER_61_960 ();
 FILLCELL_X4 FILLER_61_993 ();
 FILLCELL_X8 FILLER_61_1010 ();
 FILLCELL_X4 FILLER_61_1018 ();
 FILLCELL_X2 FILLER_61_1022 ();
 FILLCELL_X1 FILLER_61_1024 ();
 FILLCELL_X8 FILLER_61_1030 ();
 FILLCELL_X2 FILLER_61_1049 ();
 FILLCELL_X2 FILLER_61_1057 ();
 FILLCELL_X8 FILLER_61_1069 ();
 FILLCELL_X2 FILLER_61_1077 ();
 FILLCELL_X1 FILLER_61_1086 ();
 FILLCELL_X8 FILLER_61_1091 ();
 FILLCELL_X1 FILLER_61_1106 ();
 FILLCELL_X2 FILLER_61_1124 ();
 FILLCELL_X1 FILLER_61_1126 ();
 FILLCELL_X1 FILLER_61_1130 ();
 FILLCELL_X2 FILLER_61_1134 ();
 FILLCELL_X1 FILLER_61_1136 ();
 FILLCELL_X2 FILLER_61_1171 ();
 FILLCELL_X16 FILLER_61_1187 ();
 FILLCELL_X4 FILLER_61_1203 ();
 FILLCELL_X1 FILLER_61_1227 ();
 FILLCELL_X2 FILLER_61_1235 ();
 FILLCELL_X1 FILLER_61_1262 ();
 FILLCELL_X2 FILLER_61_1293 ();
 FILLCELL_X2 FILLER_61_1304 ();
 FILLCELL_X1 FILLER_61_1306 ();
 FILLCELL_X1 FILLER_61_1314 ();
 FILLCELL_X2 FILLER_61_1322 ();
 FILLCELL_X1 FILLER_61_1324 ();
 FILLCELL_X1 FILLER_61_1352 ();
 FILLCELL_X1 FILLER_61_1368 ();
 FILLCELL_X16 FILLER_61_1376 ();
 FILLCELL_X2 FILLER_61_1392 ();
 FILLCELL_X1 FILLER_61_1420 ();
 FILLCELL_X4 FILLER_61_1439 ();
 FILLCELL_X1 FILLER_61_1443 ();
 FILLCELL_X2 FILLER_61_1448 ();
 FILLCELL_X1 FILLER_61_1450 ();
 FILLCELL_X8 FILLER_61_1465 ();
 FILLCELL_X4 FILLER_61_1473 ();
 FILLCELL_X2 FILLER_61_1480 ();
 FILLCELL_X1 FILLER_61_1482 ();
 FILLCELL_X8 FILLER_61_1491 ();
 FILLCELL_X4 FILLER_61_1499 ();
 FILLCELL_X2 FILLER_61_1503 ();
 FILLCELL_X1 FILLER_61_1505 ();
 FILLCELL_X2 FILLER_61_1513 ();
 FILLCELL_X1 FILLER_61_1515 ();
 FILLCELL_X1 FILLER_61_1539 ();
 FILLCELL_X1 FILLER_61_1543 ();
 FILLCELL_X2 FILLER_61_1555 ();
 FILLCELL_X1 FILLER_61_1573 ();
 FILLCELL_X2 FILLER_61_1578 ();
 FILLCELL_X2 FILLER_61_1584 ();
 FILLCELL_X1 FILLER_61_1590 ();
 FILLCELL_X2 FILLER_61_1595 ();
 FILLCELL_X1 FILLER_61_1612 ();
 FILLCELL_X2 FILLER_61_1622 ();
 FILLCELL_X16 FILLER_61_1631 ();
 FILLCELL_X4 FILLER_61_1647 ();
 FILLCELL_X8 FILLER_62_1 ();
 FILLCELL_X4 FILLER_62_9 ();
 FILLCELL_X32 FILLER_62_16 ();
 FILLCELL_X32 FILLER_62_48 ();
 FILLCELL_X32 FILLER_62_80 ();
 FILLCELL_X16 FILLER_62_112 ();
 FILLCELL_X8 FILLER_62_128 ();
 FILLCELL_X1 FILLER_62_136 ();
 FILLCELL_X1 FILLER_62_204 ();
 FILLCELL_X2 FILLER_62_208 ();
 FILLCELL_X8 FILLER_62_231 ();
 FILLCELL_X4 FILLER_62_239 ();
 FILLCELL_X2 FILLER_62_243 ();
 FILLCELL_X2 FILLER_62_271 ();
 FILLCELL_X1 FILLER_62_273 ();
 FILLCELL_X4 FILLER_62_308 ();
 FILLCELL_X2 FILLER_62_312 ();
 FILLCELL_X4 FILLER_62_334 ();
 FILLCELL_X2 FILLER_62_350 ();
 FILLCELL_X16 FILLER_62_355 ();
 FILLCELL_X4 FILLER_62_371 ();
 FILLCELL_X1 FILLER_62_405 ();
 FILLCELL_X4 FILLER_62_415 ();
 FILLCELL_X1 FILLER_62_419 ();
 FILLCELL_X16 FILLER_62_429 ();
 FILLCELL_X2 FILLER_62_445 ();
 FILLCELL_X16 FILLER_62_451 ();
 FILLCELL_X1 FILLER_62_467 ();
 FILLCELL_X2 FILLER_62_501 ();
 FILLCELL_X2 FILLER_62_513 ();
 FILLCELL_X1 FILLER_62_558 ();
 FILLCELL_X2 FILLER_62_568 ();
 FILLCELL_X2 FILLER_62_573 ();
 FILLCELL_X2 FILLER_62_578 ();
 FILLCELL_X1 FILLER_62_580 ();
 FILLCELL_X2 FILLER_62_594 ();
 FILLCELL_X1 FILLER_62_596 ();
 FILLCELL_X4 FILLER_62_600 ();
 FILLCELL_X2 FILLER_62_604 ();
 FILLCELL_X1 FILLER_62_606 ();
 FILLCELL_X4 FILLER_62_611 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X16 FILLER_62_632 ();
 FILLCELL_X4 FILLER_62_648 ();
 FILLCELL_X4 FILLER_62_655 ();
 FILLCELL_X1 FILLER_62_659 ();
 FILLCELL_X2 FILLER_62_663 ();
 FILLCELL_X1 FILLER_62_665 ();
 FILLCELL_X1 FILLER_62_675 ();
 FILLCELL_X4 FILLER_62_680 ();
 FILLCELL_X2 FILLER_62_684 ();
 FILLCELL_X1 FILLER_62_686 ();
 FILLCELL_X4 FILLER_62_704 ();
 FILLCELL_X4 FILLER_62_712 ();
 FILLCELL_X1 FILLER_62_716 ();
 FILLCELL_X4 FILLER_62_724 ();
 FILLCELL_X2 FILLER_62_728 ();
 FILLCELL_X8 FILLER_62_740 ();
 FILLCELL_X4 FILLER_62_755 ();
 FILLCELL_X1 FILLER_62_759 ();
 FILLCELL_X2 FILLER_62_773 ();
 FILLCELL_X1 FILLER_62_783 ();
 FILLCELL_X2 FILLER_62_792 ();
 FILLCELL_X1 FILLER_62_798 ();
 FILLCELL_X2 FILLER_62_812 ();
 FILLCELL_X8 FILLER_62_821 ();
 FILLCELL_X4 FILLER_62_829 ();
 FILLCELL_X2 FILLER_62_833 ();
 FILLCELL_X16 FILLER_62_840 ();
 FILLCELL_X2 FILLER_62_856 ();
 FILLCELL_X1 FILLER_62_879 ();
 FILLCELL_X1 FILLER_62_883 ();
 FILLCELL_X16 FILLER_62_912 ();
 FILLCELL_X1 FILLER_62_928 ();
 FILLCELL_X1 FILLER_62_934 ();
 FILLCELL_X4 FILLER_62_937 ();
 FILLCELL_X2 FILLER_62_941 ();
 FILLCELL_X1 FILLER_62_943 ();
 FILLCELL_X8 FILLER_62_950 ();
 FILLCELL_X2 FILLER_62_958 ();
 FILLCELL_X1 FILLER_62_967 ();
 FILLCELL_X4 FILLER_62_973 ();
 FILLCELL_X1 FILLER_62_977 ();
 FILLCELL_X4 FILLER_62_983 ();
 FILLCELL_X2 FILLER_62_987 ();
 FILLCELL_X1 FILLER_62_989 ();
 FILLCELL_X4 FILLER_62_999 ();
 FILLCELL_X2 FILLER_62_1003 ();
 FILLCELL_X1 FILLER_62_1005 ();
 FILLCELL_X16 FILLER_62_1009 ();
 FILLCELL_X4 FILLER_62_1025 ();
 FILLCELL_X1 FILLER_62_1029 ();
 FILLCELL_X2 FILLER_62_1032 ();
 FILLCELL_X4 FILLER_62_1041 ();
 FILLCELL_X2 FILLER_62_1065 ();
 FILLCELL_X1 FILLER_62_1096 ();
 FILLCELL_X8 FILLER_62_1104 ();
 FILLCELL_X2 FILLER_62_1112 ();
 FILLCELL_X1 FILLER_62_1114 ();
 FILLCELL_X2 FILLER_62_1118 ();
 FILLCELL_X1 FILLER_62_1128 ();
 FILLCELL_X1 FILLER_62_1154 ();
 FILLCELL_X2 FILLER_62_1174 ();
 FILLCELL_X1 FILLER_62_1176 ();
 FILLCELL_X4 FILLER_62_1199 ();
 FILLCELL_X8 FILLER_62_1210 ();
 FILLCELL_X4 FILLER_62_1218 ();
 FILLCELL_X2 FILLER_62_1222 ();
 FILLCELL_X1 FILLER_62_1224 ();
 FILLCELL_X1 FILLER_62_1305 ();
 FILLCELL_X1 FILLER_62_1309 ();
 FILLCELL_X8 FILLER_62_1317 ();
 FILLCELL_X1 FILLER_62_1325 ();
 FILLCELL_X2 FILLER_62_1333 ();
 FILLCELL_X8 FILLER_62_1382 ();
 FILLCELL_X4 FILLER_62_1401 ();
 FILLCELL_X2 FILLER_62_1405 ();
 FILLCELL_X2 FILLER_62_1416 ();
 FILLCELL_X1 FILLER_62_1418 ();
 FILLCELL_X2 FILLER_62_1432 ();
 FILLCELL_X2 FILLER_62_1441 ();
 FILLCELL_X1 FILLER_62_1443 ();
 FILLCELL_X4 FILLER_62_1449 ();
 FILLCELL_X2 FILLER_62_1466 ();
 FILLCELL_X1 FILLER_62_1476 ();
 FILLCELL_X4 FILLER_62_1486 ();
 FILLCELL_X8 FILLER_62_1508 ();
 FILLCELL_X2 FILLER_62_1516 ();
 FILLCELL_X4 FILLER_62_1520 ();
 FILLCELL_X2 FILLER_62_1524 ();
 FILLCELL_X8 FILLER_62_1537 ();
 FILLCELL_X2 FILLER_62_1545 ();
 FILLCELL_X4 FILLER_62_1555 ();
 FILLCELL_X1 FILLER_62_1559 ();
 FILLCELL_X2 FILLER_62_1567 ();
 FILLCELL_X2 FILLER_62_1572 ();
 FILLCELL_X1 FILLER_62_1574 ();
 FILLCELL_X1 FILLER_62_1579 ();
 FILLCELL_X1 FILLER_62_1589 ();
 FILLCELL_X2 FILLER_62_1601 ();
 FILLCELL_X2 FILLER_62_1606 ();
 FILLCELL_X4 FILLER_62_1612 ();
 FILLCELL_X4 FILLER_62_1620 ();
 FILLCELL_X16 FILLER_62_1629 ();
 FILLCELL_X4 FILLER_62_1645 ();
 FILLCELL_X2 FILLER_62_1649 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X8 FILLER_63_129 ();
 FILLCELL_X4 FILLER_63_157 ();
 FILLCELL_X2 FILLER_63_161 ();
 FILLCELL_X4 FILLER_63_170 ();
 FILLCELL_X2 FILLER_63_174 ();
 FILLCELL_X4 FILLER_63_196 ();
 FILLCELL_X2 FILLER_63_200 ();
 FILLCELL_X8 FILLER_63_217 ();
 FILLCELL_X4 FILLER_63_225 ();
 FILLCELL_X4 FILLER_63_241 ();
 FILLCELL_X1 FILLER_63_258 ();
 FILLCELL_X4 FILLER_63_268 ();
 FILLCELL_X1 FILLER_63_272 ();
 FILLCELL_X8 FILLER_63_277 ();
 FILLCELL_X1 FILLER_63_285 ();
 FILLCELL_X1 FILLER_63_311 ();
 FILLCELL_X4 FILLER_63_316 ();
 FILLCELL_X2 FILLER_63_320 ();
 FILLCELL_X2 FILLER_63_329 ();
 FILLCELL_X1 FILLER_63_334 ();
 FILLCELL_X1 FILLER_63_338 ();
 FILLCELL_X1 FILLER_63_365 ();
 FILLCELL_X2 FILLER_63_372 ();
 FILLCELL_X1 FILLER_63_392 ();
 FILLCELL_X8 FILLER_63_423 ();
 FILLCELL_X4 FILLER_63_431 ();
 FILLCELL_X8 FILLER_63_459 ();
 FILLCELL_X2 FILLER_63_467 ();
 FILLCELL_X2 FILLER_63_480 ();
 FILLCELL_X1 FILLER_63_482 ();
 FILLCELL_X8 FILLER_63_503 ();
 FILLCELL_X4 FILLER_63_511 ();
 FILLCELL_X1 FILLER_63_515 ();
 FILLCELL_X1 FILLER_63_533 ();
 FILLCELL_X8 FILLER_63_554 ();
 FILLCELL_X4 FILLER_63_562 ();
 FILLCELL_X4 FILLER_63_589 ();
 FILLCELL_X1 FILLER_63_617 ();
 FILLCELL_X2 FILLER_63_653 ();
 FILLCELL_X1 FILLER_63_666 ();
 FILLCELL_X1 FILLER_63_678 ();
 FILLCELL_X1 FILLER_63_683 ();
 FILLCELL_X4 FILLER_63_694 ();
 FILLCELL_X1 FILLER_63_714 ();
 FILLCELL_X1 FILLER_63_719 ();
 FILLCELL_X1 FILLER_63_724 ();
 FILLCELL_X1 FILLER_63_728 ();
 FILLCELL_X1 FILLER_63_736 ();
 FILLCELL_X4 FILLER_63_769 ();
 FILLCELL_X16 FILLER_63_808 ();
 FILLCELL_X8 FILLER_63_824 ();
 FILLCELL_X2 FILLER_63_832 ();
 FILLCELL_X2 FILLER_63_838 ();
 FILLCELL_X1 FILLER_63_840 ();
 FILLCELL_X16 FILLER_63_882 ();
 FILLCELL_X2 FILLER_63_898 ();
 FILLCELL_X2 FILLER_63_943 ();
 FILLCELL_X2 FILLER_63_996 ();
 FILLCELL_X1 FILLER_63_998 ();
 FILLCELL_X2 FILLER_63_1003 ();
 FILLCELL_X1 FILLER_63_1005 ();
 FILLCELL_X2 FILLER_63_1009 ();
 FILLCELL_X1 FILLER_63_1011 ();
 FILLCELL_X4 FILLER_63_1021 ();
 FILLCELL_X2 FILLER_63_1025 ();
 FILLCELL_X4 FILLER_63_1059 ();
 FILLCELL_X2 FILLER_63_1063 ();
 FILLCELL_X1 FILLER_63_1067 ();
 FILLCELL_X1 FILLER_63_1073 ();
 FILLCELL_X1 FILLER_63_1081 ();
 FILLCELL_X1 FILLER_63_1084 ();
 FILLCELL_X2 FILLER_63_1095 ();
 FILLCELL_X8 FILLER_63_1104 ();
 FILLCELL_X2 FILLER_63_1112 ();
 FILLCELL_X1 FILLER_63_1114 ();
 FILLCELL_X8 FILLER_63_1123 ();
 FILLCELL_X4 FILLER_63_1131 ();
 FILLCELL_X2 FILLER_63_1135 ();
 FILLCELL_X1 FILLER_63_1167 ();
 FILLCELL_X1 FILLER_63_1172 ();
 FILLCELL_X1 FILLER_63_1177 ();
 FILLCELL_X2 FILLER_63_1182 ();
 FILLCELL_X1 FILLER_63_1184 ();
 FILLCELL_X4 FILLER_63_1191 ();
 FILLCELL_X4 FILLER_63_1199 ();
 FILLCELL_X1 FILLER_63_1203 ();
 FILLCELL_X1 FILLER_63_1223 ();
 FILLCELL_X2 FILLER_63_1264 ();
 FILLCELL_X1 FILLER_63_1289 ();
 FILLCELL_X2 FILLER_63_1292 ();
 FILLCELL_X2 FILLER_63_1314 ();
 FILLCELL_X1 FILLER_63_1357 ();
 FILLCELL_X8 FILLER_63_1388 ();
 FILLCELL_X4 FILLER_63_1396 ();
 FILLCELL_X2 FILLER_63_1411 ();
 FILLCELL_X1 FILLER_63_1413 ();
 FILLCELL_X1 FILLER_63_1438 ();
 FILLCELL_X2 FILLER_63_1442 ();
 FILLCELL_X2 FILLER_63_1472 ();
 FILLCELL_X1 FILLER_63_1474 ();
 FILLCELL_X2 FILLER_63_1484 ();
 FILLCELL_X1 FILLER_63_1486 ();
 FILLCELL_X8 FILLER_63_1498 ();
 FILLCELL_X4 FILLER_63_1506 ();
 FILLCELL_X2 FILLER_63_1510 ();
 FILLCELL_X1 FILLER_63_1512 ();
 FILLCELL_X1 FILLER_63_1516 ();
 FILLCELL_X1 FILLER_63_1521 ();
 FILLCELL_X1 FILLER_63_1533 ();
 FILLCELL_X2 FILLER_63_1559 ();
 FILLCELL_X1 FILLER_63_1565 ();
 FILLCELL_X8 FILLER_63_1570 ();
 FILLCELL_X1 FILLER_63_1578 ();
 FILLCELL_X1 FILLER_63_1588 ();
 FILLCELL_X1 FILLER_63_1595 ();
 FILLCELL_X2 FILLER_63_1604 ();
 FILLCELL_X2 FILLER_63_1613 ();
 FILLCELL_X16 FILLER_63_1621 ();
 FILLCELL_X8 FILLER_63_1637 ();
 FILLCELL_X4 FILLER_63_1645 ();
 FILLCELL_X2 FILLER_63_1649 ();
 FILLCELL_X8 FILLER_64_1 ();
 FILLCELL_X1 FILLER_64_9 ();
 FILLCELL_X32 FILLER_64_14 ();
 FILLCELL_X32 FILLER_64_46 ();
 FILLCELL_X32 FILLER_64_78 ();
 FILLCELL_X32 FILLER_64_110 ();
 FILLCELL_X4 FILLER_64_142 ();
 FILLCELL_X4 FILLER_64_153 ();
 FILLCELL_X2 FILLER_64_157 ();
 FILLCELL_X4 FILLER_64_179 ();
 FILLCELL_X2 FILLER_64_183 ();
 FILLCELL_X4 FILLER_64_209 ();
 FILLCELL_X2 FILLER_64_213 ();
 FILLCELL_X1 FILLER_64_215 ();
 FILLCELL_X8 FILLER_64_243 ();
 FILLCELL_X2 FILLER_64_251 ();
 FILLCELL_X2 FILLER_64_283 ();
 FILLCELL_X1 FILLER_64_292 ();
 FILLCELL_X1 FILLER_64_304 ();
 FILLCELL_X4 FILLER_64_330 ();
 FILLCELL_X2 FILLER_64_334 ();
 FILLCELL_X8 FILLER_64_343 ();
 FILLCELL_X4 FILLER_64_351 ();
 FILLCELL_X2 FILLER_64_355 ();
 FILLCELL_X2 FILLER_64_387 ();
 FILLCELL_X1 FILLER_64_403 ();
 FILLCELL_X8 FILLER_64_415 ();
 FILLCELL_X2 FILLER_64_423 ();
 FILLCELL_X4 FILLER_64_458 ();
 FILLCELL_X2 FILLER_64_462 ();
 FILLCELL_X1 FILLER_64_464 ();
 FILLCELL_X4 FILLER_64_486 ();
 FILLCELL_X2 FILLER_64_490 ();
 FILLCELL_X1 FILLER_64_492 ();
 FILLCELL_X16 FILLER_64_508 ();
 FILLCELL_X8 FILLER_64_524 ();
 FILLCELL_X2 FILLER_64_532 ();
 FILLCELL_X1 FILLER_64_534 ();
 FILLCELL_X2 FILLER_64_545 ();
 FILLCELL_X1 FILLER_64_562 ();
 FILLCELL_X4 FILLER_64_583 ();
 FILLCELL_X2 FILLER_64_587 ();
 FILLCELL_X1 FILLER_64_624 ();
 FILLCELL_X2 FILLER_64_682 ();
 FILLCELL_X1 FILLER_64_684 ();
 FILLCELL_X1 FILLER_64_691 ();
 FILLCELL_X1 FILLER_64_707 ();
 FILLCELL_X2 FILLER_64_714 ();
 FILLCELL_X4 FILLER_64_756 ();
 FILLCELL_X2 FILLER_64_763 ();
 FILLCELL_X1 FILLER_64_765 ();
 FILLCELL_X2 FILLER_64_787 ();
 FILLCELL_X2 FILLER_64_814 ();
 FILLCELL_X1 FILLER_64_841 ();
 FILLCELL_X4 FILLER_64_849 ();
 FILLCELL_X8 FILLER_64_881 ();
 FILLCELL_X2 FILLER_64_889 ();
 FILLCELL_X1 FILLER_64_911 ();
 FILLCELL_X4 FILLER_64_919 ();
 FILLCELL_X2 FILLER_64_923 ();
 FILLCELL_X1 FILLER_64_925 ();
 FILLCELL_X8 FILLER_64_928 ();
 FILLCELL_X1 FILLER_64_936 ();
 FILLCELL_X4 FILLER_64_939 ();
 FILLCELL_X2 FILLER_64_943 ();
 FILLCELL_X16 FILLER_64_976 ();
 FILLCELL_X8 FILLER_64_992 ();
 FILLCELL_X2 FILLER_64_1000 ();
 FILLCELL_X1 FILLER_64_1002 ();
 FILLCELL_X2 FILLER_64_1022 ();
 FILLCELL_X1 FILLER_64_1024 ();
 FILLCELL_X1 FILLER_64_1031 ();
 FILLCELL_X1 FILLER_64_1034 ();
 FILLCELL_X4 FILLER_64_1038 ();
 FILLCELL_X4 FILLER_64_1049 ();
 FILLCELL_X2 FILLER_64_1053 ();
 FILLCELL_X4 FILLER_64_1092 ();
 FILLCELL_X1 FILLER_64_1096 ();
 FILLCELL_X1 FILLER_64_1123 ();
 FILLCELL_X4 FILLER_64_1165 ();
 FILLCELL_X2 FILLER_64_1169 ();
 FILLCELL_X1 FILLER_64_1171 ();
 FILLCELL_X1 FILLER_64_1176 ();
 FILLCELL_X2 FILLER_64_1201 ();
 FILLCELL_X8 FILLER_64_1263 ();
 FILLCELL_X4 FILLER_64_1271 ();
 FILLCELL_X1 FILLER_64_1275 ();
 FILLCELL_X4 FILLER_64_1281 ();
 FILLCELL_X4 FILLER_64_1308 ();
 FILLCELL_X2 FILLER_64_1312 ();
 FILLCELL_X2 FILLER_64_1344 ();
 FILLCELL_X2 FILLER_64_1353 ();
 FILLCELL_X1 FILLER_64_1355 ();
 FILLCELL_X16 FILLER_64_1363 ();
 FILLCELL_X8 FILLER_64_1379 ();
 FILLCELL_X4 FILLER_64_1387 ();
 FILLCELL_X4 FILLER_64_1395 ();
 FILLCELL_X1 FILLER_64_1399 ();
 FILLCELL_X1 FILLER_64_1407 ();
 FILLCELL_X8 FILLER_64_1417 ();
 FILLCELL_X2 FILLER_64_1434 ();
 FILLCELL_X4 FILLER_64_1448 ();
 FILLCELL_X1 FILLER_64_1452 ();
 FILLCELL_X4 FILLER_64_1465 ();
 FILLCELL_X4 FILLER_64_1473 ();
 FILLCELL_X8 FILLER_64_1492 ();
 FILLCELL_X1 FILLER_64_1500 ();
 FILLCELL_X2 FILLER_64_1504 ();
 FILLCELL_X1 FILLER_64_1510 ();
 FILLCELL_X8 FILLER_64_1525 ();
 FILLCELL_X4 FILLER_64_1533 ();
 FILLCELL_X2 FILLER_64_1537 ();
 FILLCELL_X1 FILLER_64_1539 ();
 FILLCELL_X16 FILLER_64_1543 ();
 FILLCELL_X1 FILLER_64_1559 ();
 FILLCELL_X2 FILLER_64_1573 ();
 FILLCELL_X1 FILLER_64_1575 ();
 FILLCELL_X1 FILLER_64_1579 ();
 FILLCELL_X4 FILLER_64_1584 ();
 FILLCELL_X1 FILLER_64_1588 ();
 FILLCELL_X4 FILLER_64_1593 ();
 FILLCELL_X1 FILLER_64_1597 ();
 FILLCELL_X2 FILLER_64_1609 ();
 FILLCELL_X16 FILLER_64_1624 ();
 FILLCELL_X8 FILLER_64_1640 ();
 FILLCELL_X2 FILLER_64_1648 ();
 FILLCELL_X1 FILLER_64_1650 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X2 FILLER_65_129 ();
 FILLCELL_X8 FILLER_65_163 ();
 FILLCELL_X2 FILLER_65_171 ();
 FILLCELL_X1 FILLER_65_173 ();
 FILLCELL_X4 FILLER_65_181 ();
 FILLCELL_X8 FILLER_65_192 ();
 FILLCELL_X4 FILLER_65_200 ();
 FILLCELL_X2 FILLER_65_204 ();
 FILLCELL_X1 FILLER_65_209 ();
 FILLCELL_X16 FILLER_65_217 ();
 FILLCELL_X2 FILLER_65_233 ();
 FILLCELL_X1 FILLER_65_235 ();
 FILLCELL_X4 FILLER_65_244 ();
 FILLCELL_X4 FILLER_65_255 ();
 FILLCELL_X2 FILLER_65_259 ();
 FILLCELL_X1 FILLER_65_265 ();
 FILLCELL_X1 FILLER_65_270 ();
 FILLCELL_X2 FILLER_65_275 ();
 FILLCELL_X2 FILLER_65_288 ();
 FILLCELL_X1 FILLER_65_290 ();
 FILLCELL_X1 FILLER_65_298 ();
 FILLCELL_X2 FILLER_65_310 ();
 FILLCELL_X16 FILLER_65_323 ();
 FILLCELL_X4 FILLER_65_349 ();
 FILLCELL_X1 FILLER_65_353 ();
 FILLCELL_X1 FILLER_65_358 ();
 FILLCELL_X16 FILLER_65_385 ();
 FILLCELL_X8 FILLER_65_401 ();
 FILLCELL_X4 FILLER_65_409 ();
 FILLCELL_X1 FILLER_65_413 ();
 FILLCELL_X4 FILLER_65_421 ();
 FILLCELL_X2 FILLER_65_425 ();
 FILLCELL_X1 FILLER_65_427 ();
 FILLCELL_X4 FILLER_65_437 ();
 FILLCELL_X1 FILLER_65_441 ();
 FILLCELL_X2 FILLER_65_451 ();
 FILLCELL_X4 FILLER_65_460 ();
 FILLCELL_X1 FILLER_65_464 ();
 FILLCELL_X8 FILLER_65_489 ();
 FILLCELL_X4 FILLER_65_497 ();
 FILLCELL_X2 FILLER_65_513 ();
 FILLCELL_X2 FILLER_65_522 ();
 FILLCELL_X1 FILLER_65_540 ();
 FILLCELL_X8 FILLER_65_547 ();
 FILLCELL_X4 FILLER_65_566 ();
 FILLCELL_X8 FILLER_65_592 ();
 FILLCELL_X1 FILLER_65_600 ();
 FILLCELL_X8 FILLER_65_604 ();
 FILLCELL_X1 FILLER_65_612 ();
 FILLCELL_X2 FILLER_65_630 ();
 FILLCELL_X1 FILLER_65_636 ();
 FILLCELL_X4 FILLER_65_641 ();
 FILLCELL_X1 FILLER_65_645 ();
 FILLCELL_X4 FILLER_65_651 ();
 FILLCELL_X16 FILLER_65_659 ();
 FILLCELL_X2 FILLER_65_684 ();
 FILLCELL_X8 FILLER_65_690 ();
 FILLCELL_X2 FILLER_65_698 ();
 FILLCELL_X1 FILLER_65_716 ();
 FILLCELL_X2 FILLER_65_720 ();
 FILLCELL_X2 FILLER_65_726 ();
 FILLCELL_X2 FILLER_65_732 ();
 FILLCELL_X1 FILLER_65_734 ();
 FILLCELL_X16 FILLER_65_746 ();
 FILLCELL_X8 FILLER_65_762 ();
 FILLCELL_X1 FILLER_65_770 ();
 FILLCELL_X1 FILLER_65_786 ();
 FILLCELL_X1 FILLER_65_791 ();
 FILLCELL_X1 FILLER_65_801 ();
 FILLCELL_X1 FILLER_65_823 ();
 FILLCELL_X4 FILLER_65_849 ();
 FILLCELL_X1 FILLER_65_853 ();
 FILLCELL_X2 FILLER_65_858 ();
 FILLCELL_X1 FILLER_65_860 ();
 FILLCELL_X2 FILLER_65_865 ();
 FILLCELL_X2 FILLER_65_871 ();
 FILLCELL_X8 FILLER_65_880 ();
 FILLCELL_X1 FILLER_65_908 ();
 FILLCELL_X2 FILLER_65_921 ();
 FILLCELL_X1 FILLER_65_923 ();
 FILLCELL_X8 FILLER_65_939 ();
 FILLCELL_X4 FILLER_65_947 ();
 FILLCELL_X1 FILLER_65_958 ();
 FILLCELL_X4 FILLER_65_967 ();
 FILLCELL_X1 FILLER_65_971 ();
 FILLCELL_X8 FILLER_65_983 ();
 FILLCELL_X1 FILLER_65_991 ();
 FILLCELL_X2 FILLER_65_995 ();
 FILLCELL_X1 FILLER_65_997 ();
 FILLCELL_X2 FILLER_65_1005 ();
 FILLCELL_X1 FILLER_65_1007 ();
 FILLCELL_X4 FILLER_65_1011 ();
 FILLCELL_X2 FILLER_65_1015 ();
 FILLCELL_X1 FILLER_65_1025 ();
 FILLCELL_X4 FILLER_65_1056 ();
 FILLCELL_X2 FILLER_65_1060 ();
 FILLCELL_X4 FILLER_65_1065 ();
 FILLCELL_X2 FILLER_65_1069 ();
 FILLCELL_X1 FILLER_65_1071 ();
 FILLCELL_X2 FILLER_65_1078 ();
 FILLCELL_X1 FILLER_65_1095 ();
 FILLCELL_X4 FILLER_65_1109 ();
 FILLCELL_X1 FILLER_65_1113 ();
 FILLCELL_X4 FILLER_65_1120 ();
 FILLCELL_X2 FILLER_65_1124 ();
 FILLCELL_X2 FILLER_65_1132 ();
 FILLCELL_X1 FILLER_65_1134 ();
 FILLCELL_X1 FILLER_65_1141 ();
 FILLCELL_X2 FILLER_65_1145 ();
 FILLCELL_X4 FILLER_65_1159 ();
 FILLCELL_X2 FILLER_65_1163 ();
 FILLCELL_X1 FILLER_65_1165 ();
 FILLCELL_X4 FILLER_65_1178 ();
 FILLCELL_X1 FILLER_65_1202 ();
 FILLCELL_X8 FILLER_65_1230 ();
 FILLCELL_X4 FILLER_65_1238 ();
 FILLCELL_X1 FILLER_65_1242 ();
 FILLCELL_X2 FILLER_65_1264 ();
 FILLCELL_X4 FILLER_65_1273 ();
 FILLCELL_X2 FILLER_65_1284 ();
 FILLCELL_X1 FILLER_65_1286 ();
 FILLCELL_X1 FILLER_65_1292 ();
 FILLCELL_X1 FILLER_65_1306 ();
 FILLCELL_X2 FILLER_65_1327 ();
 FILLCELL_X2 FILLER_65_1336 ();
 FILLCELL_X2 FILLER_65_1358 ();
 FILLCELL_X1 FILLER_65_1360 ();
 FILLCELL_X2 FILLER_65_1392 ();
 FILLCELL_X16 FILLER_65_1401 ();
 FILLCELL_X8 FILLER_65_1417 ();
 FILLCELL_X4 FILLER_65_1425 ();
 FILLCELL_X1 FILLER_65_1429 ();
 FILLCELL_X4 FILLER_65_1444 ();
 FILLCELL_X4 FILLER_65_1451 ();
 FILLCELL_X2 FILLER_65_1474 ();
 FILLCELL_X1 FILLER_65_1476 ();
 FILLCELL_X4 FILLER_65_1497 ();
 FILLCELL_X1 FILLER_65_1501 ();
 FILLCELL_X4 FILLER_65_1510 ();
 FILLCELL_X1 FILLER_65_1514 ();
 FILLCELL_X1 FILLER_65_1525 ();
 FILLCELL_X2 FILLER_65_1533 ();
 FILLCELL_X16 FILLER_65_1545 ();
 FILLCELL_X4 FILLER_65_1561 ();
 FILLCELL_X1 FILLER_65_1565 ();
 FILLCELL_X1 FILLER_65_1599 ();
 FILLCELL_X1 FILLER_65_1611 ();
 FILLCELL_X4 FILLER_65_1616 ();
 FILLCELL_X2 FILLER_65_1620 ();
 FILLCELL_X2 FILLER_65_1625 ();
 FILLCELL_X1 FILLER_65_1627 ();
 FILLCELL_X16 FILLER_65_1631 ();
 FILLCELL_X4 FILLER_65_1647 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X2 FILLER_66_129 ();
 FILLCELL_X1 FILLER_66_131 ();
 FILLCELL_X8 FILLER_66_139 ();
 FILLCELL_X8 FILLER_66_174 ();
 FILLCELL_X4 FILLER_66_182 ();
 FILLCELL_X2 FILLER_66_186 ();
 FILLCELL_X1 FILLER_66_210 ();
 FILLCELL_X4 FILLER_66_225 ();
 FILLCELL_X4 FILLER_66_236 ();
 FILLCELL_X1 FILLER_66_240 ();
 FILLCELL_X4 FILLER_66_263 ();
 FILLCELL_X2 FILLER_66_267 ();
 FILLCELL_X1 FILLER_66_269 ();
 FILLCELL_X1 FILLER_66_273 ();
 FILLCELL_X4 FILLER_66_277 ();
 FILLCELL_X2 FILLER_66_281 ();
 FILLCELL_X8 FILLER_66_298 ();
 FILLCELL_X4 FILLER_66_315 ();
 FILLCELL_X2 FILLER_66_323 ();
 FILLCELL_X2 FILLER_66_353 ();
 FILLCELL_X8 FILLER_66_363 ();
 FILLCELL_X2 FILLER_66_371 ();
 FILLCELL_X8 FILLER_66_378 ();
 FILLCELL_X2 FILLER_66_386 ();
 FILLCELL_X1 FILLER_66_403 ();
 FILLCELL_X4 FILLER_66_408 ();
 FILLCELL_X1 FILLER_66_412 ();
 FILLCELL_X4 FILLER_66_447 ();
 FILLCELL_X1 FILLER_66_451 ();
 FILLCELL_X4 FILLER_66_470 ();
 FILLCELL_X2 FILLER_66_474 ();
 FILLCELL_X8 FILLER_66_485 ();
 FILLCELL_X4 FILLER_66_552 ();
 FILLCELL_X1 FILLER_66_556 ();
 FILLCELL_X32 FILLER_66_559 ();
 FILLCELL_X8 FILLER_66_591 ();
 FILLCELL_X8 FILLER_66_616 ();
 FILLCELL_X1 FILLER_66_624 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X2 FILLER_66_632 ();
 FILLCELL_X8 FILLER_66_637 ();
 FILLCELL_X2 FILLER_66_645 ();
 FILLCELL_X8 FILLER_66_667 ();
 FILLCELL_X1 FILLER_66_675 ();
 FILLCELL_X2 FILLER_66_686 ();
 FILLCELL_X4 FILLER_66_708 ();
 FILLCELL_X2 FILLER_66_712 ();
 FILLCELL_X1 FILLER_66_714 ();
 FILLCELL_X4 FILLER_66_720 ();
 FILLCELL_X2 FILLER_66_724 ();
 FILLCELL_X1 FILLER_66_726 ();
 FILLCELL_X2 FILLER_66_731 ();
 FILLCELL_X2 FILLER_66_736 ();
 FILLCELL_X1 FILLER_66_738 ();
 FILLCELL_X2 FILLER_66_746 ();
 FILLCELL_X1 FILLER_66_748 ();
 FILLCELL_X2 FILLER_66_756 ();
 FILLCELL_X2 FILLER_66_778 ();
 FILLCELL_X1 FILLER_66_784 ();
 FILLCELL_X2 FILLER_66_788 ();
 FILLCELL_X2 FILLER_66_801 ();
 FILLCELL_X1 FILLER_66_803 ();
 FILLCELL_X8 FILLER_66_813 ();
 FILLCELL_X4 FILLER_66_848 ();
 FILLCELL_X2 FILLER_66_877 ();
 FILLCELL_X1 FILLER_66_879 ();
 FILLCELL_X2 FILLER_66_900 ();
 FILLCELL_X1 FILLER_66_902 ();
 FILLCELL_X4 FILLER_66_917 ();
 FILLCELL_X2 FILLER_66_921 ();
 FILLCELL_X4 FILLER_66_947 ();
 FILLCELL_X1 FILLER_66_951 ();
 FILLCELL_X1 FILLER_66_964 ();
 FILLCELL_X2 FILLER_66_968 ();
 FILLCELL_X8 FILLER_66_975 ();
 FILLCELL_X1 FILLER_66_986 ();
 FILLCELL_X2 FILLER_66_1012 ();
 FILLCELL_X8 FILLER_66_1021 ();
 FILLCELL_X1 FILLER_66_1029 ();
 FILLCELL_X1 FILLER_66_1032 ();
 FILLCELL_X1 FILLER_66_1045 ();
 FILLCELL_X4 FILLER_66_1049 ();
 FILLCELL_X4 FILLER_66_1066 ();
 FILLCELL_X2 FILLER_66_1070 ();
 FILLCELL_X1 FILLER_66_1072 ();
 FILLCELL_X1 FILLER_66_1076 ();
 FILLCELL_X1 FILLER_66_1099 ();
 FILLCELL_X2 FILLER_66_1134 ();
 FILLCELL_X2 FILLER_66_1142 ();
 FILLCELL_X1 FILLER_66_1172 ();
 FILLCELL_X2 FILLER_66_1179 ();
 FILLCELL_X1 FILLER_66_1181 ();
 FILLCELL_X32 FILLER_66_1197 ();
 FILLCELL_X2 FILLER_66_1229 ();
 FILLCELL_X8 FILLER_66_1245 ();
 FILLCELL_X1 FILLER_66_1253 ();
 FILLCELL_X1 FILLER_66_1329 ();
 FILLCELL_X16 FILLER_66_1337 ();
 FILLCELL_X2 FILLER_66_1353 ();
 FILLCELL_X1 FILLER_66_1355 ();
 FILLCELL_X2 FILLER_66_1363 ();
 FILLCELL_X2 FILLER_66_1369 ();
 FILLCELL_X2 FILLER_66_1391 ();
 FILLCELL_X1 FILLER_66_1393 ();
 FILLCELL_X2 FILLER_66_1401 ();
 FILLCELL_X1 FILLER_66_1403 ();
 FILLCELL_X2 FILLER_66_1411 ();
 FILLCELL_X2 FILLER_66_1417 ();
 FILLCELL_X1 FILLER_66_1419 ();
 FILLCELL_X4 FILLER_66_1444 ();
 FILLCELL_X1 FILLER_66_1448 ();
 FILLCELL_X4 FILLER_66_1458 ();
 FILLCELL_X1 FILLER_66_1462 ();
 FILLCELL_X2 FILLER_66_1470 ();
 FILLCELL_X2 FILLER_66_1481 ();
 FILLCELL_X16 FILLER_66_1503 ();
 FILLCELL_X1 FILLER_66_1519 ();
 FILLCELL_X1 FILLER_66_1543 ();
 FILLCELL_X4 FILLER_66_1556 ();
 FILLCELL_X1 FILLER_66_1560 ();
 FILLCELL_X1 FILLER_66_1568 ();
 FILLCELL_X1 FILLER_66_1572 ();
 FILLCELL_X2 FILLER_66_1601 ();
 FILLCELL_X2 FILLER_66_1613 ();
 FILLCELL_X1 FILLER_66_1615 ();
 FILLCELL_X4 FILLER_66_1624 ();
 FILLCELL_X2 FILLER_66_1628 ();
 FILLCELL_X8 FILLER_66_1633 ();
 FILLCELL_X4 FILLER_66_1641 ();
 FILLCELL_X2 FILLER_66_1648 ();
 FILLCELL_X1 FILLER_66_1650 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X1 FILLER_67_129 ();
 FILLCELL_X8 FILLER_67_137 ();
 FILLCELL_X4 FILLER_67_145 ();
 FILLCELL_X1 FILLER_67_149 ();
 FILLCELL_X8 FILLER_67_170 ();
 FILLCELL_X8 FILLER_67_185 ();
 FILLCELL_X2 FILLER_67_200 ();
 FILLCELL_X1 FILLER_67_202 ();
 FILLCELL_X4 FILLER_67_206 ();
 FILLCELL_X1 FILLER_67_210 ();
 FILLCELL_X4 FILLER_67_220 ();
 FILLCELL_X2 FILLER_67_231 ();
 FILLCELL_X4 FILLER_67_236 ();
 FILLCELL_X1 FILLER_67_244 ();
 FILLCELL_X8 FILLER_67_261 ();
 FILLCELL_X2 FILLER_67_294 ();
 FILLCELL_X2 FILLER_67_299 ();
 FILLCELL_X1 FILLER_67_301 ();
 FILLCELL_X2 FILLER_67_313 ();
 FILLCELL_X1 FILLER_67_315 ();
 FILLCELL_X16 FILLER_67_318 ();
 FILLCELL_X1 FILLER_67_334 ();
 FILLCELL_X1 FILLER_67_367 ();
 FILLCELL_X2 FILLER_67_374 ();
 FILLCELL_X1 FILLER_67_376 ();
 FILLCELL_X8 FILLER_67_384 ();
 FILLCELL_X4 FILLER_67_392 ();
 FILLCELL_X1 FILLER_67_410 ();
 FILLCELL_X8 FILLER_67_420 ();
 FILLCELL_X4 FILLER_67_431 ();
 FILLCELL_X4 FILLER_67_438 ();
 FILLCELL_X2 FILLER_67_442 ();
 FILLCELL_X2 FILLER_67_454 ();
 FILLCELL_X16 FILLER_67_459 ();
 FILLCELL_X4 FILLER_67_475 ();
 FILLCELL_X1 FILLER_67_479 ();
 FILLCELL_X8 FILLER_67_516 ();
 FILLCELL_X2 FILLER_67_524 ();
 FILLCELL_X1 FILLER_67_562 ();
 FILLCELL_X2 FILLER_67_585 ();
 FILLCELL_X1 FILLER_67_587 ();
 FILLCELL_X2 FILLER_67_612 ();
 FILLCELL_X1 FILLER_67_614 ();
 FILLCELL_X4 FILLER_67_622 ();
 FILLCELL_X2 FILLER_67_626 ();
 FILLCELL_X4 FILLER_67_641 ();
 FILLCELL_X2 FILLER_67_645 ();
 FILLCELL_X8 FILLER_67_654 ();
 FILLCELL_X2 FILLER_67_662 ();
 FILLCELL_X1 FILLER_67_684 ();
 FILLCELL_X4 FILLER_67_718 ();
 FILLCELL_X2 FILLER_67_722 ();
 FILLCELL_X1 FILLER_67_724 ();
 FILLCELL_X1 FILLER_67_734 ();
 FILLCELL_X1 FILLER_67_739 ();
 FILLCELL_X2 FILLER_67_760 ();
 FILLCELL_X8 FILLER_67_770 ();
 FILLCELL_X2 FILLER_67_778 ();
 FILLCELL_X4 FILLER_67_787 ();
 FILLCELL_X2 FILLER_67_811 ();
 FILLCELL_X16 FILLER_67_827 ();
 FILLCELL_X8 FILLER_67_865 ();
 FILLCELL_X4 FILLER_67_873 ();
 FILLCELL_X2 FILLER_67_877 ();
 FILLCELL_X4 FILLER_67_899 ();
 FILLCELL_X4 FILLER_67_910 ();
 FILLCELL_X1 FILLER_67_914 ();
 FILLCELL_X4 FILLER_67_917 ();
 FILLCELL_X2 FILLER_67_921 ();
 FILLCELL_X1 FILLER_67_923 ();
 FILLCELL_X2 FILLER_67_934 ();
 FILLCELL_X1 FILLER_67_936 ();
 FILLCELL_X1 FILLER_67_942 ();
 FILLCELL_X4 FILLER_67_945 ();
 FILLCELL_X2 FILLER_67_949 ();
 FILLCELL_X2 FILLER_67_968 ();
 FILLCELL_X4 FILLER_67_1001 ();
 FILLCELL_X2 FILLER_67_1005 ();
 FILLCELL_X8 FILLER_67_1023 ();
 FILLCELL_X2 FILLER_67_1031 ();
 FILLCELL_X2 FILLER_67_1061 ();
 FILLCELL_X8 FILLER_67_1087 ();
 FILLCELL_X2 FILLER_67_1095 ();
 FILLCELL_X8 FILLER_67_1104 ();
 FILLCELL_X2 FILLER_67_1112 ();
 FILLCELL_X8 FILLER_67_1126 ();
 FILLCELL_X2 FILLER_67_1134 ();
 FILLCELL_X1 FILLER_67_1136 ();
 FILLCELL_X4 FILLER_67_1155 ();
 FILLCELL_X1 FILLER_67_1159 ();
 FILLCELL_X2 FILLER_67_1202 ();
 FILLCELL_X2 FILLER_67_1216 ();
 FILLCELL_X4 FILLER_67_1225 ();
 FILLCELL_X2 FILLER_67_1229 ();
 FILLCELL_X2 FILLER_67_1252 ();
 FILLCELL_X2 FILLER_67_1261 ();
 FILLCELL_X8 FILLER_67_1271 ();
 FILLCELL_X4 FILLER_67_1293 ();
 FILLCELL_X1 FILLER_67_1297 ();
 FILLCELL_X2 FILLER_67_1320 ();
 FILLCELL_X2 FILLER_67_1369 ();
 FILLCELL_X1 FILLER_67_1371 ();
 FILLCELL_X1 FILLER_67_1386 ();
 FILLCELL_X1 FILLER_67_1407 ();
 FILLCELL_X1 FILLER_67_1415 ();
 FILLCELL_X32 FILLER_67_1420 ();
 FILLCELL_X2 FILLER_67_1452 ();
 FILLCELL_X1 FILLER_67_1454 ();
 FILLCELL_X1 FILLER_67_1465 ();
 FILLCELL_X1 FILLER_67_1479 ();
 FILLCELL_X4 FILLER_67_1485 ();
 FILLCELL_X1 FILLER_67_1489 ();
 FILLCELL_X8 FILLER_67_1494 ();
 FILLCELL_X2 FILLER_67_1502 ();
 FILLCELL_X1 FILLER_67_1504 ();
 FILLCELL_X1 FILLER_67_1510 ();
 FILLCELL_X1 FILLER_67_1529 ();
 FILLCELL_X1 FILLER_67_1537 ();
 FILLCELL_X4 FILLER_67_1542 ();
 FILLCELL_X16 FILLER_67_1558 ();
 FILLCELL_X8 FILLER_67_1574 ();
 FILLCELL_X4 FILLER_67_1582 ();
 FILLCELL_X32 FILLER_67_1619 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X16 FILLER_68_97 ();
 FILLCELL_X8 FILLER_68_113 ();
 FILLCELL_X4 FILLER_68_121 ();
 FILLCELL_X2 FILLER_68_125 ();
 FILLCELL_X4 FILLER_68_147 ();
 FILLCELL_X1 FILLER_68_151 ();
 FILLCELL_X1 FILLER_68_166 ();
 FILLCELL_X1 FILLER_68_174 ();
 FILLCELL_X2 FILLER_68_195 ();
 FILLCELL_X2 FILLER_68_204 ();
 FILLCELL_X1 FILLER_68_206 ();
 FILLCELL_X1 FILLER_68_249 ();
 FILLCELL_X2 FILLER_68_257 ();
 FILLCELL_X2 FILLER_68_295 ();
 FILLCELL_X4 FILLER_68_322 ();
 FILLCELL_X2 FILLER_68_326 ();
 FILLCELL_X16 FILLER_68_332 ();
 FILLCELL_X1 FILLER_68_348 ();
 FILLCELL_X1 FILLER_68_401 ();
 FILLCELL_X1 FILLER_68_406 ();
 FILLCELL_X1 FILLER_68_411 ();
 FILLCELL_X8 FILLER_68_416 ();
 FILLCELL_X1 FILLER_68_456 ();
 FILLCELL_X1 FILLER_68_461 ();
 FILLCELL_X16 FILLER_68_472 ();
 FILLCELL_X2 FILLER_68_488 ();
 FILLCELL_X1 FILLER_68_490 ();
 FILLCELL_X2 FILLER_68_508 ();
 FILLCELL_X1 FILLER_68_510 ();
 FILLCELL_X8 FILLER_68_515 ();
 FILLCELL_X4 FILLER_68_523 ();
 FILLCELL_X1 FILLER_68_534 ();
 FILLCELL_X1 FILLER_68_543 ();
 FILLCELL_X1 FILLER_68_554 ();
 FILLCELL_X1 FILLER_68_559 ();
 FILLCELL_X2 FILLER_68_571 ();
 FILLCELL_X1 FILLER_68_573 ();
 FILLCELL_X1 FILLER_68_584 ();
 FILLCELL_X4 FILLER_68_596 ();
 FILLCELL_X1 FILLER_68_600 ();
 FILLCELL_X2 FILLER_68_604 ();
 FILLCELL_X1 FILLER_68_606 ();
 FILLCELL_X8 FILLER_68_620 ();
 FILLCELL_X2 FILLER_68_628 ();
 FILLCELL_X1 FILLER_68_630 ();
 FILLCELL_X1 FILLER_68_676 ();
 FILLCELL_X1 FILLER_68_684 ();
 FILLCELL_X4 FILLER_68_692 ();
 FILLCELL_X2 FILLER_68_720 ();
 FILLCELL_X1 FILLER_68_722 ();
 FILLCELL_X1 FILLER_68_734 ();
 FILLCELL_X1 FILLER_68_738 ();
 FILLCELL_X1 FILLER_68_748 ();
 FILLCELL_X8 FILLER_68_755 ();
 FILLCELL_X1 FILLER_68_763 ();
 FILLCELL_X2 FILLER_68_771 ();
 FILLCELL_X1 FILLER_68_773 ();
 FILLCELL_X16 FILLER_68_794 ();
 FILLCELL_X8 FILLER_68_810 ();
 FILLCELL_X2 FILLER_68_818 ();
 FILLCELL_X8 FILLER_68_823 ();
 FILLCELL_X4 FILLER_68_831 ();
 FILLCELL_X2 FILLER_68_835 ();
 FILLCELL_X8 FILLER_68_844 ();
 FILLCELL_X1 FILLER_68_852 ();
 FILLCELL_X2 FILLER_68_873 ();
 FILLCELL_X2 FILLER_68_895 ();
 FILLCELL_X1 FILLER_68_897 ();
 FILLCELL_X1 FILLER_68_903 ();
 FILLCELL_X4 FILLER_68_919 ();
 FILLCELL_X2 FILLER_68_923 ();
 FILLCELL_X1 FILLER_68_925 ();
 FILLCELL_X1 FILLER_68_931 ();
 FILLCELL_X1 FILLER_68_960 ();
 FILLCELL_X4 FILLER_68_988 ();
 FILLCELL_X2 FILLER_68_992 ();
 FILLCELL_X1 FILLER_68_994 ();
 FILLCELL_X8 FILLER_68_1013 ();
 FILLCELL_X2 FILLER_68_1021 ();
 FILLCELL_X4 FILLER_68_1038 ();
 FILLCELL_X1 FILLER_68_1042 ();
 FILLCELL_X4 FILLER_68_1049 ();
 FILLCELL_X2 FILLER_68_1053 ();
 FILLCELL_X8 FILLER_68_1058 ();
 FILLCELL_X2 FILLER_68_1066 ();
 FILLCELL_X1 FILLER_68_1068 ();
 FILLCELL_X1 FILLER_68_1077 ();
 FILLCELL_X2 FILLER_68_1085 ();
 FILLCELL_X1 FILLER_68_1087 ();
 FILLCELL_X1 FILLER_68_1091 ();
 FILLCELL_X4 FILLER_68_1112 ();
 FILLCELL_X2 FILLER_68_1126 ();
 FILLCELL_X1 FILLER_68_1128 ();
 FILLCELL_X2 FILLER_68_1133 ();
 FILLCELL_X1 FILLER_68_1135 ();
 FILLCELL_X1 FILLER_68_1145 ();
 FILLCELL_X1 FILLER_68_1152 ();
 FILLCELL_X4 FILLER_68_1166 ();
 FILLCELL_X2 FILLER_68_1170 ();
 FILLCELL_X8 FILLER_68_1190 ();
 FILLCELL_X2 FILLER_68_1198 ();
 FILLCELL_X2 FILLER_68_1214 ();
 FILLCELL_X1 FILLER_68_1216 ();
 FILLCELL_X4 FILLER_68_1237 ();
 FILLCELL_X2 FILLER_68_1241 ();
 FILLCELL_X1 FILLER_68_1250 ();
 FILLCELL_X8 FILLER_68_1267 ();
 FILLCELL_X4 FILLER_68_1275 ();
 FILLCELL_X1 FILLER_68_1279 ();
 FILLCELL_X4 FILLER_68_1287 ();
 FILLCELL_X2 FILLER_68_1303 ();
 FILLCELL_X1 FILLER_68_1305 ();
 FILLCELL_X2 FILLER_68_1326 ();
 FILLCELL_X1 FILLER_68_1328 ();
 FILLCELL_X4 FILLER_68_1336 ();
 FILLCELL_X2 FILLER_68_1340 ();
 FILLCELL_X4 FILLER_68_1362 ();
 FILLCELL_X1 FILLER_68_1366 ();
 FILLCELL_X8 FILLER_68_1387 ();
 FILLCELL_X4 FILLER_68_1395 ();
 FILLCELL_X2 FILLER_68_1399 ();
 FILLCELL_X1 FILLER_68_1401 ();
 FILLCELL_X4 FILLER_68_1406 ();
 FILLCELL_X2 FILLER_68_1410 ();
 FILLCELL_X1 FILLER_68_1412 ();
 FILLCELL_X32 FILLER_68_1417 ();
 FILLCELL_X4 FILLER_68_1449 ();
 FILLCELL_X2 FILLER_68_1453 ();
 FILLCELL_X4 FILLER_68_1462 ();
 FILLCELL_X2 FILLER_68_1466 ();
 FILLCELL_X1 FILLER_68_1468 ();
 FILLCELL_X4 FILLER_68_1473 ();
 FILLCELL_X1 FILLER_68_1477 ();
 FILLCELL_X2 FILLER_68_1482 ();
 FILLCELL_X1 FILLER_68_1484 ();
 FILLCELL_X1 FILLER_68_1491 ();
 FILLCELL_X2 FILLER_68_1496 ();
 FILLCELL_X1 FILLER_68_1498 ();
 FILLCELL_X4 FILLER_68_1508 ();
 FILLCELL_X2 FILLER_68_1512 ();
 FILLCELL_X2 FILLER_68_1518 ();
 FILLCELL_X1 FILLER_68_1520 ();
 FILLCELL_X4 FILLER_68_1530 ();
 FILLCELL_X2 FILLER_68_1534 ();
 FILLCELL_X1 FILLER_68_1536 ();
 FILLCELL_X1 FILLER_68_1544 ();
 FILLCELL_X1 FILLER_68_1552 ();
 FILLCELL_X1 FILLER_68_1558 ();
 FILLCELL_X2 FILLER_68_1562 ();
 FILLCELL_X1 FILLER_68_1578 ();
 FILLCELL_X1 FILLER_68_1584 ();
 FILLCELL_X4 FILLER_68_1630 ();
 FILLCELL_X8 FILLER_68_1637 ();
 FILLCELL_X4 FILLER_68_1645 ();
 FILLCELL_X2 FILLER_68_1649 ();
 FILLCELL_X2 FILLER_69_1 ();
 FILLCELL_X1 FILLER_69_3 ();
 FILLCELL_X32 FILLER_69_7 ();
 FILLCELL_X32 FILLER_69_39 ();
 FILLCELL_X32 FILLER_69_71 ();
 FILLCELL_X16 FILLER_69_103 ();
 FILLCELL_X4 FILLER_69_119 ();
 FILLCELL_X2 FILLER_69_123 ();
 FILLCELL_X8 FILLER_69_152 ();
 FILLCELL_X4 FILLER_69_160 ();
 FILLCELL_X1 FILLER_69_164 ();
 FILLCELL_X2 FILLER_69_223 ();
 FILLCELL_X1 FILLER_69_225 ();
 FILLCELL_X2 FILLER_69_243 ();
 FILLCELL_X1 FILLER_69_245 ();
 FILLCELL_X32 FILLER_69_260 ();
 FILLCELL_X2 FILLER_69_292 ();
 FILLCELL_X2 FILLER_69_301 ();
 FILLCELL_X1 FILLER_69_303 ();
 FILLCELL_X2 FILLER_69_328 ();
 FILLCELL_X1 FILLER_69_330 ();
 FILLCELL_X1 FILLER_69_355 ();
 FILLCELL_X1 FILLER_69_362 ();
 FILLCELL_X1 FILLER_69_372 ();
 FILLCELL_X4 FILLER_69_379 ();
 FILLCELL_X2 FILLER_69_383 ();
 FILLCELL_X4 FILLER_69_411 ();
 FILLCELL_X1 FILLER_69_418 ();
 FILLCELL_X8 FILLER_69_423 ();
 FILLCELL_X2 FILLER_69_431 ();
 FILLCELL_X1 FILLER_69_433 ();
 FILLCELL_X1 FILLER_69_443 ();
 FILLCELL_X2 FILLER_69_497 ();
 FILLCELL_X1 FILLER_69_499 ();
 FILLCELL_X8 FILLER_69_512 ();
 FILLCELL_X2 FILLER_69_520 ();
 FILLCELL_X1 FILLER_69_522 ();
 FILLCELL_X2 FILLER_69_527 ();
 FILLCELL_X1 FILLER_69_529 ();
 FILLCELL_X2 FILLER_69_550 ();
 FILLCELL_X2 FILLER_69_573 ();
 FILLCELL_X1 FILLER_69_575 ();
 FILLCELL_X8 FILLER_69_579 ();
 FILLCELL_X1 FILLER_69_587 ();
 FILLCELL_X4 FILLER_69_603 ();
 FILLCELL_X2 FILLER_69_607 ();
 FILLCELL_X16 FILLER_69_612 ();
 FILLCELL_X1 FILLER_69_631 ();
 FILLCELL_X2 FILLER_69_639 ();
 FILLCELL_X2 FILLER_69_648 ();
 FILLCELL_X4 FILLER_69_664 ();
 FILLCELL_X1 FILLER_69_668 ();
 FILLCELL_X1 FILLER_69_685 ();
 FILLCELL_X8 FILLER_69_699 ();
 FILLCELL_X4 FILLER_69_707 ();
 FILLCELL_X2 FILLER_69_711 ();
 FILLCELL_X8 FILLER_69_717 ();
 FILLCELL_X4 FILLER_69_725 ();
 FILLCELL_X1 FILLER_69_729 ();
 FILLCELL_X4 FILLER_69_734 ();
 FILLCELL_X2 FILLER_69_738 ();
 FILLCELL_X1 FILLER_69_740 ();
 FILLCELL_X4 FILLER_69_752 ();
 FILLCELL_X1 FILLER_69_759 ();
 FILLCELL_X1 FILLER_69_783 ();
 FILLCELL_X4 FILLER_69_791 ();
 FILLCELL_X2 FILLER_69_795 ();
 FILLCELL_X1 FILLER_69_797 ();
 FILLCELL_X2 FILLER_69_818 ();
 FILLCELL_X1 FILLER_69_820 ();
 FILLCELL_X1 FILLER_69_828 ();
 FILLCELL_X8 FILLER_69_856 ();
 FILLCELL_X8 FILLER_69_889 ();
 FILLCELL_X4 FILLER_69_897 ();
 FILLCELL_X2 FILLER_69_901 ();
 FILLCELL_X1 FILLER_69_903 ();
 FILLCELL_X1 FILLER_69_909 ();
 FILLCELL_X4 FILLER_69_941 ();
 FILLCELL_X1 FILLER_69_945 ();
 FILLCELL_X1 FILLER_69_948 ();
 FILLCELL_X4 FILLER_69_965 ();
 FILLCELL_X1 FILLER_69_969 ();
 FILLCELL_X4 FILLER_69_976 ();
 FILLCELL_X1 FILLER_69_980 ();
 FILLCELL_X1 FILLER_69_988 ();
 FILLCELL_X1 FILLER_69_995 ();
 FILLCELL_X4 FILLER_69_1001 ();
 FILLCELL_X1 FILLER_69_1007 ();
 FILLCELL_X1 FILLER_69_1035 ();
 FILLCELL_X2 FILLER_69_1063 ();
 FILLCELL_X1 FILLER_69_1068 ();
 FILLCELL_X4 FILLER_69_1081 ();
 FILLCELL_X4 FILLER_69_1091 ();
 FILLCELL_X1 FILLER_69_1095 ();
 FILLCELL_X8 FILLER_69_1105 ();
 FILLCELL_X1 FILLER_69_1113 ();
 FILLCELL_X1 FILLER_69_1149 ();
 FILLCELL_X8 FILLER_69_1156 ();
 FILLCELL_X2 FILLER_69_1164 ();
 FILLCELL_X2 FILLER_69_1169 ();
 FILLCELL_X2 FILLER_69_1177 ();
 FILLCELL_X1 FILLER_69_1179 ();
 FILLCELL_X2 FILLER_69_1190 ();
 FILLCELL_X1 FILLER_69_1192 ();
 FILLCELL_X2 FILLER_69_1200 ();
 FILLCELL_X1 FILLER_69_1202 ();
 FILLCELL_X2 FILLER_69_1210 ();
 FILLCELL_X1 FILLER_69_1212 ();
 FILLCELL_X2 FILLER_69_1218 ();
 FILLCELL_X1 FILLER_69_1262 ();
 FILLCELL_X1 FILLER_69_1264 ();
 FILLCELL_X2 FILLER_69_1279 ();
 FILLCELL_X1 FILLER_69_1286 ();
 FILLCELL_X1 FILLER_69_1296 ();
 FILLCELL_X2 FILLER_69_1304 ();
 FILLCELL_X2 FILLER_69_1326 ();
 FILLCELL_X2 FILLER_69_1335 ();
 FILLCELL_X2 FILLER_69_1344 ();
 FILLCELL_X1 FILLER_69_1346 ();
 FILLCELL_X8 FILLER_69_1354 ();
 FILLCELL_X4 FILLER_69_1362 ();
 FILLCELL_X2 FILLER_69_1366 ();
 FILLCELL_X1 FILLER_69_1368 ();
 FILLCELL_X32 FILLER_69_1396 ();
 FILLCELL_X32 FILLER_69_1428 ();
 FILLCELL_X8 FILLER_69_1460 ();
 FILLCELL_X4 FILLER_69_1468 ();
 FILLCELL_X8 FILLER_69_1488 ();
 FILLCELL_X2 FILLER_69_1496 ();
 FILLCELL_X1 FILLER_69_1514 ();
 FILLCELL_X4 FILLER_69_1526 ();
 FILLCELL_X1 FILLER_69_1530 ();
 FILLCELL_X8 FILLER_69_1534 ();
 FILLCELL_X2 FILLER_69_1542 ();
 FILLCELL_X1 FILLER_69_1544 ();
 FILLCELL_X1 FILLER_69_1552 ();
 FILLCELL_X2 FILLER_69_1576 ();
 FILLCELL_X2 FILLER_69_1602 ();
 FILLCELL_X4 FILLER_69_1622 ();
 FILLCELL_X2 FILLER_69_1626 ();
 FILLCELL_X16 FILLER_69_1631 ();
 FILLCELL_X4 FILLER_69_1647 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X16 FILLER_70_97 ();
 FILLCELL_X8 FILLER_70_113 ();
 FILLCELL_X4 FILLER_70_121 ();
 FILLCELL_X2 FILLER_70_125 ();
 FILLCELL_X4 FILLER_70_154 ();
 FILLCELL_X4 FILLER_70_166 ();
 FILLCELL_X8 FILLER_70_197 ();
 FILLCELL_X1 FILLER_70_205 ();
 FILLCELL_X2 FILLER_70_210 ();
 FILLCELL_X2 FILLER_70_223 ();
 FILLCELL_X8 FILLER_70_244 ();
 FILLCELL_X4 FILLER_70_252 ();
 FILLCELL_X2 FILLER_70_256 ();
 FILLCELL_X8 FILLER_70_265 ();
 FILLCELL_X4 FILLER_70_273 ();
 FILLCELL_X4 FILLER_70_291 ();
 FILLCELL_X1 FILLER_70_299 ();
 FILLCELL_X4 FILLER_70_320 ();
 FILLCELL_X2 FILLER_70_324 ();
 FILLCELL_X1 FILLER_70_333 ();
 FILLCELL_X1 FILLER_70_338 ();
 FILLCELL_X2 FILLER_70_357 ();
 FILLCELL_X1 FILLER_70_359 ();
 FILLCELL_X4 FILLER_70_377 ();
 FILLCELL_X2 FILLER_70_381 ();
 FILLCELL_X1 FILLER_70_383 ();
 FILLCELL_X16 FILLER_70_387 ();
 FILLCELL_X8 FILLER_70_403 ();
 FILLCELL_X4 FILLER_70_411 ();
 FILLCELL_X8 FILLER_70_442 ();
 FILLCELL_X4 FILLER_70_450 ();
 FILLCELL_X2 FILLER_70_478 ();
 FILLCELL_X1 FILLER_70_493 ();
 FILLCELL_X4 FILLER_70_528 ();
 FILLCELL_X8 FILLER_70_537 ();
 FILLCELL_X4 FILLER_70_545 ();
 FILLCELL_X8 FILLER_70_566 ();
 FILLCELL_X2 FILLER_70_574 ();
 FILLCELL_X1 FILLER_70_576 ();
 FILLCELL_X2 FILLER_70_586 ();
 FILLCELL_X1 FILLER_70_626 ();
 FILLCELL_X1 FILLER_70_652 ();
 FILLCELL_X1 FILLER_70_664 ();
 FILLCELL_X2 FILLER_70_668 ();
 FILLCELL_X4 FILLER_70_681 ();
 FILLCELL_X1 FILLER_70_685 ();
 FILLCELL_X2 FILLER_70_706 ();
 FILLCELL_X1 FILLER_70_708 ();
 FILLCELL_X1 FILLER_70_713 ();
 FILLCELL_X1 FILLER_70_734 ();
 FILLCELL_X1 FILLER_70_740 ();
 FILLCELL_X1 FILLER_70_771 ();
 FILLCELL_X2 FILLER_70_776 ();
 FILLCELL_X1 FILLER_70_788 ();
 FILLCELL_X2 FILLER_70_809 ();
 FILLCELL_X2 FILLER_70_818 ();
 FILLCELL_X2 FILLER_70_824 ();
 FILLCELL_X1 FILLER_70_826 ();
 FILLCELL_X16 FILLER_70_848 ();
 FILLCELL_X4 FILLER_70_864 ();
 FILLCELL_X2 FILLER_70_868 ();
 FILLCELL_X1 FILLER_70_910 ();
 FILLCELL_X4 FILLER_70_923 ();
 FILLCELL_X1 FILLER_70_947 ();
 FILLCELL_X8 FILLER_70_955 ();
 FILLCELL_X4 FILLER_70_963 ();
 FILLCELL_X2 FILLER_70_967 ();
 FILLCELL_X1 FILLER_70_969 ();
 FILLCELL_X8 FILLER_70_1017 ();
 FILLCELL_X2 FILLER_70_1025 ();
 FILLCELL_X16 FILLER_70_1050 ();
 FILLCELL_X2 FILLER_70_1072 ();
 FILLCELL_X1 FILLER_70_1096 ();
 FILLCELL_X4 FILLER_70_1107 ();
 FILLCELL_X2 FILLER_70_1111 ();
 FILLCELL_X2 FILLER_70_1149 ();
 FILLCELL_X1 FILLER_70_1161 ();
 FILLCELL_X1 FILLER_70_1175 ();
 FILLCELL_X8 FILLER_70_1188 ();
 FILLCELL_X1 FILLER_70_1196 ();
 FILLCELL_X8 FILLER_70_1204 ();
 FILLCELL_X4 FILLER_70_1212 ();
 FILLCELL_X2 FILLER_70_1216 ();
 FILLCELL_X4 FILLER_70_1225 ();
 FILLCELL_X1 FILLER_70_1229 ();
 FILLCELL_X4 FILLER_70_1237 ();
 FILLCELL_X1 FILLER_70_1241 ();
 FILLCELL_X2 FILLER_70_1262 ();
 FILLCELL_X1 FILLER_70_1268 ();
 FILLCELL_X1 FILLER_70_1274 ();
 FILLCELL_X4 FILLER_70_1297 ();
 FILLCELL_X8 FILLER_70_1310 ();
 FILLCELL_X2 FILLER_70_1318 ();
 FILLCELL_X1 FILLER_70_1320 ();
 FILLCELL_X4 FILLER_70_1328 ();
 FILLCELL_X2 FILLER_70_1332 ();
 FILLCELL_X1 FILLER_70_1334 ();
 FILLCELL_X4 FILLER_70_1355 ();
 FILLCELL_X1 FILLER_70_1359 ();
 FILLCELL_X4 FILLER_70_1388 ();
 FILLCELL_X2 FILLER_70_1392 ();
 FILLCELL_X1 FILLER_70_1394 ();
 FILLCELL_X32 FILLER_70_1415 ();
 FILLCELL_X16 FILLER_70_1447 ();
 FILLCELL_X8 FILLER_70_1463 ();
 FILLCELL_X2 FILLER_70_1471 ();
 FILLCELL_X4 FILLER_70_1491 ();
 FILLCELL_X1 FILLER_70_1495 ();
 FILLCELL_X2 FILLER_70_1514 ();
 FILLCELL_X1 FILLER_70_1516 ();
 FILLCELL_X4 FILLER_70_1530 ();
 FILLCELL_X1 FILLER_70_1534 ();
 FILLCELL_X2 FILLER_70_1544 ();
 FILLCELL_X4 FILLER_70_1553 ();
 FILLCELL_X2 FILLER_70_1557 ();
 FILLCELL_X4 FILLER_70_1575 ();
 FILLCELL_X1 FILLER_70_1579 ();
 FILLCELL_X1 FILLER_70_1591 ();
 FILLCELL_X1 FILLER_70_1598 ();
 FILLCELL_X2 FILLER_70_1612 ();
 FILLCELL_X16 FILLER_70_1623 ();
 FILLCELL_X8 FILLER_70_1639 ();
 FILLCELL_X4 FILLER_70_1647 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X4 FILLER_71_129 ();
 FILLCELL_X2 FILLER_71_133 ();
 FILLCELL_X1 FILLER_71_135 ();
 FILLCELL_X2 FILLER_71_143 ();
 FILLCELL_X1 FILLER_71_145 ();
 FILLCELL_X32 FILLER_71_173 ();
 FILLCELL_X4 FILLER_71_205 ();
 FILLCELL_X1 FILLER_71_209 ();
 FILLCELL_X8 FILLER_71_213 ();
 FILLCELL_X1 FILLER_71_221 ();
 FILLCELL_X2 FILLER_71_229 ();
 FILLCELL_X2 FILLER_71_242 ();
 FILLCELL_X1 FILLER_71_244 ();
 FILLCELL_X8 FILLER_71_250 ();
 FILLCELL_X4 FILLER_71_272 ();
 FILLCELL_X1 FILLER_71_276 ();
 FILLCELL_X1 FILLER_71_284 ();
 FILLCELL_X2 FILLER_71_299 ();
 FILLCELL_X2 FILLER_71_316 ();
 FILLCELL_X4 FILLER_71_342 ();
 FILLCELL_X1 FILLER_71_346 ();
 FILLCELL_X1 FILLER_71_357 ();
 FILLCELL_X1 FILLER_71_367 ();
 FILLCELL_X8 FILLER_71_397 ();
 FILLCELL_X4 FILLER_71_405 ();
 FILLCELL_X2 FILLER_71_409 ();
 FILLCELL_X1 FILLER_71_411 ();
 FILLCELL_X4 FILLER_71_419 ();
 FILLCELL_X2 FILLER_71_423 ();
 FILLCELL_X1 FILLER_71_425 ();
 FILLCELL_X16 FILLER_71_440 ();
 FILLCELL_X2 FILLER_71_456 ();
 FILLCELL_X1 FILLER_71_458 ();
 FILLCELL_X8 FILLER_71_464 ();
 FILLCELL_X4 FILLER_71_472 ();
 FILLCELL_X2 FILLER_71_486 ();
 FILLCELL_X2 FILLER_71_492 ();
 FILLCELL_X8 FILLER_71_501 ();
 FILLCELL_X1 FILLER_71_509 ();
 FILLCELL_X8 FILLER_71_528 ();
 FILLCELL_X4 FILLER_71_536 ();
 FILLCELL_X2 FILLER_71_560 ();
 FILLCELL_X2 FILLER_71_572 ();
 FILLCELL_X8 FILLER_71_578 ();
 FILLCELL_X1 FILLER_71_586 ();
 FILLCELL_X4 FILLER_71_597 ();
 FILLCELL_X1 FILLER_71_601 ();
 FILLCELL_X4 FILLER_71_622 ();
 FILLCELL_X1 FILLER_71_626 ();
 FILLCELL_X2 FILLER_71_649 ();
 FILLCELL_X1 FILLER_71_651 ();
 FILLCELL_X2 FILLER_71_677 ();
 FILLCELL_X1 FILLER_71_679 ();
 FILLCELL_X4 FILLER_71_684 ();
 FILLCELL_X1 FILLER_71_705 ();
 FILLCELL_X1 FILLER_71_708 ();
 FILLCELL_X4 FILLER_71_719 ();
 FILLCELL_X2 FILLER_71_723 ();
 FILLCELL_X1 FILLER_71_725 ();
 FILLCELL_X1 FILLER_71_743 ();
 FILLCELL_X1 FILLER_71_755 ();
 FILLCELL_X1 FILLER_71_774 ();
 FILLCELL_X2 FILLER_71_802 ();
 FILLCELL_X2 FILLER_71_808 ();
 FILLCELL_X2 FILLER_71_813 ();
 FILLCELL_X1 FILLER_71_815 ();
 FILLCELL_X1 FILLER_71_842 ();
 FILLCELL_X4 FILLER_71_867 ();
 FILLCELL_X2 FILLER_71_871 ();
 FILLCELL_X1 FILLER_71_873 ();
 FILLCELL_X1 FILLER_71_879 ();
 FILLCELL_X1 FILLER_71_887 ();
 FILLCELL_X2 FILLER_71_959 ();
 FILLCELL_X1 FILLER_71_961 ();
 FILLCELL_X8 FILLER_71_966 ();
 FILLCELL_X1 FILLER_71_974 ();
 FILLCELL_X1 FILLER_71_997 ();
 FILLCELL_X2 FILLER_71_1001 ();
 FILLCELL_X16 FILLER_71_1013 ();
 FILLCELL_X4 FILLER_71_1029 ();
 FILLCELL_X2 FILLER_71_1033 ();
 FILLCELL_X1 FILLER_71_1042 ();
 FILLCELL_X2 FILLER_71_1066 ();
 FILLCELL_X8 FILLER_71_1077 ();
 FILLCELL_X1 FILLER_71_1085 ();
 FILLCELL_X4 FILLER_71_1090 ();
 FILLCELL_X4 FILLER_71_1098 ();
 FILLCELL_X1 FILLER_71_1108 ();
 FILLCELL_X1 FILLER_71_1121 ();
 FILLCELL_X2 FILLER_71_1128 ();
 FILLCELL_X1 FILLER_71_1130 ();
 FILLCELL_X8 FILLER_71_1137 ();
 FILLCELL_X4 FILLER_71_1145 ();
 FILLCELL_X2 FILLER_71_1149 ();
 FILLCELL_X4 FILLER_71_1171 ();
 FILLCELL_X16 FILLER_71_1188 ();
 FILLCELL_X1 FILLER_71_1204 ();
 FILLCELL_X8 FILLER_71_1212 ();
 FILLCELL_X1 FILLER_71_1220 ();
 FILLCELL_X1 FILLER_71_1334 ();
 FILLCELL_X4 FILLER_71_1340 ();
 FILLCELL_X2 FILLER_71_1344 ();
 FILLCELL_X1 FILLER_71_1346 ();
 FILLCELL_X4 FILLER_71_1354 ();
 FILLCELL_X4 FILLER_71_1385 ();
 FILLCELL_X2 FILLER_71_1389 ();
 FILLCELL_X1 FILLER_71_1391 ();
 FILLCELL_X2 FILLER_71_1396 ();
 FILLCELL_X16 FILLER_71_1405 ();
 FILLCELL_X1 FILLER_71_1421 ();
 FILLCELL_X1 FILLER_71_1426 ();
 FILLCELL_X16 FILLER_71_1443 ();
 FILLCELL_X4 FILLER_71_1459 ();
 FILLCELL_X32 FILLER_71_1476 ();
 FILLCELL_X8 FILLER_71_1508 ();
 FILLCELL_X2 FILLER_71_1516 ();
 FILLCELL_X4 FILLER_71_1527 ();
 FILLCELL_X1 FILLER_71_1552 ();
 FILLCELL_X32 FILLER_71_1567 ();
 FILLCELL_X32 FILLER_71_1599 ();
 FILLCELL_X16 FILLER_71_1631 ();
 FILLCELL_X4 FILLER_71_1647 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X16 FILLER_72_97 ();
 FILLCELL_X8 FILLER_72_113 ();
 FILLCELL_X2 FILLER_72_121 ();
 FILLCELL_X4 FILLER_72_143 ();
 FILLCELL_X2 FILLER_72_147 ();
 FILLCELL_X4 FILLER_72_191 ();
 FILLCELL_X1 FILLER_72_195 ();
 FILLCELL_X2 FILLER_72_216 ();
 FILLCELL_X16 FILLER_72_238 ();
 FILLCELL_X4 FILLER_72_254 ();
 FILLCELL_X4 FILLER_72_310 ();
 FILLCELL_X2 FILLER_72_314 ();
 FILLCELL_X1 FILLER_72_316 ();
 FILLCELL_X4 FILLER_72_326 ();
 FILLCELL_X1 FILLER_72_337 ();
 FILLCELL_X4 FILLER_72_348 ();
 FILLCELL_X1 FILLER_72_370 ();
 FILLCELL_X8 FILLER_72_379 ();
 FILLCELL_X2 FILLER_72_387 ();
 FILLCELL_X1 FILLER_72_413 ();
 FILLCELL_X1 FILLER_72_421 ();
 FILLCELL_X1 FILLER_72_436 ();
 FILLCELL_X1 FILLER_72_444 ();
 FILLCELL_X2 FILLER_72_452 ();
 FILLCELL_X2 FILLER_72_495 ();
 FILLCELL_X8 FILLER_72_501 ();
 FILLCELL_X4 FILLER_72_509 ();
 FILLCELL_X16 FILLER_72_526 ();
 FILLCELL_X8 FILLER_72_549 ();
 FILLCELL_X2 FILLER_72_557 ();
 FILLCELL_X2 FILLER_72_586 ();
 FILLCELL_X8 FILLER_72_602 ();
 FILLCELL_X1 FILLER_72_610 ();
 FILLCELL_X4 FILLER_72_614 ();
 FILLCELL_X2 FILLER_72_618 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X8 FILLER_72_632 ();
 FILLCELL_X4 FILLER_72_640 ();
 FILLCELL_X1 FILLER_72_666 ();
 FILLCELL_X1 FILLER_72_682 ();
 FILLCELL_X1 FILLER_72_690 ();
 FILLCELL_X4 FILLER_72_709 ();
 FILLCELL_X2 FILLER_72_717 ();
 FILLCELL_X2 FILLER_72_739 ();
 FILLCELL_X1 FILLER_72_741 ();
 FILLCELL_X8 FILLER_72_752 ();
 FILLCELL_X2 FILLER_72_763 ();
 FILLCELL_X2 FILLER_72_771 ();
 FILLCELL_X1 FILLER_72_773 ();
 FILLCELL_X1 FILLER_72_800 ();
 FILLCELL_X8 FILLER_72_822 ();
 FILLCELL_X1 FILLER_72_834 ();
 FILLCELL_X16 FILLER_72_848 ();
 FILLCELL_X8 FILLER_72_864 ();
 FILLCELL_X2 FILLER_72_872 ();
 FILLCELL_X1 FILLER_72_917 ();
 FILLCELL_X8 FILLER_72_926 ();
 FILLCELL_X4 FILLER_72_934 ();
 FILLCELL_X2 FILLER_72_945 ();
 FILLCELL_X4 FILLER_72_973 ();
 FILLCELL_X2 FILLER_72_977 ();
 FILLCELL_X1 FILLER_72_979 ();
 FILLCELL_X16 FILLER_72_987 ();
 FILLCELL_X4 FILLER_72_1003 ();
 FILLCELL_X2 FILLER_72_1018 ();
 FILLCELL_X4 FILLER_72_1053 ();
 FILLCELL_X2 FILLER_72_1091 ();
 FILLCELL_X2 FILLER_72_1096 ();
 FILLCELL_X1 FILLER_72_1098 ();
 FILLCELL_X2 FILLER_72_1120 ();
 FILLCELL_X1 FILLER_72_1122 ();
 FILLCELL_X1 FILLER_72_1129 ();
 FILLCELL_X4 FILLER_72_1154 ();
 FILLCELL_X2 FILLER_72_1158 ();
 FILLCELL_X1 FILLER_72_1188 ();
 FILLCELL_X1 FILLER_72_1199 ();
 FILLCELL_X1 FILLER_72_1207 ();
 FILLCELL_X8 FILLER_72_1228 ();
 FILLCELL_X2 FILLER_72_1236 ();
 FILLCELL_X1 FILLER_72_1245 ();
 FILLCELL_X4 FILLER_72_1253 ();
 FILLCELL_X1 FILLER_72_1265 ();
 FILLCELL_X1 FILLER_72_1276 ();
 FILLCELL_X1 FILLER_72_1304 ();
 FILLCELL_X1 FILLER_72_1349 ();
 FILLCELL_X1 FILLER_72_1357 ();
 FILLCELL_X1 FILLER_72_1378 ();
 FILLCELL_X1 FILLER_72_1399 ();
 FILLCELL_X8 FILLER_72_1407 ();
 FILLCELL_X4 FILLER_72_1415 ();
 FILLCELL_X1 FILLER_72_1419 ();
 FILLCELL_X2 FILLER_72_1443 ();
 FILLCELL_X8 FILLER_72_1472 ();
 FILLCELL_X2 FILLER_72_1480 ();
 FILLCELL_X8 FILLER_72_1491 ();
 FILLCELL_X4 FILLER_72_1499 ();
 FILLCELL_X32 FILLER_72_1510 ();
 FILLCELL_X8 FILLER_72_1542 ();
 FILLCELL_X8 FILLER_72_1555 ();
 FILLCELL_X4 FILLER_72_1563 ();
 FILLCELL_X2 FILLER_72_1567 ();
 FILLCELL_X32 FILLER_72_1587 ();
 FILLCELL_X4 FILLER_72_1619 ();
 FILLCELL_X1 FILLER_72_1623 ();
 FILLCELL_X16 FILLER_72_1627 ();
 FILLCELL_X8 FILLER_72_1643 ();
 FILLCELL_X8 FILLER_73_1 ();
 FILLCELL_X4 FILLER_73_9 ();
 FILLCELL_X2 FILLER_73_13 ();
 FILLCELL_X1 FILLER_73_15 ();
 FILLCELL_X32 FILLER_73_19 ();
 FILLCELL_X32 FILLER_73_51 ();
 FILLCELL_X32 FILLER_73_83 ();
 FILLCELL_X8 FILLER_73_115 ();
 FILLCELL_X2 FILLER_73_123 ();
 FILLCELL_X8 FILLER_73_132 ();
 FILLCELL_X4 FILLER_73_140 ();
 FILLCELL_X2 FILLER_73_144 ();
 FILLCELL_X16 FILLER_73_153 ();
 FILLCELL_X4 FILLER_73_169 ();
 FILLCELL_X4 FILLER_73_180 ();
 FILLCELL_X1 FILLER_73_184 ();
 FILLCELL_X2 FILLER_73_207 ();
 FILLCELL_X1 FILLER_73_216 ();
 FILLCELL_X1 FILLER_73_223 ();
 FILLCELL_X1 FILLER_73_229 ();
 FILLCELL_X1 FILLER_73_236 ();
 FILLCELL_X4 FILLER_73_243 ();
 FILLCELL_X2 FILLER_73_247 ();
 FILLCELL_X8 FILLER_73_276 ();
 FILLCELL_X4 FILLER_73_284 ();
 FILLCELL_X2 FILLER_73_288 ();
 FILLCELL_X1 FILLER_73_297 ();
 FILLCELL_X2 FILLER_73_302 ();
 FILLCELL_X1 FILLER_73_304 ();
 FILLCELL_X2 FILLER_73_320 ();
 FILLCELL_X1 FILLER_73_322 ();
 FILLCELL_X4 FILLER_73_346 ();
 FILLCELL_X1 FILLER_73_365 ();
 FILLCELL_X8 FILLER_73_369 ();
 FILLCELL_X2 FILLER_73_377 ();
 FILLCELL_X1 FILLER_73_379 ();
 FILLCELL_X2 FILLER_73_460 ();
 FILLCELL_X1 FILLER_73_484 ();
 FILLCELL_X4 FILLER_73_495 ();
 FILLCELL_X2 FILLER_73_499 ();
 FILLCELL_X4 FILLER_73_527 ();
 FILLCELL_X2 FILLER_73_531 ();
 FILLCELL_X2 FILLER_73_562 ();
 FILLCELL_X4 FILLER_73_570 ();
 FILLCELL_X2 FILLER_73_574 ();
 FILLCELL_X4 FILLER_73_579 ();
 FILLCELL_X1 FILLER_73_583 ();
 FILLCELL_X4 FILLER_73_608 ();
 FILLCELL_X1 FILLER_73_612 ();
 FILLCELL_X1 FILLER_73_617 ();
 FILLCELL_X1 FILLER_73_620 ();
 FILLCELL_X8 FILLER_73_630 ();
 FILLCELL_X4 FILLER_73_638 ();
 FILLCELL_X2 FILLER_73_660 ();
 FILLCELL_X8 FILLER_73_718 ();
 FILLCELL_X1 FILLER_73_726 ();
 FILLCELL_X16 FILLER_73_755 ();
 FILLCELL_X1 FILLER_73_771 ();
 FILLCELL_X2 FILLER_73_784 ();
 FILLCELL_X32 FILLER_73_847 ();
 FILLCELL_X16 FILLER_73_879 ();
 FILLCELL_X4 FILLER_73_895 ();
 FILLCELL_X2 FILLER_73_899 ();
 FILLCELL_X2 FILLER_73_923 ();
 FILLCELL_X1 FILLER_73_936 ();
 FILLCELL_X2 FILLER_73_944 ();
 FILLCELL_X1 FILLER_73_962 ();
 FILLCELL_X4 FILLER_73_967 ();
 FILLCELL_X2 FILLER_73_971 ();
 FILLCELL_X2 FILLER_73_998 ();
 FILLCELL_X4 FILLER_73_1027 ();
 FILLCELL_X2 FILLER_73_1056 ();
 FILLCELL_X1 FILLER_73_1058 ();
 FILLCELL_X2 FILLER_73_1075 ();
 FILLCELL_X1 FILLER_73_1083 ();
 FILLCELL_X2 FILLER_73_1090 ();
 FILLCELL_X2 FILLER_73_1099 ();
 FILLCELL_X2 FILLER_73_1114 ();
 FILLCELL_X1 FILLER_73_1116 ();
 FILLCELL_X8 FILLER_73_1123 ();
 FILLCELL_X1 FILLER_73_1131 ();
 FILLCELL_X2 FILLER_73_1141 ();
 FILLCELL_X16 FILLER_73_1149 ();
 FILLCELL_X8 FILLER_73_1165 ();
 FILLCELL_X1 FILLER_73_1173 ();
 FILLCELL_X8 FILLER_73_1181 ();
 FILLCELL_X2 FILLER_73_1189 ();
 FILLCELL_X8 FILLER_73_1205 ();
 FILLCELL_X4 FILLER_73_1213 ();
 FILLCELL_X1 FILLER_73_1217 ();
 FILLCELL_X4 FILLER_73_1225 ();
 FILLCELL_X1 FILLER_73_1229 ();
 FILLCELL_X8 FILLER_73_1252 ();
 FILLCELL_X2 FILLER_73_1260 ();
 FILLCELL_X1 FILLER_73_1262 ();
 FILLCELL_X2 FILLER_73_1264 ();
 FILLCELL_X1 FILLER_73_1276 ();
 FILLCELL_X4 FILLER_73_1287 ();
 FILLCELL_X2 FILLER_73_1311 ();
 FILLCELL_X1 FILLER_73_1313 ();
 FILLCELL_X16 FILLER_73_1334 ();
 FILLCELL_X2 FILLER_73_1350 ();
 FILLCELL_X1 FILLER_73_1352 ();
 FILLCELL_X8 FILLER_73_1380 ();
 FILLCELL_X1 FILLER_73_1388 ();
 FILLCELL_X16 FILLER_73_1413 ();
 FILLCELL_X8 FILLER_73_1429 ();
 FILLCELL_X1 FILLER_73_1462 ();
 FILLCELL_X4 FILLER_73_1470 ();
 FILLCELL_X1 FILLER_73_1483 ();
 FILLCELL_X2 FILLER_73_1493 ();
 FILLCELL_X2 FILLER_73_1498 ();
 FILLCELL_X1 FILLER_73_1512 ();
 FILLCELL_X1 FILLER_73_1540 ();
 FILLCELL_X32 FILLER_73_1545 ();
 FILLCELL_X32 FILLER_73_1577 ();
 FILLCELL_X32 FILLER_73_1609 ();
 FILLCELL_X8 FILLER_73_1641 ();
 FILLCELL_X2 FILLER_73_1649 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X1 FILLER_74_129 ();
 FILLCELL_X2 FILLER_74_157 ();
 FILLCELL_X4 FILLER_74_181 ();
 FILLCELL_X1 FILLER_74_185 ();
 FILLCELL_X4 FILLER_74_191 ();
 FILLCELL_X2 FILLER_74_195 ();
 FILLCELL_X1 FILLER_74_197 ();
 FILLCELL_X1 FILLER_74_213 ();
 FILLCELL_X2 FILLER_74_220 ();
 FILLCELL_X2 FILLER_74_248 ();
 FILLCELL_X8 FILLER_74_257 ();
 FILLCELL_X4 FILLER_74_265 ();
 FILLCELL_X2 FILLER_74_269 ();
 FILLCELL_X1 FILLER_74_271 ();
 FILLCELL_X4 FILLER_74_293 ();
 FILLCELL_X2 FILLER_74_297 ();
 FILLCELL_X1 FILLER_74_299 ();
 FILLCELL_X16 FILLER_74_337 ();
 FILLCELL_X1 FILLER_74_353 ();
 FILLCELL_X4 FILLER_74_375 ();
 FILLCELL_X2 FILLER_74_379 ();
 FILLCELL_X4 FILLER_74_388 ();
 FILLCELL_X8 FILLER_74_399 ();
 FILLCELL_X4 FILLER_74_407 ();
 FILLCELL_X2 FILLER_74_411 ();
 FILLCELL_X2 FILLER_74_420 ();
 FILLCELL_X1 FILLER_74_422 ();
 FILLCELL_X1 FILLER_74_452 ();
 FILLCELL_X8 FILLER_74_456 ();
 FILLCELL_X4 FILLER_74_464 ();
 FILLCELL_X8 FILLER_74_475 ();
 FILLCELL_X1 FILLER_74_483 ();
 FILLCELL_X4 FILLER_74_493 ();
 FILLCELL_X2 FILLER_74_497 ();
 FILLCELL_X1 FILLER_74_499 ();
 FILLCELL_X1 FILLER_74_520 ();
 FILLCELL_X16 FILLER_74_524 ();
 FILLCELL_X2 FILLER_74_540 ();
 FILLCELL_X1 FILLER_74_542 ();
 FILLCELL_X2 FILLER_74_561 ();
 FILLCELL_X2 FILLER_74_572 ();
 FILLCELL_X1 FILLER_74_574 ();
 FILLCELL_X4 FILLER_74_602 ();
 FILLCELL_X2 FILLER_74_606 ();
 FILLCELL_X1 FILLER_74_615 ();
 FILLCELL_X2 FILLER_74_628 ();
 FILLCELL_X1 FILLER_74_630 ();
 FILLCELL_X16 FILLER_74_661 ();
 FILLCELL_X8 FILLER_74_677 ();
 FILLCELL_X2 FILLER_74_685 ();
 FILLCELL_X2 FILLER_74_691 ();
 FILLCELL_X1 FILLER_74_704 ();
 FILLCELL_X2 FILLER_74_734 ();
 FILLCELL_X1 FILLER_74_736 ();
 FILLCELL_X8 FILLER_74_746 ();
 FILLCELL_X1 FILLER_74_754 ();
 FILLCELL_X1 FILLER_74_757 ();
 FILLCELL_X8 FILLER_74_767 ();
 FILLCELL_X2 FILLER_74_775 ();
 FILLCELL_X1 FILLER_74_777 ();
 FILLCELL_X2 FILLER_74_785 ();
 FILLCELL_X1 FILLER_74_787 ();
 FILLCELL_X2 FILLER_74_791 ();
 FILLCELL_X1 FILLER_74_797 ();
 FILLCELL_X2 FILLER_74_801 ();
 FILLCELL_X2 FILLER_74_823 ();
 FILLCELL_X1 FILLER_74_825 ();
 FILLCELL_X8 FILLER_74_853 ();
 FILLCELL_X4 FILLER_74_861 ();
 FILLCELL_X1 FILLER_74_890 ();
 FILLCELL_X4 FILLER_74_898 ();
 FILLCELL_X2 FILLER_74_902 ();
 FILLCELL_X8 FILLER_74_906 ();
 FILLCELL_X4 FILLER_74_916 ();
 FILLCELL_X2 FILLER_74_920 ();
 FILLCELL_X1 FILLER_74_922 ();
 FILLCELL_X4 FILLER_74_928 ();
 FILLCELL_X1 FILLER_74_932 ();
 FILLCELL_X16 FILLER_74_964 ();
 FILLCELL_X8 FILLER_74_980 ();
 FILLCELL_X4 FILLER_74_988 ();
 FILLCELL_X2 FILLER_74_992 ();
 FILLCELL_X1 FILLER_74_994 ();
 FILLCELL_X8 FILLER_74_1023 ();
 FILLCELL_X4 FILLER_74_1031 ();
 FILLCELL_X2 FILLER_74_1035 ();
 FILLCELL_X4 FILLER_74_1047 ();
 FILLCELL_X1 FILLER_74_1051 ();
 FILLCELL_X8 FILLER_74_1069 ();
 FILLCELL_X2 FILLER_74_1077 ();
 FILLCELL_X4 FILLER_74_1095 ();
 FILLCELL_X1 FILLER_74_1099 ();
 FILLCELL_X1 FILLER_74_1107 ();
 FILLCELL_X8 FILLER_74_1115 ();
 FILLCELL_X4 FILLER_74_1123 ();
 FILLCELL_X2 FILLER_74_1153 ();
 FILLCELL_X1 FILLER_74_1155 ();
 FILLCELL_X4 FILLER_74_1163 ();
 FILLCELL_X2 FILLER_74_1167 ();
 FILLCELL_X16 FILLER_74_1173 ();
 FILLCELL_X8 FILLER_74_1189 ();
 FILLCELL_X2 FILLER_74_1225 ();
 FILLCELL_X8 FILLER_74_1247 ();
 FILLCELL_X4 FILLER_74_1255 ();
 FILLCELL_X2 FILLER_74_1298 ();
 FILLCELL_X1 FILLER_74_1300 ();
 FILLCELL_X1 FILLER_74_1308 ();
 FILLCELL_X2 FILLER_74_1316 ();
 FILLCELL_X1 FILLER_74_1318 ();
 FILLCELL_X2 FILLER_74_1326 ();
 FILLCELL_X1 FILLER_74_1328 ();
 FILLCELL_X2 FILLER_74_1336 ();
 FILLCELL_X1 FILLER_74_1338 ();
 FILLCELL_X2 FILLER_74_1359 ();
 FILLCELL_X1 FILLER_74_1361 ();
 FILLCELL_X4 FILLER_74_1369 ();
 FILLCELL_X1 FILLER_74_1373 ();
 FILLCELL_X4 FILLER_74_1381 ();
 FILLCELL_X1 FILLER_74_1385 ();
 FILLCELL_X4 FILLER_74_1390 ();
 FILLCELL_X2 FILLER_74_1401 ();
 FILLCELL_X2 FILLER_74_1423 ();
 FILLCELL_X1 FILLER_74_1425 ();
 FILLCELL_X8 FILLER_74_1433 ();
 FILLCELL_X2 FILLER_74_1441 ();
 FILLCELL_X1 FILLER_74_1506 ();
 FILLCELL_X1 FILLER_74_1510 ();
 FILLCELL_X2 FILLER_74_1520 ();
 FILLCELL_X2 FILLER_74_1531 ();
 FILLCELL_X1 FILLER_74_1533 ();
 FILLCELL_X2 FILLER_74_1537 ();
 FILLCELL_X1 FILLER_74_1539 ();
 FILLCELL_X2 FILLER_74_1551 ();
 FILLCELL_X1 FILLER_74_1558 ();
 FILLCELL_X1 FILLER_74_1566 ();
 FILLCELL_X2 FILLER_74_1579 ();
 FILLCELL_X1 FILLER_74_1581 ();
 FILLCELL_X32 FILLER_74_1598 ();
 FILLCELL_X16 FILLER_74_1630 ();
 FILLCELL_X4 FILLER_74_1646 ();
 FILLCELL_X1 FILLER_74_1650 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X2 FILLER_75_129 ();
 FILLCELL_X2 FILLER_75_138 ();
 FILLCELL_X8 FILLER_75_148 ();
 FILLCELL_X1 FILLER_75_156 ();
 FILLCELL_X8 FILLER_75_186 ();
 FILLCELL_X4 FILLER_75_194 ();
 FILLCELL_X2 FILLER_75_198 ();
 FILLCELL_X1 FILLER_75_200 ();
 FILLCELL_X2 FILLER_75_207 ();
 FILLCELL_X4 FILLER_75_221 ();
 FILLCELL_X2 FILLER_75_225 ();
 FILLCELL_X8 FILLER_75_231 ();
 FILLCELL_X4 FILLER_75_239 ();
 FILLCELL_X1 FILLER_75_243 ();
 FILLCELL_X2 FILLER_75_253 ();
 FILLCELL_X1 FILLER_75_255 ();
 FILLCELL_X4 FILLER_75_263 ();
 FILLCELL_X2 FILLER_75_267 ();
 FILLCELL_X1 FILLER_75_269 ();
 FILLCELL_X4 FILLER_75_277 ();
 FILLCELL_X2 FILLER_75_281 ();
 FILLCELL_X1 FILLER_75_283 ();
 FILLCELL_X8 FILLER_75_358 ();
 FILLCELL_X1 FILLER_75_373 ();
 FILLCELL_X1 FILLER_75_381 ();
 FILLCELL_X2 FILLER_75_409 ();
 FILLCELL_X1 FILLER_75_411 ();
 FILLCELL_X2 FILLER_75_419 ();
 FILLCELL_X16 FILLER_75_429 ();
 FILLCELL_X4 FILLER_75_445 ();
 FILLCELL_X1 FILLER_75_459 ();
 FILLCELL_X4 FILLER_75_470 ();
 FILLCELL_X1 FILLER_75_474 ();
 FILLCELL_X8 FILLER_75_493 ();
 FILLCELL_X1 FILLER_75_531 ();
 FILLCELL_X8 FILLER_75_538 ();
 FILLCELL_X4 FILLER_75_546 ();
 FILLCELL_X16 FILLER_75_557 ();
 FILLCELL_X1 FILLER_75_573 ();
 FILLCELL_X4 FILLER_75_599 ();
 FILLCELL_X2 FILLER_75_603 ();
 FILLCELL_X1 FILLER_75_605 ();
 FILLCELL_X1 FILLER_75_612 ();
 FILLCELL_X2 FILLER_75_616 ();
 FILLCELL_X2 FILLER_75_627 ();
 FILLCELL_X2 FILLER_75_635 ();
 FILLCELL_X1 FILLER_75_637 ();
 FILLCELL_X2 FILLER_75_645 ();
 FILLCELL_X1 FILLER_75_647 ();
 FILLCELL_X4 FILLER_75_651 ();
 FILLCELL_X2 FILLER_75_655 ();
 FILLCELL_X8 FILLER_75_678 ();
 FILLCELL_X2 FILLER_75_686 ();
 FILLCELL_X1 FILLER_75_688 ();
 FILLCELL_X2 FILLER_75_698 ();
 FILLCELL_X2 FILLER_75_713 ();
 FILLCELL_X2 FILLER_75_718 ();
 FILLCELL_X1 FILLER_75_720 ();
 FILLCELL_X4 FILLER_75_724 ();
 FILLCELL_X2 FILLER_75_728 ();
 FILLCELL_X8 FILLER_75_739 ();
 FILLCELL_X1 FILLER_75_747 ();
 FILLCELL_X2 FILLER_75_751 ();
 FILLCELL_X8 FILLER_75_814 ();
 FILLCELL_X8 FILLER_75_827 ();
 FILLCELL_X2 FILLER_75_835 ();
 FILLCELL_X8 FILLER_75_883 ();
 FILLCELL_X4 FILLER_75_891 ();
 FILLCELL_X1 FILLER_75_895 ();
 FILLCELL_X8 FILLER_75_913 ();
 FILLCELL_X4 FILLER_75_921 ();
 FILLCELL_X2 FILLER_75_928 ();
 FILLCELL_X4 FILLER_75_936 ();
 FILLCELL_X1 FILLER_75_940 ();
 FILLCELL_X1 FILLER_75_946 ();
 FILLCELL_X2 FILLER_75_950 ();
 FILLCELL_X1 FILLER_75_952 ();
 FILLCELL_X1 FILLER_75_957 ();
 FILLCELL_X2 FILLER_75_971 ();
 FILLCELL_X1 FILLER_75_976 ();
 FILLCELL_X2 FILLER_75_984 ();
 FILLCELL_X2 FILLER_75_1020 ();
 FILLCELL_X4 FILLER_75_1028 ();
 FILLCELL_X4 FILLER_75_1039 ();
 FILLCELL_X1 FILLER_75_1043 ();
 FILLCELL_X1 FILLER_75_1053 ();
 FILLCELL_X8 FILLER_75_1057 ();
 FILLCELL_X1 FILLER_75_1065 ();
 FILLCELL_X4 FILLER_75_1072 ();
 FILLCELL_X1 FILLER_75_1076 ();
 FILLCELL_X4 FILLER_75_1106 ();
 FILLCELL_X2 FILLER_75_1110 ();
 FILLCELL_X2 FILLER_75_1131 ();
 FILLCELL_X2 FILLER_75_1137 ();
 FILLCELL_X2 FILLER_75_1148 ();
 FILLCELL_X8 FILLER_75_1188 ();
 FILLCELL_X2 FILLER_75_1196 ();
 FILLCELL_X1 FILLER_75_1198 ();
 FILLCELL_X4 FILLER_75_1213 ();
 FILLCELL_X2 FILLER_75_1217 ();
 FILLCELL_X8 FILLER_75_1226 ();
 FILLCELL_X2 FILLER_75_1257 ();
 FILLCELL_X2 FILLER_75_1293 ();
 FILLCELL_X4 FILLER_75_1315 ();
 FILLCELL_X2 FILLER_75_1319 ();
 FILLCELL_X1 FILLER_75_1321 ();
 FILLCELL_X4 FILLER_75_1336 ();
 FILLCELL_X4 FILLER_75_1360 ();
 FILLCELL_X1 FILLER_75_1364 ();
 FILLCELL_X2 FILLER_75_1368 ();
 FILLCELL_X1 FILLER_75_1370 ();
 FILLCELL_X4 FILLER_75_1378 ();
 FILLCELL_X2 FILLER_75_1382 ();
 FILLCELL_X1 FILLER_75_1384 ();
 FILLCELL_X16 FILLER_75_1392 ();
 FILLCELL_X8 FILLER_75_1408 ();
 FILLCELL_X2 FILLER_75_1416 ();
 FILLCELL_X1 FILLER_75_1418 ();
 FILLCELL_X4 FILLER_75_1424 ();
 FILLCELL_X1 FILLER_75_1428 ();
 FILLCELL_X4 FILLER_75_1438 ();
 FILLCELL_X2 FILLER_75_1442 ();
 FILLCELL_X1 FILLER_75_1444 ();
 FILLCELL_X8 FILLER_75_1452 ();
 FILLCELL_X4 FILLER_75_1460 ();
 FILLCELL_X2 FILLER_75_1464 ();
 FILLCELL_X1 FILLER_75_1466 ();
 FILLCELL_X1 FILLER_75_1476 ();
 FILLCELL_X2 FILLER_75_1482 ();
 FILLCELL_X16 FILLER_75_1489 ();
 FILLCELL_X1 FILLER_75_1505 ();
 FILLCELL_X2 FILLER_75_1509 ();
 FILLCELL_X1 FILLER_75_1511 ();
 FILLCELL_X1 FILLER_75_1539 ();
 FILLCELL_X1 FILLER_75_1544 ();
 FILLCELL_X1 FILLER_75_1554 ();
 FILLCELL_X4 FILLER_75_1564 ();
 FILLCELL_X8 FILLER_75_1593 ();
 FILLCELL_X8 FILLER_75_1610 ();
 FILLCELL_X2 FILLER_75_1618 ();
 FILLCELL_X4 FILLER_75_1625 ();
 FILLCELL_X2 FILLER_75_1629 ();
 FILLCELL_X16 FILLER_75_1634 ();
 FILLCELL_X1 FILLER_75_1650 ();
 FILLCELL_X16 FILLER_76_1 ();
 FILLCELL_X4 FILLER_76_17 ();
 FILLCELL_X2 FILLER_76_21 ();
 FILLCELL_X32 FILLER_76_27 ();
 FILLCELL_X32 FILLER_76_59 ();
 FILLCELL_X32 FILLER_76_91 ();
 FILLCELL_X2 FILLER_76_143 ();
 FILLCELL_X1 FILLER_76_145 ();
 FILLCELL_X4 FILLER_76_153 ();
 FILLCELL_X2 FILLER_76_157 ();
 FILLCELL_X4 FILLER_76_166 ();
 FILLCELL_X2 FILLER_76_170 ();
 FILLCELL_X4 FILLER_76_179 ();
 FILLCELL_X1 FILLER_76_183 ();
 FILLCELL_X1 FILLER_76_204 ();
 FILLCELL_X2 FILLER_76_215 ();
 FILLCELL_X4 FILLER_76_221 ();
 FILLCELL_X2 FILLER_76_242 ();
 FILLCELL_X1 FILLER_76_244 ();
 FILLCELL_X4 FILLER_76_251 ();
 FILLCELL_X8 FILLER_76_260 ();
 FILLCELL_X4 FILLER_76_268 ();
 FILLCELL_X8 FILLER_76_285 ();
 FILLCELL_X4 FILLER_76_293 ();
 FILLCELL_X1 FILLER_76_297 ();
 FILLCELL_X16 FILLER_76_343 ();
 FILLCELL_X1 FILLER_76_359 ();
 FILLCELL_X1 FILLER_76_383 ();
 FILLCELL_X2 FILLER_76_427 ();
 FILLCELL_X1 FILLER_76_429 ();
 FILLCELL_X8 FILLER_76_437 ();
 FILLCELL_X1 FILLER_76_445 ();
 FILLCELL_X4 FILLER_76_466 ();
 FILLCELL_X2 FILLER_76_470 ();
 FILLCELL_X4 FILLER_76_502 ();
 FILLCELL_X2 FILLER_76_506 ();
 FILLCELL_X2 FILLER_76_515 ();
 FILLCELL_X1 FILLER_76_517 ();
 FILLCELL_X1 FILLER_76_551 ();
 FILLCELL_X16 FILLER_76_569 ();
 FILLCELL_X1 FILLER_76_585 ();
 FILLCELL_X2 FILLER_76_595 ();
 FILLCELL_X8 FILLER_76_620 ();
 FILLCELL_X2 FILLER_76_628 ();
 FILLCELL_X1 FILLER_76_630 ();
 FILLCELL_X2 FILLER_76_632 ();
 FILLCELL_X1 FILLER_76_634 ();
 FILLCELL_X4 FILLER_76_638 ();
 FILLCELL_X8 FILLER_76_646 ();
 FILLCELL_X2 FILLER_76_654 ();
 FILLCELL_X2 FILLER_76_680 ();
 FILLCELL_X8 FILLER_76_690 ();
 FILLCELL_X4 FILLER_76_698 ();
 FILLCELL_X2 FILLER_76_702 ();
 FILLCELL_X2 FILLER_76_780 ();
 FILLCELL_X1 FILLER_76_786 ();
 FILLCELL_X2 FILLER_76_827 ();
 FILLCELL_X4 FILLER_76_841 ();
 FILLCELL_X2 FILLER_76_845 ();
 FILLCELL_X1 FILLER_76_847 ();
 FILLCELL_X8 FILLER_76_861 ();
 FILLCELL_X4 FILLER_76_869 ();
 FILLCELL_X1 FILLER_76_873 ();
 FILLCELL_X4 FILLER_76_891 ();
 FILLCELL_X1 FILLER_76_895 ();
 FILLCELL_X4 FILLER_76_930 ();
 FILLCELL_X2 FILLER_76_934 ();
 FILLCELL_X1 FILLER_76_936 ();
 FILLCELL_X4 FILLER_76_940 ();
 FILLCELL_X2 FILLER_76_944 ();
 FILLCELL_X1 FILLER_76_946 ();
 FILLCELL_X1 FILLER_76_953 ();
 FILLCELL_X2 FILLER_76_992 ();
 FILLCELL_X1 FILLER_76_1009 ();
 FILLCELL_X2 FILLER_76_1019 ();
 FILLCELL_X2 FILLER_76_1051 ();
 FILLCELL_X1 FILLER_76_1053 ();
 FILLCELL_X8 FILLER_76_1061 ();
 FILLCELL_X4 FILLER_76_1069 ();
 FILLCELL_X1 FILLER_76_1073 ();
 FILLCELL_X8 FILLER_76_1096 ();
 FILLCELL_X4 FILLER_76_1104 ();
 FILLCELL_X2 FILLER_76_1108 ();
 FILLCELL_X1 FILLER_76_1110 ();
 FILLCELL_X16 FILLER_76_1133 ();
 FILLCELL_X2 FILLER_76_1160 ();
 FILLCELL_X1 FILLER_76_1162 ();
 FILLCELL_X4 FILLER_76_1170 ();
 FILLCELL_X1 FILLER_76_1174 ();
 FILLCELL_X2 FILLER_76_1184 ();
 FILLCELL_X4 FILLER_76_1195 ();
 FILLCELL_X1 FILLER_76_1199 ();
 FILLCELL_X4 FILLER_76_1271 ();
 FILLCELL_X2 FILLER_76_1275 ();
 FILLCELL_X2 FILLER_76_1302 ();
 FILLCELL_X8 FILLER_76_1311 ();
 FILLCELL_X2 FILLER_76_1319 ();
 FILLCELL_X4 FILLER_76_1348 ();
 FILLCELL_X1 FILLER_76_1359 ();
 FILLCELL_X2 FILLER_76_1385 ();
 FILLCELL_X1 FILLER_76_1387 ();
 FILLCELL_X16 FILLER_76_1408 ();
 FILLCELL_X1 FILLER_76_1424 ();
 FILLCELL_X4 FILLER_76_1434 ();
 FILLCELL_X2 FILLER_76_1438 ();
 FILLCELL_X1 FILLER_76_1449 ();
 FILLCELL_X1 FILLER_76_1454 ();
 FILLCELL_X4 FILLER_76_1464 ();
 FILLCELL_X2 FILLER_76_1468 ();
 FILLCELL_X2 FILLER_76_1502 ();
 FILLCELL_X1 FILLER_76_1527 ();
 FILLCELL_X2 FILLER_76_1532 ();
 FILLCELL_X2 FILLER_76_1538 ();
 FILLCELL_X1 FILLER_76_1540 ();
 FILLCELL_X4 FILLER_76_1566 ();
 FILLCELL_X2 FILLER_76_1570 ();
 FILLCELL_X4 FILLER_76_1583 ();
 FILLCELL_X2 FILLER_76_1603 ();
 FILLCELL_X1 FILLER_76_1605 ();
 FILLCELL_X8 FILLER_76_1609 ();
 FILLCELL_X4 FILLER_76_1620 ();
 FILLCELL_X2 FILLER_76_1624 ();
 FILLCELL_X1 FILLER_76_1629 ();
 FILLCELL_X16 FILLER_76_1634 ();
 FILLCELL_X1 FILLER_76_1650 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X16 FILLER_77_97 ();
 FILLCELL_X8 FILLER_77_113 ();
 FILLCELL_X1 FILLER_77_121 ();
 FILLCELL_X2 FILLER_77_169 ();
 FILLCELL_X1 FILLER_77_171 ();
 FILLCELL_X1 FILLER_77_186 ();
 FILLCELL_X4 FILLER_77_211 ();
 FILLCELL_X2 FILLER_77_215 ();
 FILLCELL_X1 FILLER_77_237 ();
 FILLCELL_X4 FILLER_77_268 ();
 FILLCELL_X2 FILLER_77_272 ();
 FILLCELL_X4 FILLER_77_278 ();
 FILLCELL_X2 FILLER_77_282 ();
 FILLCELL_X1 FILLER_77_284 ();
 FILLCELL_X4 FILLER_77_301 ();
 FILLCELL_X2 FILLER_77_305 ();
 FILLCELL_X1 FILLER_77_307 ();
 FILLCELL_X16 FILLER_77_315 ();
 FILLCELL_X4 FILLER_77_331 ();
 FILLCELL_X2 FILLER_77_335 ();
 FILLCELL_X1 FILLER_77_337 ();
 FILLCELL_X1 FILLER_77_351 ();
 FILLCELL_X2 FILLER_77_379 ();
 FILLCELL_X1 FILLER_77_381 ();
 FILLCELL_X8 FILLER_77_389 ();
 FILLCELL_X16 FILLER_77_402 ();
 FILLCELL_X1 FILLER_77_418 ();
 FILLCELL_X8 FILLER_77_426 ();
 FILLCELL_X4 FILLER_77_434 ();
 FILLCELL_X2 FILLER_77_438 ();
 FILLCELL_X1 FILLER_77_440 ();
 FILLCELL_X1 FILLER_77_496 ();
 FILLCELL_X8 FILLER_77_501 ();
 FILLCELL_X4 FILLER_77_509 ();
 FILLCELL_X2 FILLER_77_513 ();
 FILLCELL_X1 FILLER_77_515 ();
 FILLCELL_X8 FILLER_77_522 ();
 FILLCELL_X2 FILLER_77_530 ();
 FILLCELL_X16 FILLER_77_536 ();
 FILLCELL_X4 FILLER_77_572 ();
 FILLCELL_X1 FILLER_77_576 ();
 FILLCELL_X2 FILLER_77_593 ();
 FILLCELL_X8 FILLER_77_615 ();
 FILLCELL_X4 FILLER_77_652 ();
 FILLCELL_X2 FILLER_77_666 ();
 FILLCELL_X2 FILLER_77_694 ();
 FILLCELL_X2 FILLER_77_717 ();
 FILLCELL_X4 FILLER_77_726 ();
 FILLCELL_X2 FILLER_77_730 ();
 FILLCELL_X4 FILLER_77_742 ();
 FILLCELL_X2 FILLER_77_746 ();
 FILLCELL_X4 FILLER_77_752 ();
 FILLCELL_X2 FILLER_77_756 ();
 FILLCELL_X1 FILLER_77_758 ();
 FILLCELL_X1 FILLER_77_764 ();
 FILLCELL_X2 FILLER_77_785 ();
 FILLCELL_X2 FILLER_77_793 ();
 FILLCELL_X32 FILLER_77_798 ();
 FILLCELL_X32 FILLER_77_830 ();
 FILLCELL_X16 FILLER_77_862 ();
 FILLCELL_X2 FILLER_77_878 ();
 FILLCELL_X1 FILLER_77_880 ();
 FILLCELL_X4 FILLER_77_901 ();
 FILLCELL_X2 FILLER_77_905 ();
 FILLCELL_X1 FILLER_77_907 ();
 FILLCELL_X8 FILLER_77_910 ();
 FILLCELL_X1 FILLER_77_918 ();
 FILLCELL_X8 FILLER_77_923 ();
 FILLCELL_X4 FILLER_77_931 ();
 FILLCELL_X8 FILLER_77_940 ();
 FILLCELL_X4 FILLER_77_948 ();
 FILLCELL_X2 FILLER_77_952 ();
 FILLCELL_X1 FILLER_77_954 ();
 FILLCELL_X32 FILLER_77_962 ();
 FILLCELL_X4 FILLER_77_1003 ();
 FILLCELL_X1 FILLER_77_1007 ();
 FILLCELL_X2 FILLER_77_1021 ();
 FILLCELL_X16 FILLER_77_1033 ();
 FILLCELL_X2 FILLER_77_1049 ();
 FILLCELL_X4 FILLER_77_1084 ();
 FILLCELL_X4 FILLER_77_1097 ();
 FILLCELL_X1 FILLER_77_1101 ();
 FILLCELL_X4 FILLER_77_1106 ();
 FILLCELL_X8 FILLER_77_1126 ();
 FILLCELL_X4 FILLER_77_1134 ();
 FILLCELL_X1 FILLER_77_1138 ();
 FILLCELL_X2 FILLER_77_1172 ();
 FILLCELL_X1 FILLER_77_1174 ();
 FILLCELL_X4 FILLER_77_1207 ();
 FILLCELL_X1 FILLER_77_1211 ();
 FILLCELL_X4 FILLER_77_1233 ();
 FILLCELL_X1 FILLER_77_1237 ();
 FILLCELL_X16 FILLER_77_1264 ();
 FILLCELL_X4 FILLER_77_1280 ();
 FILLCELL_X2 FILLER_77_1284 ();
 FILLCELL_X1 FILLER_77_1286 ();
 FILLCELL_X2 FILLER_77_1307 ();
 FILLCELL_X1 FILLER_77_1309 ();
 FILLCELL_X1 FILLER_77_1337 ();
 FILLCELL_X4 FILLER_77_1345 ();
 FILLCELL_X4 FILLER_77_1376 ();
 FILLCELL_X1 FILLER_77_1380 ();
 FILLCELL_X2 FILLER_77_1388 ();
 FILLCELL_X1 FILLER_77_1390 ();
 FILLCELL_X4 FILLER_77_1411 ();
 FILLCELL_X4 FILLER_77_1424 ();
 FILLCELL_X2 FILLER_77_1428 ();
 FILLCELL_X4 FILLER_77_1435 ();
 FILLCELL_X2 FILLER_77_1439 ();
 FILLCELL_X1 FILLER_77_1441 ();
 FILLCELL_X1 FILLER_77_1451 ();
 FILLCELL_X2 FILLER_77_1456 ();
 FILLCELL_X1 FILLER_77_1458 ();
 FILLCELL_X4 FILLER_77_1483 ();
 FILLCELL_X4 FILLER_77_1494 ();
 FILLCELL_X2 FILLER_77_1501 ();
 FILLCELL_X1 FILLER_77_1503 ();
 FILLCELL_X1 FILLER_77_1515 ();
 FILLCELL_X2 FILLER_77_1520 ();
 FILLCELL_X1 FILLER_77_1531 ();
 FILLCELL_X2 FILLER_77_1536 ();
 FILLCELL_X1 FILLER_77_1542 ();
 FILLCELL_X4 FILLER_77_1558 ();
 FILLCELL_X2 FILLER_77_1570 ();
 FILLCELL_X1 FILLER_77_1572 ();
 FILLCELL_X8 FILLER_77_1576 ();
 FILLCELL_X2 FILLER_77_1584 ();
 FILLCELL_X8 FILLER_77_1590 ();
 FILLCELL_X4 FILLER_77_1598 ();
 FILLCELL_X2 FILLER_77_1602 ();
 FILLCELL_X1 FILLER_77_1604 ();
 FILLCELL_X4 FILLER_77_1619 ();
 FILLCELL_X2 FILLER_77_1623 ();
 FILLCELL_X16 FILLER_77_1631 ();
 FILLCELL_X4 FILLER_77_1647 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X16 FILLER_78_97 ();
 FILLCELL_X8 FILLER_78_113 ();
 FILLCELL_X4 FILLER_78_121 ();
 FILLCELL_X2 FILLER_78_125 ();
 FILLCELL_X1 FILLER_78_127 ();
 FILLCELL_X4 FILLER_78_142 ();
 FILLCELL_X2 FILLER_78_146 ();
 FILLCELL_X1 FILLER_78_148 ();
 FILLCELL_X8 FILLER_78_156 ();
 FILLCELL_X2 FILLER_78_164 ();
 FILLCELL_X1 FILLER_78_195 ();
 FILLCELL_X2 FILLER_78_216 ();
 FILLCELL_X1 FILLER_78_225 ();
 FILLCELL_X1 FILLER_78_241 ();
 FILLCELL_X1 FILLER_78_244 ();
 FILLCELL_X2 FILLER_78_249 ();
 FILLCELL_X1 FILLER_78_251 ();
 FILLCELL_X8 FILLER_78_303 ();
 FILLCELL_X2 FILLER_78_311 ();
 FILLCELL_X8 FILLER_78_327 ();
 FILLCELL_X2 FILLER_78_344 ();
 FILLCELL_X1 FILLER_78_346 ();
 FILLCELL_X8 FILLER_78_384 ();
 FILLCELL_X4 FILLER_78_392 ();
 FILLCELL_X4 FILLER_78_417 ();
 FILLCELL_X2 FILLER_78_421 ();
 FILLCELL_X16 FILLER_78_443 ();
 FILLCELL_X2 FILLER_78_459 ();
 FILLCELL_X1 FILLER_78_473 ();
 FILLCELL_X1 FILLER_78_480 ();
 FILLCELL_X1 FILLER_78_485 ();
 FILLCELL_X2 FILLER_78_506 ();
 FILLCELL_X4 FILLER_78_535 ();
 FILLCELL_X2 FILLER_78_539 ();
 FILLCELL_X8 FILLER_78_545 ();
 FILLCELL_X4 FILLER_78_553 ();
 FILLCELL_X1 FILLER_78_557 ();
 FILLCELL_X1 FILLER_78_565 ();
 FILLCELL_X2 FILLER_78_586 ();
 FILLCELL_X16 FILLER_78_615 ();
 FILLCELL_X2 FILLER_78_673 ();
 FILLCELL_X1 FILLER_78_678 ();
 FILLCELL_X4 FILLER_78_697 ();
 FILLCELL_X4 FILLER_78_704 ();
 FILLCELL_X2 FILLER_78_708 ();
 FILLCELL_X1 FILLER_78_723 ();
 FILLCELL_X4 FILLER_78_731 ();
 FILLCELL_X8 FILLER_78_740 ();
 FILLCELL_X2 FILLER_78_748 ();
 FILLCELL_X1 FILLER_78_750 ();
 FILLCELL_X2 FILLER_78_758 ();
 FILLCELL_X4 FILLER_78_762 ();
 FILLCELL_X8 FILLER_78_782 ();
 FILLCELL_X4 FILLER_78_790 ();
 FILLCELL_X2 FILLER_78_794 ();
 FILLCELL_X1 FILLER_78_796 ();
 FILLCELL_X1 FILLER_78_804 ();
 FILLCELL_X32 FILLER_78_845 ();
 FILLCELL_X16 FILLER_78_877 ();
 FILLCELL_X8 FILLER_78_893 ();
 FILLCELL_X4 FILLER_78_901 ();
 FILLCELL_X2 FILLER_78_905 ();
 FILLCELL_X1 FILLER_78_907 ();
 FILLCELL_X8 FILLER_78_913 ();
 FILLCELL_X1 FILLER_78_921 ();
 FILLCELL_X4 FILLER_78_925 ();
 FILLCELL_X1 FILLER_78_932 ();
 FILLCELL_X1 FILLER_78_937 ();
 FILLCELL_X1 FILLER_78_958 ();
 FILLCELL_X4 FILLER_78_967 ();
 FILLCELL_X1 FILLER_78_971 ();
 FILLCELL_X1 FILLER_78_987 ();
 FILLCELL_X8 FILLER_78_990 ();
 FILLCELL_X2 FILLER_78_1005 ();
 FILLCELL_X1 FILLER_78_1013 ();
 FILLCELL_X8 FILLER_78_1023 ();
 FILLCELL_X2 FILLER_78_1031 ();
 FILLCELL_X4 FILLER_78_1049 ();
 FILLCELL_X4 FILLER_78_1059 ();
 FILLCELL_X1 FILLER_78_1063 ();
 FILLCELL_X2 FILLER_78_1093 ();
 FILLCELL_X2 FILLER_78_1101 ();
 FILLCELL_X1 FILLER_78_1103 ();
 FILLCELL_X1 FILLER_78_1122 ();
 FILLCELL_X4 FILLER_78_1139 ();
 FILLCELL_X1 FILLER_78_1143 ();
 FILLCELL_X16 FILLER_78_1153 ();
 FILLCELL_X4 FILLER_78_1169 ();
 FILLCELL_X2 FILLER_78_1173 ();
 FILLCELL_X1 FILLER_78_1175 ();
 FILLCELL_X2 FILLER_78_1185 ();
 FILLCELL_X1 FILLER_78_1203 ();
 FILLCELL_X16 FILLER_78_1211 ();
 FILLCELL_X2 FILLER_78_1227 ();
 FILLCELL_X2 FILLER_78_1232 ();
 FILLCELL_X2 FILLER_78_1241 ();
 FILLCELL_X4 FILLER_78_1263 ();
 FILLCELL_X8 FILLER_78_1287 ();
 FILLCELL_X4 FILLER_78_1295 ();
 FILLCELL_X2 FILLER_78_1299 ();
 FILLCELL_X1 FILLER_78_1328 ();
 FILLCELL_X1 FILLER_78_1336 ();
 FILLCELL_X1 FILLER_78_1357 ();
 FILLCELL_X32 FILLER_78_1378 ();
 FILLCELL_X8 FILLER_78_1410 ();
 FILLCELL_X2 FILLER_78_1418 ();
 FILLCELL_X1 FILLER_78_1420 ();
 FILLCELL_X4 FILLER_78_1426 ();
 FILLCELL_X8 FILLER_78_1437 ();
 FILLCELL_X4 FILLER_78_1445 ();
 FILLCELL_X1 FILLER_78_1449 ();
 FILLCELL_X2 FILLER_78_1470 ();
 FILLCELL_X4 FILLER_78_1489 ();
 FILLCELL_X1 FILLER_78_1493 ();
 FILLCELL_X8 FILLER_78_1499 ();
 FILLCELL_X2 FILLER_78_1507 ();
 FILLCELL_X1 FILLER_78_1509 ();
 FILLCELL_X2 FILLER_78_1513 ();
 FILLCELL_X1 FILLER_78_1515 ();
 FILLCELL_X4 FILLER_78_1520 ();
 FILLCELL_X1 FILLER_78_1535 ();
 FILLCELL_X2 FILLER_78_1542 ();
 FILLCELL_X4 FILLER_78_1547 ();
 FILLCELL_X2 FILLER_78_1551 ();
 FILLCELL_X1 FILLER_78_1553 ();
 FILLCELL_X2 FILLER_78_1559 ();
 FILLCELL_X4 FILLER_78_1587 ();
 FILLCELL_X8 FILLER_78_1595 ();
 FILLCELL_X4 FILLER_78_1603 ();
 FILLCELL_X2 FILLER_78_1611 ();
 FILLCELL_X1 FILLER_78_1613 ();
 FILLCELL_X16 FILLER_78_1617 ();
 FILLCELL_X2 FILLER_78_1633 ();
 FILLCELL_X1 FILLER_78_1641 ();
 FILLCELL_X2 FILLER_78_1648 ();
 FILLCELL_X1 FILLER_78_1650 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X8 FILLER_79_129 ();
 FILLCELL_X4 FILLER_79_137 ();
 FILLCELL_X2 FILLER_79_161 ();
 FILLCELL_X8 FILLER_79_170 ();
 FILLCELL_X4 FILLER_79_178 ();
 FILLCELL_X1 FILLER_79_182 ();
 FILLCELL_X16 FILLER_79_185 ();
 FILLCELL_X4 FILLER_79_201 ();
 FILLCELL_X2 FILLER_79_205 ();
 FILLCELL_X1 FILLER_79_207 ();
 FILLCELL_X2 FILLER_79_213 ();
 FILLCELL_X1 FILLER_79_215 ();
 FILLCELL_X4 FILLER_79_220 ();
 FILLCELL_X2 FILLER_79_224 ();
 FILLCELL_X2 FILLER_79_233 ();
 FILLCELL_X1 FILLER_79_235 ();
 FILLCELL_X1 FILLER_79_253 ();
 FILLCELL_X2 FILLER_79_258 ();
 FILLCELL_X2 FILLER_79_263 ();
 FILLCELL_X1 FILLER_79_265 ();
 FILLCELL_X4 FILLER_79_273 ();
 FILLCELL_X2 FILLER_79_277 ();
 FILLCELL_X1 FILLER_79_282 ();
 FILLCELL_X1 FILLER_79_287 ();
 FILLCELL_X1 FILLER_79_292 ();
 FILLCELL_X1 FILLER_79_304 ();
 FILLCELL_X2 FILLER_79_308 ();
 FILLCELL_X1 FILLER_79_317 ();
 FILLCELL_X2 FILLER_79_322 ();
 FILLCELL_X4 FILLER_79_338 ();
 FILLCELL_X1 FILLER_79_342 ();
 FILLCELL_X4 FILLER_79_360 ();
 FILLCELL_X2 FILLER_79_364 ();
 FILLCELL_X1 FILLER_79_396 ();
 FILLCELL_X4 FILLER_79_404 ();
 FILLCELL_X1 FILLER_79_408 ();
 FILLCELL_X4 FILLER_79_429 ();
 FILLCELL_X2 FILLER_79_467 ();
 FILLCELL_X1 FILLER_79_480 ();
 FILLCELL_X2 FILLER_79_485 ();
 FILLCELL_X2 FILLER_79_501 ();
 FILLCELL_X16 FILLER_79_505 ();
 FILLCELL_X4 FILLER_79_521 ();
 FILLCELL_X4 FILLER_79_547 ();
 FILLCELL_X2 FILLER_79_551 ();
 FILLCELL_X1 FILLER_79_553 ();
 FILLCELL_X1 FILLER_79_567 ();
 FILLCELL_X1 FILLER_79_575 ();
 FILLCELL_X1 FILLER_79_603 ();
 FILLCELL_X4 FILLER_79_614 ();
 FILLCELL_X2 FILLER_79_618 ();
 FILLCELL_X1 FILLER_79_620 ();
 FILLCELL_X4 FILLER_79_630 ();
 FILLCELL_X2 FILLER_79_634 ();
 FILLCELL_X1 FILLER_79_636 ();
 FILLCELL_X8 FILLER_79_644 ();
 FILLCELL_X4 FILLER_79_652 ();
 FILLCELL_X16 FILLER_79_663 ();
 FILLCELL_X1 FILLER_79_679 ();
 FILLCELL_X8 FILLER_79_686 ();
 FILLCELL_X4 FILLER_79_694 ();
 FILLCELL_X2 FILLER_79_698 ();
 FILLCELL_X1 FILLER_79_709 ();
 FILLCELL_X2 FILLER_79_714 ();
 FILLCELL_X2 FILLER_79_721 ();
 FILLCELL_X1 FILLER_79_723 ();
 FILLCELL_X4 FILLER_79_726 ();
 FILLCELL_X1 FILLER_79_730 ();
 FILLCELL_X1 FILLER_79_758 ();
 FILLCELL_X8 FILLER_79_779 ();
 FILLCELL_X4 FILLER_79_787 ();
 FILLCELL_X2 FILLER_79_791 ();
 FILLCELL_X8 FILLER_79_816 ();
 FILLCELL_X2 FILLER_79_824 ();
 FILLCELL_X1 FILLER_79_826 ();
 FILLCELL_X8 FILLER_79_831 ();
 FILLCELL_X2 FILLER_79_839 ();
 FILLCELL_X4 FILLER_79_863 ();
 FILLCELL_X2 FILLER_79_867 ();
 FILLCELL_X1 FILLER_79_869 ();
 FILLCELL_X8 FILLER_79_892 ();
 FILLCELL_X2 FILLER_79_900 ();
 FILLCELL_X2 FILLER_79_909 ();
 FILLCELL_X4 FILLER_79_915 ();
 FILLCELL_X4 FILLER_79_939 ();
 FILLCELL_X1 FILLER_79_954 ();
 FILLCELL_X16 FILLER_79_959 ();
 FILLCELL_X4 FILLER_79_975 ();
 FILLCELL_X2 FILLER_79_979 ();
 FILLCELL_X1 FILLER_79_981 ();
 FILLCELL_X16 FILLER_79_1012 ();
 FILLCELL_X4 FILLER_79_1028 ();
 FILLCELL_X1 FILLER_79_1038 ();
 FILLCELL_X8 FILLER_79_1045 ();
 FILLCELL_X4 FILLER_79_1065 ();
 FILLCELL_X2 FILLER_79_1069 ();
 FILLCELL_X4 FILLER_79_1084 ();
 FILLCELL_X2 FILLER_79_1095 ();
 FILLCELL_X1 FILLER_79_1097 ();
 FILLCELL_X2 FILLER_79_1105 ();
 FILLCELL_X2 FILLER_79_1110 ();
 FILLCELL_X1 FILLER_79_1112 ();
 FILLCELL_X2 FILLER_79_1123 ();
 FILLCELL_X1 FILLER_79_1125 ();
 FILLCELL_X1 FILLER_79_1135 ();
 FILLCELL_X8 FILLER_79_1169 ();
 FILLCELL_X8 FILLER_79_1195 ();
 FILLCELL_X4 FILLER_79_1203 ();
 FILLCELL_X4 FILLER_79_1213 ();
 FILLCELL_X2 FILLER_79_1217 ();
 FILLCELL_X1 FILLER_79_1219 ();
 FILLCELL_X2 FILLER_79_1234 ();
 FILLCELL_X2 FILLER_79_1239 ();
 FILLCELL_X2 FILLER_79_1248 ();
 FILLCELL_X16 FILLER_79_1264 ();
 FILLCELL_X4 FILLER_79_1287 ();
 FILLCELL_X1 FILLER_79_1291 ();
 FILLCELL_X2 FILLER_79_1306 ();
 FILLCELL_X1 FILLER_79_1308 ();
 FILLCELL_X2 FILLER_79_1316 ();
 FILLCELL_X8 FILLER_79_1338 ();
 FILLCELL_X8 FILLER_79_1353 ();
 FILLCELL_X4 FILLER_79_1381 ();
 FILLCELL_X1 FILLER_79_1385 ();
 FILLCELL_X32 FILLER_79_1406 ();
 FILLCELL_X1 FILLER_79_1438 ();
 FILLCELL_X1 FILLER_79_1455 ();
 FILLCELL_X4 FILLER_79_1465 ();
 FILLCELL_X2 FILLER_79_1469 ();
 FILLCELL_X1 FILLER_79_1487 ();
 FILLCELL_X2 FILLER_79_1492 ();
 FILLCELL_X2 FILLER_79_1526 ();
 FILLCELL_X1 FILLER_79_1533 ();
 FILLCELL_X1 FILLER_79_1538 ();
 FILLCELL_X2 FILLER_79_1543 ();
 FILLCELL_X2 FILLER_79_1550 ();
 FILLCELL_X1 FILLER_79_1552 ();
 FILLCELL_X2 FILLER_79_1564 ();
 FILLCELL_X1 FILLER_79_1566 ();
 FILLCELL_X8 FILLER_79_1588 ();
 FILLCELL_X4 FILLER_79_1596 ();
 FILLCELL_X1 FILLER_79_1604 ();
 FILLCELL_X4 FILLER_79_1617 ();
 FILLCELL_X1 FILLER_79_1621 ();
 FILLCELL_X4 FILLER_79_1627 ();
 FILLCELL_X2 FILLER_79_1631 ();
 FILLCELL_X1 FILLER_79_1633 ();
 FILLCELL_X2 FILLER_79_1637 ();
 FILLCELL_X1 FILLER_79_1639 ();
 FILLCELL_X2 FILLER_79_1648 ();
 FILLCELL_X1 FILLER_79_1650 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X16 FILLER_80_97 ();
 FILLCELL_X8 FILLER_80_113 ();
 FILLCELL_X4 FILLER_80_121 ();
 FILLCELL_X2 FILLER_80_125 ();
 FILLCELL_X1 FILLER_80_127 ();
 FILLCELL_X8 FILLER_80_158 ();
 FILLCELL_X1 FILLER_80_186 ();
 FILLCELL_X1 FILLER_80_207 ();
 FILLCELL_X1 FILLER_80_212 ();
 FILLCELL_X1 FILLER_80_216 ();
 FILLCELL_X1 FILLER_80_224 ();
 FILLCELL_X2 FILLER_80_229 ();
 FILLCELL_X4 FILLER_80_238 ();
 FILLCELL_X2 FILLER_80_281 ();
 FILLCELL_X4 FILLER_80_294 ();
 FILLCELL_X2 FILLER_80_300 ();
 FILLCELL_X1 FILLER_80_302 ();
 FILLCELL_X8 FILLER_80_308 ();
 FILLCELL_X2 FILLER_80_316 ();
 FILLCELL_X2 FILLER_80_321 ();
 FILLCELL_X2 FILLER_80_330 ();
 FILLCELL_X1 FILLER_80_357 ();
 FILLCELL_X2 FILLER_80_365 ();
 FILLCELL_X1 FILLER_80_367 ();
 FILLCELL_X1 FILLER_80_374 ();
 FILLCELL_X4 FILLER_80_409 ();
 FILLCELL_X2 FILLER_80_413 ();
 FILLCELL_X1 FILLER_80_415 ();
 FILLCELL_X1 FILLER_80_419 ();
 FILLCELL_X8 FILLER_80_425 ();
 FILLCELL_X2 FILLER_80_433 ();
 FILLCELL_X1 FILLER_80_442 ();
 FILLCELL_X1 FILLER_80_452 ();
 FILLCELL_X1 FILLER_80_464 ();
 FILLCELL_X1 FILLER_80_469 ();
 FILLCELL_X1 FILLER_80_474 ();
 FILLCELL_X2 FILLER_80_498 ();
 FILLCELL_X16 FILLER_80_504 ();
 FILLCELL_X4 FILLER_80_520 ();
 FILLCELL_X2 FILLER_80_524 ();
 FILLCELL_X8 FILLER_80_541 ();
 FILLCELL_X1 FILLER_80_549 ();
 FILLCELL_X2 FILLER_80_578 ();
 FILLCELL_X4 FILLER_80_593 ();
 FILLCELL_X4 FILLER_80_600 ();
 FILLCELL_X1 FILLER_80_604 ();
 FILLCELL_X8 FILLER_80_622 ();
 FILLCELL_X1 FILLER_80_630 ();
 FILLCELL_X4 FILLER_80_632 ();
 FILLCELL_X1 FILLER_80_636 ();
 FILLCELL_X8 FILLER_80_652 ();
 FILLCELL_X2 FILLER_80_691 ();
 FILLCELL_X2 FILLER_80_703 ();
 FILLCELL_X1 FILLER_80_715 ();
 FILLCELL_X8 FILLER_80_744 ();
 FILLCELL_X1 FILLER_80_752 ();
 FILLCELL_X4 FILLER_80_789 ();
 FILLCELL_X2 FILLER_80_793 ();
 FILLCELL_X2 FILLER_80_835 ();
 FILLCELL_X1 FILLER_80_837 ();
 FILLCELL_X16 FILLER_80_845 ();
 FILLCELL_X2 FILLER_80_861 ();
 FILLCELL_X1 FILLER_80_870 ();
 FILLCELL_X1 FILLER_80_883 ();
 FILLCELL_X8 FILLER_80_906 ();
 FILLCELL_X2 FILLER_80_914 ();
 FILLCELL_X16 FILLER_80_920 ();
 FILLCELL_X8 FILLER_80_936 ();
 FILLCELL_X2 FILLER_80_944 ();
 FILLCELL_X4 FILLER_80_956 ();
 FILLCELL_X2 FILLER_80_960 ();
 FILLCELL_X1 FILLER_80_962 ();
 FILLCELL_X2 FILLER_80_968 ();
 FILLCELL_X16 FILLER_80_980 ();
 FILLCELL_X2 FILLER_80_996 ();
 FILLCELL_X1 FILLER_80_998 ();
 FILLCELL_X8 FILLER_80_1004 ();
 FILLCELL_X4 FILLER_80_1012 ();
 FILLCELL_X8 FILLER_80_1023 ();
 FILLCELL_X1 FILLER_80_1031 ();
 FILLCELL_X4 FILLER_80_1042 ();
 FILLCELL_X2 FILLER_80_1046 ();
 FILLCELL_X2 FILLER_80_1055 ();
 FILLCELL_X1 FILLER_80_1057 ();
 FILLCELL_X4 FILLER_80_1062 ();
 FILLCELL_X4 FILLER_80_1076 ();
 FILLCELL_X2 FILLER_80_1080 ();
 FILLCELL_X1 FILLER_80_1082 ();
 FILLCELL_X8 FILLER_80_1115 ();
 FILLCELL_X4 FILLER_80_1123 ();
 FILLCELL_X8 FILLER_80_1133 ();
 FILLCELL_X4 FILLER_80_1141 ();
 FILLCELL_X2 FILLER_80_1145 ();
 FILLCELL_X1 FILLER_80_1147 ();
 FILLCELL_X32 FILLER_80_1150 ();
 FILLCELL_X16 FILLER_80_1182 ();
 FILLCELL_X1 FILLER_80_1198 ();
 FILLCELL_X1 FILLER_80_1206 ();
 FILLCELL_X2 FILLER_80_1210 ();
 FILLCELL_X8 FILLER_80_1269 ();
 FILLCELL_X4 FILLER_80_1277 ();
 FILLCELL_X1 FILLER_80_1281 ();
 FILLCELL_X16 FILLER_80_1316 ();
 FILLCELL_X8 FILLER_80_1332 ();
 FILLCELL_X2 FILLER_80_1340 ();
 FILLCELL_X16 FILLER_80_1352 ();
 FILLCELL_X1 FILLER_80_1368 ();
 FILLCELL_X16 FILLER_80_1389 ();
 FILLCELL_X4 FILLER_80_1405 ();
 FILLCELL_X1 FILLER_80_1409 ();
 FILLCELL_X4 FILLER_80_1429 ();
 FILLCELL_X2 FILLER_80_1433 ();
 FILLCELL_X1 FILLER_80_1435 ();
 FILLCELL_X2 FILLER_80_1468 ();
 FILLCELL_X2 FILLER_80_1474 ();
 FILLCELL_X2 FILLER_80_1493 ();
 FILLCELL_X2 FILLER_80_1502 ();
 FILLCELL_X1 FILLER_80_1504 ();
 FILLCELL_X4 FILLER_80_1508 ();
 FILLCELL_X2 FILLER_80_1512 ();
 FILLCELL_X4 FILLER_80_1529 ();
 FILLCELL_X2 FILLER_80_1533 ();
 FILLCELL_X2 FILLER_80_1539 ();
 FILLCELL_X1 FILLER_80_1541 ();
 FILLCELL_X4 FILLER_80_1574 ();
 FILLCELL_X2 FILLER_80_1578 ();
 FILLCELL_X4 FILLER_80_1594 ();
 FILLCELL_X2 FILLER_80_1598 ();
 FILLCELL_X1 FILLER_80_1600 ();
 FILLCELL_X1 FILLER_80_1609 ();
 FILLCELL_X16 FILLER_80_1614 ();
 FILLCELL_X8 FILLER_80_1630 ();
 FILLCELL_X2 FILLER_80_1638 ();
 FILLCELL_X1 FILLER_80_1640 ();
 FILLCELL_X4 FILLER_80_1644 ();
 FILLCELL_X2 FILLER_80_1648 ();
 FILLCELL_X1 FILLER_80_1650 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X16 FILLER_81_129 ();
 FILLCELL_X2 FILLER_81_145 ();
 FILLCELL_X1 FILLER_81_147 ();
 FILLCELL_X4 FILLER_81_180 ();
 FILLCELL_X2 FILLER_81_184 ();
 FILLCELL_X1 FILLER_81_186 ();
 FILLCELL_X2 FILLER_81_222 ();
 FILLCELL_X1 FILLER_81_224 ();
 FILLCELL_X2 FILLER_81_230 ();
 FILLCELL_X1 FILLER_81_232 ();
 FILLCELL_X2 FILLER_81_239 ();
 FILLCELL_X1 FILLER_81_241 ();
 FILLCELL_X2 FILLER_81_262 ();
 FILLCELL_X4 FILLER_81_294 ();
 FILLCELL_X1 FILLER_81_304 ();
 FILLCELL_X2 FILLER_81_310 ();
 FILLCELL_X1 FILLER_81_339 ();
 FILLCELL_X2 FILLER_81_380 ();
 FILLCELL_X1 FILLER_81_396 ();
 FILLCELL_X1 FILLER_81_436 ();
 FILLCELL_X2 FILLER_81_444 ();
 FILLCELL_X1 FILLER_81_446 ();
 FILLCELL_X2 FILLER_81_465 ();
 FILLCELL_X1 FILLER_81_467 ();
 FILLCELL_X4 FILLER_81_481 ();
 FILLCELL_X2 FILLER_81_485 ();
 FILLCELL_X1 FILLER_81_487 ();
 FILLCELL_X4 FILLER_81_509 ();
 FILLCELL_X4 FILLER_81_519 ();
 FILLCELL_X2 FILLER_81_523 ();
 FILLCELL_X4 FILLER_81_535 ();
 FILLCELL_X4 FILLER_81_545 ();
 FILLCELL_X2 FILLER_81_562 ();
 FILLCELL_X2 FILLER_81_576 ();
 FILLCELL_X8 FILLER_81_595 ();
 FILLCELL_X2 FILLER_81_603 ();
 FILLCELL_X1 FILLER_81_620 ();
 FILLCELL_X2 FILLER_81_626 ();
 FILLCELL_X2 FILLER_81_640 ();
 FILLCELL_X1 FILLER_81_642 ();
 FILLCELL_X2 FILLER_81_690 ();
 FILLCELL_X1 FILLER_81_692 ();
 FILLCELL_X1 FILLER_81_713 ();
 FILLCELL_X4 FILLER_81_720 ();
 FILLCELL_X1 FILLER_81_724 ();
 FILLCELL_X1 FILLER_81_744 ();
 FILLCELL_X1 FILLER_81_761 ();
 FILLCELL_X8 FILLER_81_788 ();
 FILLCELL_X2 FILLER_81_796 ();
 FILLCELL_X1 FILLER_81_804 ();
 FILLCELL_X1 FILLER_81_809 ();
 FILLCELL_X1 FILLER_81_814 ();
 FILLCELL_X8 FILLER_81_830 ();
 FILLCELL_X1 FILLER_81_838 ();
 FILLCELL_X2 FILLER_81_861 ();
 FILLCELL_X1 FILLER_81_863 ();
 FILLCELL_X16 FILLER_81_893 ();
 FILLCELL_X2 FILLER_81_909 ();
 FILLCELL_X1 FILLER_81_911 ();
 FILLCELL_X16 FILLER_81_929 ();
 FILLCELL_X8 FILLER_81_945 ();
 FILLCELL_X4 FILLER_81_953 ();
 FILLCELL_X2 FILLER_81_965 ();
 FILLCELL_X1 FILLER_81_967 ();
 FILLCELL_X2 FILLER_81_975 ();
 FILLCELL_X16 FILLER_81_981 ();
 FILLCELL_X8 FILLER_81_1004 ();
 FILLCELL_X1 FILLER_81_1039 ();
 FILLCELL_X2 FILLER_81_1060 ();
 FILLCELL_X2 FILLER_81_1068 ();
 FILLCELL_X2 FILLER_81_1077 ();
 FILLCELL_X1 FILLER_81_1086 ();
 FILLCELL_X32 FILLER_81_1096 ();
 FILLCELL_X4 FILLER_81_1128 ();
 FILLCELL_X4 FILLER_81_1145 ();
 FILLCELL_X4 FILLER_81_1208 ();
 FILLCELL_X2 FILLER_81_1212 ();
 FILLCELL_X1 FILLER_81_1214 ();
 FILLCELL_X4 FILLER_81_1257 ();
 FILLCELL_X2 FILLER_81_1261 ();
 FILLCELL_X1 FILLER_81_1264 ();
 FILLCELL_X1 FILLER_81_1315 ();
 FILLCELL_X2 FILLER_81_1323 ();
 FILLCELL_X2 FILLER_81_1339 ();
 FILLCELL_X1 FILLER_81_1355 ();
 FILLCELL_X2 FILLER_81_1372 ();
 FILLCELL_X8 FILLER_81_1384 ();
 FILLCELL_X4 FILLER_81_1392 ();
 FILLCELL_X1 FILLER_81_1396 ();
 FILLCELL_X4 FILLER_81_1417 ();
 FILLCELL_X1 FILLER_81_1421 ();
 FILLCELL_X1 FILLER_81_1467 ();
 FILLCELL_X2 FILLER_81_1475 ();
 FILLCELL_X2 FILLER_81_1485 ();
 FILLCELL_X1 FILLER_81_1487 ();
 FILLCELL_X4 FILLER_81_1513 ();
 FILLCELL_X2 FILLER_81_1517 ();
 FILLCELL_X1 FILLER_81_1519 ();
 FILLCELL_X8 FILLER_81_1525 ();
 FILLCELL_X1 FILLER_81_1533 ();
 FILLCELL_X2 FILLER_81_1539 ();
 FILLCELL_X1 FILLER_81_1541 ();
 FILLCELL_X8 FILLER_81_1545 ();
 FILLCELL_X1 FILLER_81_1553 ();
 FILLCELL_X4 FILLER_81_1558 ();
 FILLCELL_X1 FILLER_81_1562 ();
 FILLCELL_X4 FILLER_81_1568 ();
 FILLCELL_X2 FILLER_81_1584 ();
 FILLCELL_X2 FILLER_81_1605 ();
 FILLCELL_X1 FILLER_81_1607 ();
 FILLCELL_X2 FILLER_81_1613 ();
 FILLCELL_X8 FILLER_81_1629 ();
 FILLCELL_X2 FILLER_81_1637 ();
 FILLCELL_X8 FILLER_81_1643 ();
 FILLCELL_X4 FILLER_82_1 ();
 FILLCELL_X2 FILLER_82_5 ();
 FILLCELL_X16 FILLER_82_11 ();
 FILLCELL_X1 FILLER_82_27 ();
 FILLCELL_X4 FILLER_82_31 ();
 FILLCELL_X1 FILLER_82_35 ();
 FILLCELL_X32 FILLER_82_39 ();
 FILLCELL_X32 FILLER_82_71 ();
 FILLCELL_X16 FILLER_82_103 ();
 FILLCELL_X8 FILLER_82_119 ();
 FILLCELL_X4 FILLER_82_127 ();
 FILLCELL_X4 FILLER_82_138 ();
 FILLCELL_X1 FILLER_82_162 ();
 FILLCELL_X1 FILLER_82_197 ();
 FILLCELL_X1 FILLER_82_234 ();
 FILLCELL_X8 FILLER_82_245 ();
 FILLCELL_X4 FILLER_82_253 ();
 FILLCELL_X2 FILLER_82_257 ();
 FILLCELL_X1 FILLER_82_274 ();
 FILLCELL_X1 FILLER_82_282 ();
 FILLCELL_X4 FILLER_82_299 ();
 FILLCELL_X8 FILLER_82_314 ();
 FILLCELL_X8 FILLER_82_332 ();
 FILLCELL_X2 FILLER_82_340 ();
 FILLCELL_X16 FILLER_82_349 ();
 FILLCELL_X4 FILLER_82_365 ();
 FILLCELL_X1 FILLER_82_369 ();
 FILLCELL_X4 FILLER_82_377 ();
 FILLCELL_X1 FILLER_82_412 ();
 FILLCELL_X1 FILLER_82_418 ();
 FILLCELL_X1 FILLER_82_427 ();
 FILLCELL_X1 FILLER_82_431 ();
 FILLCELL_X8 FILLER_82_440 ();
 FILLCELL_X32 FILLER_82_452 ();
 FILLCELL_X4 FILLER_82_484 ();
 FILLCELL_X1 FILLER_82_488 ();
 FILLCELL_X2 FILLER_82_492 ();
 FILLCELL_X1 FILLER_82_504 ();
 FILLCELL_X2 FILLER_82_525 ();
 FILLCELL_X1 FILLER_82_539 ();
 FILLCELL_X1 FILLER_82_546 ();
 FILLCELL_X1 FILLER_82_556 ();
 FILLCELL_X2 FILLER_82_560 ();
 FILLCELL_X1 FILLER_82_566 ();
 FILLCELL_X2 FILLER_82_574 ();
 FILLCELL_X1 FILLER_82_580 ();
 FILLCELL_X1 FILLER_82_588 ();
 FILLCELL_X2 FILLER_82_595 ();
 FILLCELL_X1 FILLER_82_597 ();
 FILLCELL_X4 FILLER_82_632 ();
 FILLCELL_X2 FILLER_82_636 ();
 FILLCELL_X1 FILLER_82_638 ();
 FILLCELL_X8 FILLER_82_647 ();
 FILLCELL_X2 FILLER_82_655 ();
 FILLCELL_X1 FILLER_82_657 ();
 FILLCELL_X2 FILLER_82_671 ();
 FILLCELL_X1 FILLER_82_673 ();
 FILLCELL_X16 FILLER_82_678 ();
 FILLCELL_X4 FILLER_82_694 ();
 FILLCELL_X2 FILLER_82_698 ();
 FILLCELL_X16 FILLER_82_709 ();
 FILLCELL_X4 FILLER_82_725 ();
 FILLCELL_X2 FILLER_82_729 ();
 FILLCELL_X8 FILLER_82_737 ();
 FILLCELL_X4 FILLER_82_745 ();
 FILLCELL_X2 FILLER_82_749 ();
 FILLCELL_X1 FILLER_82_751 ();
 FILLCELL_X2 FILLER_82_769 ();
 FILLCELL_X2 FILLER_82_802 ();
 FILLCELL_X4 FILLER_82_818 ();
 FILLCELL_X2 FILLER_82_822 ();
 FILLCELL_X1 FILLER_82_824 ();
 FILLCELL_X8 FILLER_82_845 ();
 FILLCELL_X4 FILLER_82_853 ();
 FILLCELL_X1 FILLER_82_857 ();
 FILLCELL_X8 FILLER_82_917 ();
 FILLCELL_X2 FILLER_82_925 ();
 FILLCELL_X1 FILLER_82_927 ();
 FILLCELL_X4 FILLER_82_932 ();
 FILLCELL_X2 FILLER_82_936 ();
 FILLCELL_X1 FILLER_82_938 ();
 FILLCELL_X1 FILLER_82_944 ();
 FILLCELL_X1 FILLER_82_952 ();
 FILLCELL_X16 FILLER_82_964 ();
 FILLCELL_X8 FILLER_82_980 ();
 FILLCELL_X4 FILLER_82_993 ();
 FILLCELL_X16 FILLER_82_1001 ();
 FILLCELL_X1 FILLER_82_1017 ();
 FILLCELL_X16 FILLER_82_1026 ();
 FILLCELL_X8 FILLER_82_1042 ();
 FILLCELL_X4 FILLER_82_1050 ();
 FILLCELL_X2 FILLER_82_1054 ();
 FILLCELL_X2 FILLER_82_1063 ();
 FILLCELL_X8 FILLER_82_1071 ();
 FILLCELL_X4 FILLER_82_1079 ();
 FILLCELL_X2 FILLER_82_1083 ();
 FILLCELL_X1 FILLER_82_1085 ();
 FILLCELL_X4 FILLER_82_1090 ();
 FILLCELL_X2 FILLER_82_1109 ();
 FILLCELL_X1 FILLER_82_1111 ();
 FILLCELL_X4 FILLER_82_1122 ();
 FILLCELL_X2 FILLER_82_1126 ();
 FILLCELL_X1 FILLER_82_1128 ();
 FILLCELL_X4 FILLER_82_1139 ();
 FILLCELL_X2 FILLER_82_1143 ();
 FILLCELL_X1 FILLER_82_1145 ();
 FILLCELL_X32 FILLER_82_1182 ();
 FILLCELL_X2 FILLER_82_1214 ();
 FILLCELL_X1 FILLER_82_1216 ();
 FILLCELL_X2 FILLER_82_1240 ();
 FILLCELL_X1 FILLER_82_1242 ();
 FILLCELL_X1 FILLER_82_1247 ();
 FILLCELL_X2 FILLER_82_1275 ();
 FILLCELL_X1 FILLER_82_1277 ();
 FILLCELL_X1 FILLER_82_1292 ();
 FILLCELL_X1 FILLER_82_1314 ();
 FILLCELL_X1 FILLER_82_1322 ();
 FILLCELL_X2 FILLER_82_1330 ();
 FILLCELL_X2 FILLER_82_1346 ();
 FILLCELL_X2 FILLER_82_1376 ();
 FILLCELL_X1 FILLER_82_1378 ();
 FILLCELL_X1 FILLER_82_1382 ();
 FILLCELL_X4 FILLER_82_1390 ();
 FILLCELL_X2 FILLER_82_1394 ();
 FILLCELL_X16 FILLER_82_1400 ();
 FILLCELL_X2 FILLER_82_1416 ();
 FILLCELL_X1 FILLER_82_1418 ();
 FILLCELL_X4 FILLER_82_1428 ();
 FILLCELL_X1 FILLER_82_1457 ();
 FILLCELL_X2 FILLER_82_1463 ();
 FILLCELL_X2 FILLER_82_1470 ();
 FILLCELL_X4 FILLER_82_1490 ();
 FILLCELL_X2 FILLER_82_1494 ();
 FILLCELL_X2 FILLER_82_1499 ();
 FILLCELL_X2 FILLER_82_1510 ();
 FILLCELL_X1 FILLER_82_1512 ();
 FILLCELL_X8 FILLER_82_1537 ();
 FILLCELL_X2 FILLER_82_1545 ();
 FILLCELL_X1 FILLER_82_1547 ();
 FILLCELL_X2 FILLER_82_1560 ();
 FILLCELL_X1 FILLER_82_1562 ();
 FILLCELL_X1 FILLER_82_1587 ();
 FILLCELL_X2 FILLER_82_1594 ();
 FILLCELL_X2 FILLER_82_1605 ();
 FILLCELL_X8 FILLER_82_1616 ();
 FILLCELL_X4 FILLER_82_1624 ();
 FILLCELL_X2 FILLER_82_1638 ();
 FILLCELL_X1 FILLER_82_1640 ();
 FILLCELL_X4 FILLER_82_1646 ();
 FILLCELL_X1 FILLER_82_1650 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X2 FILLER_83_129 ();
 FILLCELL_X1 FILLER_83_131 ();
 FILLCELL_X1 FILLER_83_159 ();
 FILLCELL_X16 FILLER_83_167 ();
 FILLCELL_X2 FILLER_83_183 ();
 FILLCELL_X4 FILLER_83_241 ();
 FILLCELL_X2 FILLER_83_245 ();
 FILLCELL_X1 FILLER_83_247 ();
 FILLCELL_X2 FILLER_83_275 ();
 FILLCELL_X1 FILLER_83_297 ();
 FILLCELL_X2 FILLER_83_323 ();
 FILLCELL_X2 FILLER_83_337 ();
 FILLCELL_X2 FILLER_83_357 ();
 FILLCELL_X1 FILLER_83_366 ();
 FILLCELL_X2 FILLER_83_371 ();
 FILLCELL_X2 FILLER_83_377 ();
 FILLCELL_X2 FILLER_83_399 ();
 FILLCELL_X1 FILLER_83_401 ();
 FILLCELL_X8 FILLER_83_408 ();
 FILLCELL_X4 FILLER_83_416 ();
 FILLCELL_X2 FILLER_83_420 ();
 FILLCELL_X2 FILLER_83_459 ();
 FILLCELL_X1 FILLER_83_464 ();
 FILLCELL_X1 FILLER_83_468 ();
 FILLCELL_X1 FILLER_83_480 ();
 FILLCELL_X1 FILLER_83_484 ();
 FILLCELL_X1 FILLER_83_495 ();
 FILLCELL_X1 FILLER_83_519 ();
 FILLCELL_X1 FILLER_83_524 ();
 FILLCELL_X1 FILLER_83_533 ();
 FILLCELL_X4 FILLER_83_548 ();
 FILLCELL_X2 FILLER_83_552 ();
 FILLCELL_X1 FILLER_83_554 ();
 FILLCELL_X8 FILLER_83_578 ();
 FILLCELL_X2 FILLER_83_586 ();
 FILLCELL_X8 FILLER_83_600 ();
 FILLCELL_X1 FILLER_83_608 ();
 FILLCELL_X2 FILLER_83_625 ();
 FILLCELL_X1 FILLER_83_627 ();
 FILLCELL_X1 FILLER_83_639 ();
 FILLCELL_X2 FILLER_83_660 ();
 FILLCELL_X2 FILLER_83_669 ();
 FILLCELL_X2 FILLER_83_678 ();
 FILLCELL_X2 FILLER_83_684 ();
 FILLCELL_X2 FILLER_83_707 ();
 FILLCELL_X8 FILLER_83_712 ();
 FILLCELL_X1 FILLER_83_720 ();
 FILLCELL_X1 FILLER_83_753 ();
 FILLCELL_X4 FILLER_83_774 ();
 FILLCELL_X8 FILLER_83_798 ();
 FILLCELL_X2 FILLER_83_813 ();
 FILLCELL_X1 FILLER_83_815 ();
 FILLCELL_X8 FILLER_83_824 ();
 FILLCELL_X2 FILLER_83_832 ();
 FILLCELL_X1 FILLER_83_863 ();
 FILLCELL_X4 FILLER_83_878 ();
 FILLCELL_X2 FILLER_83_882 ();
 FILLCELL_X1 FILLER_83_884 ();
 FILLCELL_X2 FILLER_83_927 ();
 FILLCELL_X1 FILLER_83_929 ();
 FILLCELL_X1 FILLER_83_958 ();
 FILLCELL_X16 FILLER_83_967 ();
 FILLCELL_X8 FILLER_83_983 ();
 FILLCELL_X2 FILLER_83_991 ();
 FILLCELL_X4 FILLER_83_1001 ();
 FILLCELL_X2 FILLER_83_1005 ();
 FILLCELL_X2 FILLER_83_1015 ();
 FILLCELL_X16 FILLER_83_1022 ();
 FILLCELL_X2 FILLER_83_1038 ();
 FILLCELL_X4 FILLER_83_1047 ();
 FILLCELL_X2 FILLER_83_1051 ();
 FILLCELL_X1 FILLER_83_1053 ();
 FILLCELL_X32 FILLER_83_1059 ();
 FILLCELL_X8 FILLER_83_1091 ();
 FILLCELL_X4 FILLER_83_1099 ();
 FILLCELL_X1 FILLER_83_1103 ();
 FILLCELL_X2 FILLER_83_1111 ();
 FILLCELL_X2 FILLER_83_1122 ();
 FILLCELL_X2 FILLER_83_1134 ();
 FILLCELL_X1 FILLER_83_1136 ();
 FILLCELL_X4 FILLER_83_1156 ();
 FILLCELL_X4 FILLER_83_1186 ();
 FILLCELL_X2 FILLER_83_1190 ();
 FILLCELL_X8 FILLER_83_1198 ();
 FILLCELL_X4 FILLER_83_1206 ();
 FILLCELL_X2 FILLER_83_1210 ();
 FILLCELL_X2 FILLER_83_1236 ();
 FILLCELL_X1 FILLER_83_1238 ();
 FILLCELL_X1 FILLER_83_1264 ();
 FILLCELL_X1 FILLER_83_1267 ();
 FILLCELL_X2 FILLER_83_1275 ();
 FILLCELL_X1 FILLER_83_1277 ();
 FILLCELL_X4 FILLER_83_1316 ();
 FILLCELL_X1 FILLER_83_1323 ();
 FILLCELL_X2 FILLER_83_1338 ();
 FILLCELL_X1 FILLER_83_1343 ();
 FILLCELL_X2 FILLER_83_1351 ();
 FILLCELL_X2 FILLER_83_1370 ();
 FILLCELL_X16 FILLER_83_1382 ();
 FILLCELL_X1 FILLER_83_1398 ();
 FILLCELL_X8 FILLER_83_1429 ();
 FILLCELL_X1 FILLER_83_1437 ();
 FILLCELL_X1 FILLER_83_1443 ();
 FILLCELL_X1 FILLER_83_1449 ();
 FILLCELL_X4 FILLER_83_1471 ();
 FILLCELL_X1 FILLER_83_1475 ();
 FILLCELL_X8 FILLER_83_1485 ();
 FILLCELL_X2 FILLER_83_1493 ();
 FILLCELL_X1 FILLER_83_1495 ();
 FILLCELL_X4 FILLER_83_1518 ();
 FILLCELL_X1 FILLER_83_1531 ();
 FILLCELL_X1 FILLER_83_1536 ();
 FILLCELL_X1 FILLER_83_1541 ();
 FILLCELL_X4 FILLER_83_1570 ();
 FILLCELL_X1 FILLER_83_1574 ();
 FILLCELL_X2 FILLER_83_1594 ();
 FILLCELL_X1 FILLER_83_1608 ();
 FILLCELL_X1 FILLER_83_1619 ();
 FILLCELL_X4 FILLER_83_1627 ();
 FILLCELL_X1 FILLER_83_1631 ();
 FILLCELL_X4 FILLER_83_1635 ();
 FILLCELL_X1 FILLER_83_1639 ();
 FILLCELL_X4 FILLER_83_1644 ();
 FILLCELL_X2 FILLER_83_1648 ();
 FILLCELL_X1 FILLER_83_1650 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X16 FILLER_84_129 ();
 FILLCELL_X4 FILLER_84_145 ();
 FILLCELL_X1 FILLER_84_149 ();
 FILLCELL_X2 FILLER_84_157 ();
 FILLCELL_X2 FILLER_84_179 ();
 FILLCELL_X1 FILLER_84_181 ();
 FILLCELL_X4 FILLER_84_189 ();
 FILLCELL_X1 FILLER_84_193 ();
 FILLCELL_X8 FILLER_84_196 ();
 FILLCELL_X1 FILLER_84_204 ();
 FILLCELL_X2 FILLER_84_222 ();
 FILLCELL_X1 FILLER_84_224 ();
 FILLCELL_X2 FILLER_84_232 ();
 FILLCELL_X1 FILLER_84_240 ();
 FILLCELL_X4 FILLER_84_246 ();
 FILLCELL_X1 FILLER_84_250 ();
 FILLCELL_X4 FILLER_84_255 ();
 FILLCELL_X1 FILLER_84_259 ();
 FILLCELL_X4 FILLER_84_267 ();
 FILLCELL_X1 FILLER_84_285 ();
 FILLCELL_X1 FILLER_84_294 ();
 FILLCELL_X2 FILLER_84_305 ();
 FILLCELL_X2 FILLER_84_323 ();
 FILLCELL_X4 FILLER_84_331 ();
 FILLCELL_X2 FILLER_84_335 ();
 FILLCELL_X4 FILLER_84_344 ();
 FILLCELL_X2 FILLER_84_348 ();
 FILLCELL_X1 FILLER_84_350 ();
 FILLCELL_X1 FILLER_84_358 ();
 FILLCELL_X4 FILLER_84_388 ();
 FILLCELL_X2 FILLER_84_396 ();
 FILLCELL_X2 FILLER_84_403 ();
 FILLCELL_X2 FILLER_84_411 ();
 FILLCELL_X2 FILLER_84_420 ();
 FILLCELL_X1 FILLER_84_422 ();
 FILLCELL_X8 FILLER_84_436 ();
 FILLCELL_X4 FILLER_84_447 ();
 FILLCELL_X1 FILLER_84_465 ();
 FILLCELL_X1 FILLER_84_472 ();
 FILLCELL_X2 FILLER_84_513 ();
 FILLCELL_X2 FILLER_84_524 ();
 FILLCELL_X4 FILLER_84_555 ();
 FILLCELL_X2 FILLER_84_559 ();
 FILLCELL_X2 FILLER_84_565 ();
 FILLCELL_X1 FILLER_84_567 ();
 FILLCELL_X2 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_605 ();
 FILLCELL_X1 FILLER_84_621 ();
 FILLCELL_X2 FILLER_84_654 ();
 FILLCELL_X1 FILLER_84_656 ();
 FILLCELL_X1 FILLER_84_696 ();
 FILLCELL_X2 FILLER_84_700 ();
 FILLCELL_X2 FILLER_84_739 ();
 FILLCELL_X8 FILLER_84_797 ();
 FILLCELL_X2 FILLER_84_805 ();
 FILLCELL_X4 FILLER_84_834 ();
 FILLCELL_X32 FILLER_84_858 ();
 FILLCELL_X4 FILLER_84_890 ();
 FILLCELL_X2 FILLER_84_894 ();
 FILLCELL_X4 FILLER_84_903 ();
 FILLCELL_X2 FILLER_84_907 ();
 FILLCELL_X1 FILLER_84_909 ();
 FILLCELL_X4 FILLER_84_937 ();
 FILLCELL_X2 FILLER_84_941 ();
 FILLCELL_X1 FILLER_84_949 ();
 FILLCELL_X4 FILLER_84_954 ();
 FILLCELL_X1 FILLER_84_958 ();
 FILLCELL_X1 FILLER_84_971 ();
 FILLCELL_X16 FILLER_84_977 ();
 FILLCELL_X8 FILLER_84_993 ();
 FILLCELL_X4 FILLER_84_1001 ();
 FILLCELL_X1 FILLER_84_1005 ();
 FILLCELL_X2 FILLER_84_1011 ();
 FILLCELL_X8 FILLER_84_1018 ();
 FILLCELL_X1 FILLER_84_1035 ();
 FILLCELL_X8 FILLER_84_1056 ();
 FILLCELL_X4 FILLER_84_1064 ();
 FILLCELL_X2 FILLER_84_1068 ();
 FILLCELL_X1 FILLER_84_1070 ();
 FILLCELL_X8 FILLER_84_1093 ();
 FILLCELL_X4 FILLER_84_1101 ();
 FILLCELL_X2 FILLER_84_1105 ();
 FILLCELL_X1 FILLER_84_1107 ();
 FILLCELL_X4 FILLER_84_1117 ();
 FILLCELL_X1 FILLER_84_1121 ();
 FILLCELL_X2 FILLER_84_1157 ();
 FILLCELL_X8 FILLER_84_1162 ();
 FILLCELL_X4 FILLER_84_1199 ();
 FILLCELL_X1 FILLER_84_1203 ();
 FILLCELL_X8 FILLER_84_1210 ();
 FILLCELL_X1 FILLER_84_1218 ();
 FILLCELL_X1 FILLER_84_1225 ();
 FILLCELL_X2 FILLER_84_1236 ();
 FILLCELL_X1 FILLER_84_1297 ();
 FILLCELL_X2 FILLER_84_1312 ();
 FILLCELL_X4 FILLER_84_1321 ();
 FILLCELL_X2 FILLER_84_1328 ();
 FILLCELL_X1 FILLER_84_1330 ();
 FILLCELL_X32 FILLER_84_1338 ();
 FILLCELL_X32 FILLER_84_1370 ();
 FILLCELL_X16 FILLER_84_1402 ();
 FILLCELL_X4 FILLER_84_1418 ();
 FILLCELL_X1 FILLER_84_1422 ();
 FILLCELL_X2 FILLER_84_1453 ();
 FILLCELL_X1 FILLER_84_1485 ();
 FILLCELL_X8 FILLER_84_1491 ();
 FILLCELL_X2 FILLER_84_1499 ();
 FILLCELL_X1 FILLER_84_1511 ();
 FILLCELL_X16 FILLER_84_1524 ();
 FILLCELL_X1 FILLER_84_1540 ();
 FILLCELL_X4 FILLER_84_1551 ();
 FILLCELL_X2 FILLER_84_1555 ();
 FILLCELL_X1 FILLER_84_1557 ();
 FILLCELL_X4 FILLER_84_1562 ();
 FILLCELL_X1 FILLER_84_1574 ();
 FILLCELL_X4 FILLER_84_1579 ();
 FILLCELL_X2 FILLER_84_1583 ();
 FILLCELL_X1 FILLER_84_1585 ();
 FILLCELL_X2 FILLER_84_1590 ();
 FILLCELL_X1 FILLER_84_1596 ();
 FILLCELL_X1 FILLER_84_1601 ();
 FILLCELL_X1 FILLER_84_1605 ();
 FILLCELL_X1 FILLER_84_1610 ();
 FILLCELL_X4 FILLER_84_1614 ();
 FILLCELL_X2 FILLER_84_1627 ();
 FILLCELL_X2 FILLER_84_1636 ();
 FILLCELL_X4 FILLER_84_1644 ();
 FILLCELL_X8 FILLER_85_10 ();
 FILLCELL_X4 FILLER_85_18 ();
 FILLCELL_X2 FILLER_85_22 ();
 FILLCELL_X32 FILLER_85_28 ();
 FILLCELL_X32 FILLER_85_60 ();
 FILLCELL_X32 FILLER_85_92 ();
 FILLCELL_X16 FILLER_85_124 ();
 FILLCELL_X8 FILLER_85_140 ();
 FILLCELL_X4 FILLER_85_148 ();
 FILLCELL_X2 FILLER_85_152 ();
 FILLCELL_X2 FILLER_85_161 ();
 FILLCELL_X16 FILLER_85_170 ();
 FILLCELL_X2 FILLER_85_186 ();
 FILLCELL_X1 FILLER_85_188 ();
 FILLCELL_X8 FILLER_85_194 ();
 FILLCELL_X4 FILLER_85_202 ();
 FILLCELL_X1 FILLER_85_222 ();
 FILLCELL_X2 FILLER_85_240 ();
 FILLCELL_X1 FILLER_85_242 ();
 FILLCELL_X2 FILLER_85_265 ();
 FILLCELL_X16 FILLER_85_290 ();
 FILLCELL_X8 FILLER_85_306 ();
 FILLCELL_X2 FILLER_85_314 ();
 FILLCELL_X1 FILLER_85_360 ();
 FILLCELL_X1 FILLER_85_363 ();
 FILLCELL_X2 FILLER_85_381 ();
 FILLCELL_X1 FILLER_85_406 ();
 FILLCELL_X8 FILLER_85_429 ();
 FILLCELL_X2 FILLER_85_437 ();
 FILLCELL_X1 FILLER_85_461 ();
 FILLCELL_X1 FILLER_85_476 ();
 FILLCELL_X2 FILLER_85_482 ();
 FILLCELL_X4 FILLER_85_490 ();
 FILLCELL_X2 FILLER_85_494 ();
 FILLCELL_X8 FILLER_85_516 ();
 FILLCELL_X1 FILLER_85_524 ();
 FILLCELL_X4 FILLER_85_532 ();
 FILLCELL_X8 FILLER_85_538 ();
 FILLCELL_X2 FILLER_85_546 ();
 FILLCELL_X2 FILLER_85_559 ();
 FILLCELL_X1 FILLER_85_561 ();
 FILLCELL_X4 FILLER_85_569 ();
 FILLCELL_X2 FILLER_85_573 ();
 FILLCELL_X2 FILLER_85_622 ();
 FILLCELL_X8 FILLER_85_637 ();
 FILLCELL_X2 FILLER_85_645 ();
 FILLCELL_X1 FILLER_85_647 ();
 FILLCELL_X1 FILLER_85_682 ();
 FILLCELL_X8 FILLER_85_710 ();
 FILLCELL_X4 FILLER_85_718 ();
 FILLCELL_X2 FILLER_85_722 ();
 FILLCELL_X4 FILLER_85_737 ();
 FILLCELL_X1 FILLER_85_741 ();
 FILLCELL_X1 FILLER_85_783 ();
 FILLCELL_X1 FILLER_85_790 ();
 FILLCELL_X8 FILLER_85_825 ();
 FILLCELL_X2 FILLER_85_833 ();
 FILLCELL_X2 FILLER_85_842 ();
 FILLCELL_X4 FILLER_85_851 ();
 FILLCELL_X2 FILLER_85_862 ();
 FILLCELL_X1 FILLER_85_864 ();
 FILLCELL_X16 FILLER_85_887 ();
 FILLCELL_X4 FILLER_85_903 ();
 FILLCELL_X8 FILLER_85_919 ();
 FILLCELL_X1 FILLER_85_927 ();
 FILLCELL_X32 FILLER_85_936 ();
 FILLCELL_X8 FILLER_85_968 ();
 FILLCELL_X4 FILLER_85_976 ();
 FILLCELL_X2 FILLER_85_980 ();
 FILLCELL_X1 FILLER_85_982 ();
 FILLCELL_X8 FILLER_85_1000 ();
 FILLCELL_X2 FILLER_85_1008 ();
 FILLCELL_X2 FILLER_85_1013 ();
 FILLCELL_X4 FILLER_85_1018 ();
 FILLCELL_X2 FILLER_85_1022 ();
 FILLCELL_X8 FILLER_85_1031 ();
 FILLCELL_X4 FILLER_85_1039 ();
 FILLCELL_X2 FILLER_85_1043 ();
 FILLCELL_X2 FILLER_85_1052 ();
 FILLCELL_X16 FILLER_85_1059 ();
 FILLCELL_X4 FILLER_85_1075 ();
 FILLCELL_X4 FILLER_85_1086 ();
 FILLCELL_X1 FILLER_85_1109 ();
 FILLCELL_X4 FILLER_85_1113 ();
 FILLCELL_X2 FILLER_85_1117 ();
 FILLCELL_X2 FILLER_85_1121 ();
 FILLCELL_X2 FILLER_85_1128 ();
 FILLCELL_X4 FILLER_85_1136 ();
 FILLCELL_X2 FILLER_85_1140 ();
 FILLCELL_X1 FILLER_85_1146 ();
 FILLCELL_X2 FILLER_85_1152 ();
 FILLCELL_X4 FILLER_85_1161 ();
 FILLCELL_X16 FILLER_85_1177 ();
 FILLCELL_X2 FILLER_85_1193 ();
 FILLCELL_X8 FILLER_85_1204 ();
 FILLCELL_X2 FILLER_85_1212 ();
 FILLCELL_X1 FILLER_85_1214 ();
 FILLCELL_X4 FILLER_85_1224 ();
 FILLCELL_X8 FILLER_85_1242 ();
 FILLCELL_X2 FILLER_85_1250 ();
 FILLCELL_X1 FILLER_85_1262 ();
 FILLCELL_X1 FILLER_85_1264 ();
 FILLCELL_X4 FILLER_85_1287 ();
 FILLCELL_X1 FILLER_85_1291 ();
 FILLCELL_X32 FILLER_85_1320 ();
 FILLCELL_X16 FILLER_85_1352 ();
 FILLCELL_X8 FILLER_85_1368 ();
 FILLCELL_X2 FILLER_85_1376 ();
 FILLCELL_X1 FILLER_85_1378 ();
 FILLCELL_X2 FILLER_85_1397 ();
 FILLCELL_X16 FILLER_85_1405 ();
 FILLCELL_X8 FILLER_85_1421 ();
 FILLCELL_X4 FILLER_85_1429 ();
 FILLCELL_X4 FILLER_85_1442 ();
 FILLCELL_X2 FILLER_85_1449 ();
 FILLCELL_X1 FILLER_85_1451 ();
 FILLCELL_X2 FILLER_85_1464 ();
 FILLCELL_X4 FILLER_85_1474 ();
 FILLCELL_X1 FILLER_85_1478 ();
 FILLCELL_X4 FILLER_85_1486 ();
 FILLCELL_X1 FILLER_85_1506 ();
 FILLCELL_X4 FILLER_85_1526 ();
 FILLCELL_X4 FILLER_85_1534 ();
 FILLCELL_X1 FILLER_85_1538 ();
 FILLCELL_X16 FILLER_85_1548 ();
 FILLCELL_X2 FILLER_85_1564 ();
 FILLCELL_X1 FILLER_85_1566 ();
 FILLCELL_X4 FILLER_85_1571 ();
 FILLCELL_X2 FILLER_85_1579 ();
 FILLCELL_X4 FILLER_85_1592 ();
 FILLCELL_X2 FILLER_85_1596 ();
 FILLCELL_X4 FILLER_85_1602 ();
 FILLCELL_X1 FILLER_85_1606 ();
 FILLCELL_X8 FILLER_85_1613 ();
 FILLCELL_X4 FILLER_85_1621 ();
 FILLCELL_X8 FILLER_85_1628 ();
 FILLCELL_X2 FILLER_85_1636 ();
 FILLCELL_X1 FILLER_85_1638 ();
 FILLCELL_X4 FILLER_85_1647 ();
 FILLCELL_X16 FILLER_86_1 ();
 FILLCELL_X4 FILLER_86_17 ();
 FILLCELL_X2 FILLER_86_21 ();
 FILLCELL_X1 FILLER_86_31 ();
 FILLCELL_X32 FILLER_86_36 ();
 FILLCELL_X32 FILLER_86_68 ();
 FILLCELL_X32 FILLER_86_100 ();
 FILLCELL_X16 FILLER_86_132 ();
 FILLCELL_X4 FILLER_86_185 ();
 FILLCELL_X8 FILLER_86_209 ();
 FILLCELL_X4 FILLER_86_217 ();
 FILLCELL_X2 FILLER_86_221 ();
 FILLCELL_X8 FILLER_86_244 ();
 FILLCELL_X1 FILLER_86_260 ();
 FILLCELL_X1 FILLER_86_264 ();
 FILLCELL_X1 FILLER_86_294 ();
 FILLCELL_X2 FILLER_86_315 ();
 FILLCELL_X1 FILLER_86_317 ();
 FILLCELL_X16 FILLER_86_325 ();
 FILLCELL_X8 FILLER_86_341 ();
 FILLCELL_X2 FILLER_86_349 ();
 FILLCELL_X1 FILLER_86_361 ();
 FILLCELL_X2 FILLER_86_368 ();
 FILLCELL_X1 FILLER_86_370 ();
 FILLCELL_X16 FILLER_86_373 ();
 FILLCELL_X4 FILLER_86_389 ();
 FILLCELL_X4 FILLER_86_405 ();
 FILLCELL_X2 FILLER_86_409 ();
 FILLCELL_X1 FILLER_86_411 ();
 FILLCELL_X4 FILLER_86_445 ();
 FILLCELL_X2 FILLER_86_449 ();
 FILLCELL_X2 FILLER_86_457 ();
 FILLCELL_X4 FILLER_86_466 ();
 FILLCELL_X1 FILLER_86_470 ();
 FILLCELL_X8 FILLER_86_494 ();
 FILLCELL_X2 FILLER_86_502 ();
 FILLCELL_X8 FILLER_86_514 ();
 FILLCELL_X1 FILLER_86_522 ();
 FILLCELL_X1 FILLER_86_567 ();
 FILLCELL_X4 FILLER_86_572 ();
 FILLCELL_X1 FILLER_86_576 ();
 FILLCELL_X2 FILLER_86_602 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X2 FILLER_86_625 ();
 FILLCELL_X8 FILLER_86_632 ();
 FILLCELL_X4 FILLER_86_640 ();
 FILLCELL_X1 FILLER_86_644 ();
 FILLCELL_X4 FILLER_86_655 ();
 FILLCELL_X1 FILLER_86_659 ();
 FILLCELL_X2 FILLER_86_669 ();
 FILLCELL_X1 FILLER_86_671 ();
 FILLCELL_X4 FILLER_86_686 ();
 FILLCELL_X2 FILLER_86_694 ();
 FILLCELL_X2 FILLER_86_706 ();
 FILLCELL_X1 FILLER_86_732 ();
 FILLCELL_X2 FILLER_86_740 ();
 FILLCELL_X1 FILLER_86_742 ();
 FILLCELL_X4 FILLER_86_746 ();
 FILLCELL_X1 FILLER_86_750 ();
 FILLCELL_X32 FILLER_86_781 ();
 FILLCELL_X2 FILLER_86_813 ();
 FILLCELL_X1 FILLER_86_815 ();
 FILLCELL_X2 FILLER_86_918 ();
 FILLCELL_X1 FILLER_86_920 ();
 FILLCELL_X4 FILLER_86_927 ();
 FILLCELL_X2 FILLER_86_931 ();
 FILLCELL_X8 FILLER_86_935 ();
 FILLCELL_X4 FILLER_86_943 ();
 FILLCELL_X1 FILLER_86_947 ();
 FILLCELL_X8 FILLER_86_958 ();
 FILLCELL_X4 FILLER_86_966 ();
 FILLCELL_X2 FILLER_86_970 ();
 FILLCELL_X1 FILLER_86_972 ();
 FILLCELL_X2 FILLER_86_1000 ();
 FILLCELL_X1 FILLER_86_1002 ();
 FILLCELL_X4 FILLER_86_1030 ();
 FILLCELL_X1 FILLER_86_1034 ();
 FILLCELL_X8 FILLER_86_1049 ();
 FILLCELL_X2 FILLER_86_1057 ();
 FILLCELL_X2 FILLER_86_1066 ();
 FILLCELL_X1 FILLER_86_1068 ();
 FILLCELL_X2 FILLER_86_1075 ();
 FILLCELL_X4 FILLER_86_1092 ();
 FILLCELL_X2 FILLER_86_1096 ();
 FILLCELL_X1 FILLER_86_1098 ();
 FILLCELL_X4 FILLER_86_1109 ();
 FILLCELL_X1 FILLER_86_1113 ();
 FILLCELL_X1 FILLER_86_1133 ();
 FILLCELL_X2 FILLER_86_1156 ();
 FILLCELL_X1 FILLER_86_1167 ();
 FILLCELL_X4 FILLER_86_1195 ();
 FILLCELL_X1 FILLER_86_1199 ();
 FILLCELL_X2 FILLER_86_1225 ();
 FILLCELL_X2 FILLER_86_1240 ();
 FILLCELL_X1 FILLER_86_1242 ();
 FILLCELL_X4 FILLER_86_1297 ();
 FILLCELL_X1 FILLER_86_1301 ();
 FILLCELL_X8 FILLER_86_1309 ();
 FILLCELL_X4 FILLER_86_1317 ();
 FILLCELL_X2 FILLER_86_1321 ();
 FILLCELL_X8 FILLER_86_1345 ();
 FILLCELL_X2 FILLER_86_1353 ();
 FILLCELL_X1 FILLER_86_1355 ();
 FILLCELL_X1 FILLER_86_1391 ();
 FILLCELL_X2 FILLER_86_1404 ();
 FILLCELL_X1 FILLER_86_1406 ();
 FILLCELL_X16 FILLER_86_1417 ();
 FILLCELL_X8 FILLER_86_1433 ();
 FILLCELL_X4 FILLER_86_1441 ();
 FILLCELL_X8 FILLER_86_1454 ();
 FILLCELL_X2 FILLER_86_1462 ();
 FILLCELL_X1 FILLER_86_1474 ();
 FILLCELL_X2 FILLER_86_1479 ();
 FILLCELL_X2 FILLER_86_1485 ();
 FILLCELL_X2 FILLER_86_1500 ();
 FILLCELL_X1 FILLER_86_1502 ();
 FILLCELL_X4 FILLER_86_1510 ();
 FILLCELL_X1 FILLER_86_1514 ();
 FILLCELL_X4 FILLER_86_1558 ();
 FILLCELL_X1 FILLER_86_1562 ();
 FILLCELL_X16 FILLER_86_1576 ();
 FILLCELL_X8 FILLER_86_1592 ();
 FILLCELL_X2 FILLER_86_1615 ();
 FILLCELL_X16 FILLER_86_1625 ();
 FILLCELL_X8 FILLER_86_1641 ();
 FILLCELL_X2 FILLER_86_1649 ();
 FILLCELL_X8 FILLER_87_1 ();
 FILLCELL_X4 FILLER_87_9 ();
 FILLCELL_X2 FILLER_87_13 ();
 FILLCELL_X32 FILLER_87_19 ();
 FILLCELL_X32 FILLER_87_51 ();
 FILLCELL_X32 FILLER_87_83 ();
 FILLCELL_X32 FILLER_87_115 ();
 FILLCELL_X4 FILLER_87_147 ();
 FILLCELL_X1 FILLER_87_151 ();
 FILLCELL_X1 FILLER_87_159 ();
 FILLCELL_X2 FILLER_87_175 ();
 FILLCELL_X2 FILLER_87_197 ();
 FILLCELL_X1 FILLER_87_232 ();
 FILLCELL_X2 FILLER_87_242 ();
 FILLCELL_X1 FILLER_87_244 ();
 FILLCELL_X2 FILLER_87_248 ();
 FILLCELL_X1 FILLER_87_250 ();
 FILLCELL_X1 FILLER_87_258 ();
 FILLCELL_X4 FILLER_87_265 ();
 FILLCELL_X1 FILLER_87_269 ();
 FILLCELL_X8 FILLER_87_273 ();
 FILLCELL_X4 FILLER_87_281 ();
 FILLCELL_X1 FILLER_87_294 ();
 FILLCELL_X8 FILLER_87_302 ();
 FILLCELL_X2 FILLER_87_341 ();
 FILLCELL_X1 FILLER_87_343 ();
 FILLCELL_X1 FILLER_87_347 ();
 FILLCELL_X2 FILLER_87_355 ();
 FILLCELL_X1 FILLER_87_357 ();
 FILLCELL_X4 FILLER_87_381 ();
 FILLCELL_X1 FILLER_87_385 ();
 FILLCELL_X8 FILLER_87_404 ();
 FILLCELL_X4 FILLER_87_419 ();
 FILLCELL_X2 FILLER_87_423 ();
 FILLCELL_X1 FILLER_87_425 ();
 FILLCELL_X8 FILLER_87_428 ();
 FILLCELL_X4 FILLER_87_436 ();
 FILLCELL_X2 FILLER_87_460 ();
 FILLCELL_X1 FILLER_87_462 ();
 FILLCELL_X1 FILLER_87_483 ();
 FILLCELL_X2 FILLER_87_497 ();
 FILLCELL_X1 FILLER_87_499 ();
 FILLCELL_X8 FILLER_87_525 ();
 FILLCELL_X4 FILLER_87_533 ();
 FILLCELL_X1 FILLER_87_537 ();
 FILLCELL_X4 FILLER_87_542 ();
 FILLCELL_X8 FILLER_87_574 ();
 FILLCELL_X2 FILLER_87_582 ();
 FILLCELL_X4 FILLER_87_596 ();
 FILLCELL_X2 FILLER_87_600 ();
 FILLCELL_X1 FILLER_87_626 ();
 FILLCELL_X1 FILLER_87_631 ();
 FILLCELL_X1 FILLER_87_643 ();
 FILLCELL_X4 FILLER_87_651 ();
 FILLCELL_X1 FILLER_87_655 ();
 FILLCELL_X2 FILLER_87_688 ();
 FILLCELL_X1 FILLER_87_707 ();
 FILLCELL_X2 FILLER_87_725 ();
 FILLCELL_X8 FILLER_87_747 ();
 FILLCELL_X4 FILLER_87_755 ();
 FILLCELL_X2 FILLER_87_759 ();
 FILLCELL_X16 FILLER_87_766 ();
 FILLCELL_X1 FILLER_87_787 ();
 FILLCELL_X16 FILLER_87_817 ();
 FILLCELL_X8 FILLER_87_833 ();
 FILLCELL_X4 FILLER_87_841 ();
 FILLCELL_X1 FILLER_87_845 ();
 FILLCELL_X16 FILLER_87_851 ();
 FILLCELL_X2 FILLER_87_867 ();
 FILLCELL_X4 FILLER_87_883 ();
 FILLCELL_X2 FILLER_87_887 ();
 FILLCELL_X1 FILLER_87_889 ();
 FILLCELL_X4 FILLER_87_897 ();
 FILLCELL_X16 FILLER_87_909 ();
 FILLCELL_X2 FILLER_87_925 ();
 FILLCELL_X1 FILLER_87_927 ();
 FILLCELL_X4 FILLER_87_939 ();
 FILLCELL_X1 FILLER_87_943 ();
 FILLCELL_X1 FILLER_87_968 ();
 FILLCELL_X8 FILLER_87_984 ();
 FILLCELL_X2 FILLER_87_992 ();
 FILLCELL_X8 FILLER_87_998 ();
 FILLCELL_X4 FILLER_87_1006 ();
 FILLCELL_X2 FILLER_87_1010 ();
 FILLCELL_X16 FILLER_87_1019 ();
 FILLCELL_X4 FILLER_87_1035 ();
 FILLCELL_X1 FILLER_87_1039 ();
 FILLCELL_X8 FILLER_87_1050 ();
 FILLCELL_X4 FILLER_87_1058 ();
 FILLCELL_X2 FILLER_87_1062 ();
 FILLCELL_X4 FILLER_87_1084 ();
 FILLCELL_X1 FILLER_87_1088 ();
 FILLCELL_X1 FILLER_87_1108 ();
 FILLCELL_X2 FILLER_87_1112 ();
 FILLCELL_X1 FILLER_87_1124 ();
 FILLCELL_X1 FILLER_87_1130 ();
 FILLCELL_X1 FILLER_87_1133 ();
 FILLCELL_X8 FILLER_87_1139 ();
 FILLCELL_X2 FILLER_87_1147 ();
 FILLCELL_X1 FILLER_87_1149 ();
 FILLCELL_X1 FILLER_87_1164 ();
 FILLCELL_X16 FILLER_87_1172 ();
 FILLCELL_X8 FILLER_87_1188 ();
 FILLCELL_X4 FILLER_87_1196 ();
 FILLCELL_X2 FILLER_87_1200 ();
 FILLCELL_X8 FILLER_87_1231 ();
 FILLCELL_X2 FILLER_87_1239 ();
 FILLCELL_X4 FILLER_87_1250 ();
 FILLCELL_X4 FILLER_87_1264 ();
 FILLCELL_X1 FILLER_87_1268 ();
 FILLCELL_X1 FILLER_87_1273 ();
 FILLCELL_X8 FILLER_87_1277 ();
 FILLCELL_X8 FILLER_87_1306 ();
 FILLCELL_X1 FILLER_87_1314 ();
 FILLCELL_X2 FILLER_87_1318 ();
 FILLCELL_X1 FILLER_87_1324 ();
 FILLCELL_X8 FILLER_87_1334 ();
 FILLCELL_X2 FILLER_87_1342 ();
 FILLCELL_X1 FILLER_87_1344 ();
 FILLCELL_X1 FILLER_87_1365 ();
 FILLCELL_X2 FILLER_87_1376 ();
 FILLCELL_X1 FILLER_87_1384 ();
 FILLCELL_X2 FILLER_87_1395 ();
 FILLCELL_X2 FILLER_87_1403 ();
 FILLCELL_X2 FILLER_87_1415 ();
 FILLCELL_X1 FILLER_87_1417 ();
 FILLCELL_X16 FILLER_87_1428 ();
 FILLCELL_X4 FILLER_87_1444 ();
 FILLCELL_X1 FILLER_87_1448 ();
 FILLCELL_X2 FILLER_87_1452 ();
 FILLCELL_X1 FILLER_87_1454 ();
 FILLCELL_X1 FILLER_87_1475 ();
 FILLCELL_X1 FILLER_87_1489 ();
 FILLCELL_X16 FILLER_87_1498 ();
 FILLCELL_X8 FILLER_87_1514 ();
 FILLCELL_X4 FILLER_87_1522 ();
 FILLCELL_X1 FILLER_87_1552 ();
 FILLCELL_X1 FILLER_87_1558 ();
 FILLCELL_X4 FILLER_87_1576 ();
 FILLCELL_X2 FILLER_87_1580 ();
 FILLCELL_X2 FILLER_87_1605 ();
 FILLCELL_X1 FILLER_87_1611 ();
 FILLCELL_X4 FILLER_87_1616 ();
 FILLCELL_X1 FILLER_87_1620 ();
 FILLCELL_X16 FILLER_87_1632 ();
 FILLCELL_X2 FILLER_87_1648 ();
 FILLCELL_X1 FILLER_87_1650 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X16 FILLER_88_129 ();
 FILLCELL_X8 FILLER_88_145 ();
 FILLCELL_X2 FILLER_88_202 ();
 FILLCELL_X8 FILLER_88_211 ();
 FILLCELL_X2 FILLER_88_247 ();
 FILLCELL_X4 FILLER_88_273 ();
 FILLCELL_X4 FILLER_88_301 ();
 FILLCELL_X1 FILLER_88_305 ();
 FILLCELL_X8 FILLER_88_325 ();
 FILLCELL_X4 FILLER_88_333 ();
 FILLCELL_X2 FILLER_88_365 ();
 FILLCELL_X2 FILLER_88_371 ();
 FILLCELL_X4 FILLER_88_380 ();
 FILLCELL_X1 FILLER_88_384 ();
 FILLCELL_X16 FILLER_88_407 ();
 FILLCELL_X1 FILLER_88_423 ();
 FILLCELL_X4 FILLER_88_431 ();
 FILLCELL_X1 FILLER_88_435 ();
 FILLCELL_X1 FILLER_88_479 ();
 FILLCELL_X1 FILLER_88_537 ();
 FILLCELL_X16 FILLER_88_558 ();
 FILLCELL_X2 FILLER_88_574 ();
 FILLCELL_X1 FILLER_88_576 ();
 FILLCELL_X2 FILLER_88_586 ();
 FILLCELL_X8 FILLER_88_603 ();
 FILLCELL_X4 FILLER_88_611 ();
 FILLCELL_X1 FILLER_88_615 ();
 FILLCELL_X1 FILLER_88_619 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X2 FILLER_88_688 ();
 FILLCELL_X8 FILLER_88_723 ();
 FILLCELL_X1 FILLER_88_731 ();
 FILLCELL_X1 FILLER_88_759 ();
 FILLCELL_X2 FILLER_88_780 ();
 FILLCELL_X2 FILLER_88_802 ();
 FILLCELL_X1 FILLER_88_804 ();
 FILLCELL_X4 FILLER_88_841 ();
 FILLCELL_X2 FILLER_88_867 ();
 FILLCELL_X1 FILLER_88_869 ();
 FILLCELL_X4 FILLER_88_921 ();
 FILLCELL_X2 FILLER_88_925 ();
 FILLCELL_X1 FILLER_88_929 ();
 FILLCELL_X4 FILLER_88_940 ();
 FILLCELL_X2 FILLER_88_944 ();
 FILLCELL_X16 FILLER_88_950 ();
 FILLCELL_X8 FILLER_88_966 ();
 FILLCELL_X4 FILLER_88_974 ();
 FILLCELL_X4 FILLER_88_984 ();
 FILLCELL_X2 FILLER_88_988 ();
 FILLCELL_X1 FILLER_88_990 ();
 FILLCELL_X1 FILLER_88_996 ();
 FILLCELL_X4 FILLER_88_1002 ();
 FILLCELL_X1 FILLER_88_1006 ();
 FILLCELL_X8 FILLER_88_1012 ();
 FILLCELL_X4 FILLER_88_1020 ();
 FILLCELL_X1 FILLER_88_1024 ();
 FILLCELL_X16 FILLER_88_1034 ();
 FILLCELL_X4 FILLER_88_1050 ();
 FILLCELL_X1 FILLER_88_1054 ();
 FILLCELL_X2 FILLER_88_1065 ();
 FILLCELL_X2 FILLER_88_1072 ();
 FILLCELL_X1 FILLER_88_1074 ();
 FILLCELL_X8 FILLER_88_1080 ();
 FILLCELL_X2 FILLER_88_1088 ();
 FILLCELL_X1 FILLER_88_1090 ();
 FILLCELL_X2 FILLER_88_1098 ();
 FILLCELL_X1 FILLER_88_1100 ();
 FILLCELL_X1 FILLER_88_1108 ();
 FILLCELL_X4 FILLER_88_1116 ();
 FILLCELL_X2 FILLER_88_1127 ();
 FILLCELL_X1 FILLER_88_1129 ();
 FILLCELL_X2 FILLER_88_1143 ();
 FILLCELL_X1 FILLER_88_1145 ();
 FILLCELL_X4 FILLER_88_1168 ();
 FILLCELL_X1 FILLER_88_1253 ();
 FILLCELL_X1 FILLER_88_1257 ();
 FILLCELL_X4 FILLER_88_1265 ();
 FILLCELL_X2 FILLER_88_1269 ();
 FILLCELL_X4 FILLER_88_1274 ();
 FILLCELL_X8 FILLER_88_1282 ();
 FILLCELL_X2 FILLER_88_1290 ();
 FILLCELL_X1 FILLER_88_1292 ();
 FILLCELL_X4 FILLER_88_1299 ();
 FILLCELL_X1 FILLER_88_1303 ();
 FILLCELL_X8 FILLER_88_1324 ();
 FILLCELL_X1 FILLER_88_1369 ();
 FILLCELL_X1 FILLER_88_1376 ();
 FILLCELL_X8 FILLER_88_1383 ();
 FILLCELL_X2 FILLER_88_1419 ();
 FILLCELL_X1 FILLER_88_1421 ();
 FILLCELL_X16 FILLER_88_1428 ();
 FILLCELL_X4 FILLER_88_1444 ();
 FILLCELL_X2 FILLER_88_1448 ();
 FILLCELL_X8 FILLER_88_1457 ();
 FILLCELL_X4 FILLER_88_1476 ();
 FILLCELL_X2 FILLER_88_1480 ();
 FILLCELL_X1 FILLER_88_1482 ();
 FILLCELL_X8 FILLER_88_1486 ();
 FILLCELL_X2 FILLER_88_1494 ();
 FILLCELL_X1 FILLER_88_1496 ();
 FILLCELL_X8 FILLER_88_1527 ();
 FILLCELL_X4 FILLER_88_1535 ();
 FILLCELL_X2 FILLER_88_1539 ();
 FILLCELL_X2 FILLER_88_1548 ();
 FILLCELL_X4 FILLER_88_1559 ();
 FILLCELL_X2 FILLER_88_1563 ();
 FILLCELL_X1 FILLER_88_1565 ();
 FILLCELL_X4 FILLER_88_1569 ();
 FILLCELL_X2 FILLER_88_1580 ();
 FILLCELL_X1 FILLER_88_1582 ();
 FILLCELL_X16 FILLER_88_1587 ();
 FILLCELL_X1 FILLER_88_1603 ();
 FILLCELL_X2 FILLER_88_1616 ();
 FILLCELL_X1 FILLER_88_1622 ();
 FILLCELL_X16 FILLER_88_1633 ();
 FILLCELL_X2 FILLER_88_1649 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X16 FILLER_89_161 ();
 FILLCELL_X4 FILLER_89_184 ();
 FILLCELL_X2 FILLER_89_188 ();
 FILLCELL_X1 FILLER_89_190 ();
 FILLCELL_X16 FILLER_89_233 ();
 FILLCELL_X4 FILLER_89_249 ();
 FILLCELL_X2 FILLER_89_253 ();
 FILLCELL_X2 FILLER_89_265 ();
 FILLCELL_X1 FILLER_89_267 ();
 FILLCELL_X4 FILLER_89_281 ();
 FILLCELL_X2 FILLER_89_285 ();
 FILLCELL_X2 FILLER_89_324 ();
 FILLCELL_X16 FILLER_89_333 ();
 FILLCELL_X2 FILLER_89_349 ();
 FILLCELL_X1 FILLER_89_351 ();
 FILLCELL_X4 FILLER_89_405 ();
 FILLCELL_X1 FILLER_89_409 ();
 FILLCELL_X2 FILLER_89_437 ();
 FILLCELL_X8 FILLER_89_461 ();
 FILLCELL_X2 FILLER_89_469 ();
 FILLCELL_X1 FILLER_89_471 ();
 FILLCELL_X4 FILLER_89_501 ();
 FILLCELL_X2 FILLER_89_505 ();
 FILLCELL_X1 FILLER_89_507 ();
 FILLCELL_X4 FILLER_89_515 ();
 FILLCELL_X1 FILLER_89_519 ();
 FILLCELL_X2 FILLER_89_527 ();
 FILLCELL_X1 FILLER_89_529 ();
 FILLCELL_X16 FILLER_89_550 ();
 FILLCELL_X1 FILLER_89_566 ();
 FILLCELL_X8 FILLER_89_574 ();
 FILLCELL_X2 FILLER_89_582 ();
 FILLCELL_X2 FILLER_89_601 ();
 FILLCELL_X2 FILLER_89_610 ();
 FILLCELL_X2 FILLER_89_629 ();
 FILLCELL_X1 FILLER_89_631 ();
 FILLCELL_X1 FILLER_89_636 ();
 FILLCELL_X2 FILLER_89_657 ();
 FILLCELL_X1 FILLER_89_659 ();
 FILLCELL_X16 FILLER_89_680 ();
 FILLCELL_X1 FILLER_89_701 ();
 FILLCELL_X4 FILLER_89_709 ();
 FILLCELL_X2 FILLER_89_713 ();
 FILLCELL_X8 FILLER_89_722 ();
 FILLCELL_X4 FILLER_89_730 ();
 FILLCELL_X2 FILLER_89_734 ();
 FILLCELL_X1 FILLER_89_736 ();
 FILLCELL_X4 FILLER_89_748 ();
 FILLCELL_X2 FILLER_89_759 ();
 FILLCELL_X1 FILLER_89_761 ();
 FILLCELL_X2 FILLER_89_769 ();
 FILLCELL_X2 FILLER_89_798 ();
 FILLCELL_X4 FILLER_89_807 ();
 FILLCELL_X1 FILLER_89_811 ();
 FILLCELL_X4 FILLER_89_819 ();
 FILLCELL_X2 FILLER_89_823 ();
 FILLCELL_X2 FILLER_89_856 ();
 FILLCELL_X1 FILLER_89_858 ();
 FILLCELL_X8 FILLER_89_881 ();
 FILLCELL_X2 FILLER_89_889 ();
 FILLCELL_X1 FILLER_89_891 ();
 FILLCELL_X4 FILLER_89_914 ();
 FILLCELL_X2 FILLER_89_918 ();
 FILLCELL_X4 FILLER_89_924 ();
 FILLCELL_X2 FILLER_89_928 ();
 FILLCELL_X1 FILLER_89_930 ();
 FILLCELL_X8 FILLER_89_945 ();
 FILLCELL_X4 FILLER_89_953 ();
 FILLCELL_X2 FILLER_89_957 ();
 FILLCELL_X8 FILLER_89_966 ();
 FILLCELL_X2 FILLER_89_974 ();
 FILLCELL_X1 FILLER_89_976 ();
 FILLCELL_X16 FILLER_89_981 ();
 FILLCELL_X8 FILLER_89_997 ();
 FILLCELL_X2 FILLER_89_1005 ();
 FILLCELL_X32 FILLER_89_1033 ();
 FILLCELL_X1 FILLER_89_1065 ();
 FILLCELL_X8 FILLER_89_1083 ();
 FILLCELL_X2 FILLER_89_1091 ();
 FILLCELL_X1 FILLER_89_1093 ();
 FILLCELL_X4 FILLER_89_1107 ();
 FILLCELL_X1 FILLER_89_1111 ();
 FILLCELL_X8 FILLER_89_1129 ();
 FILLCELL_X1 FILLER_89_1137 ();
 FILLCELL_X4 FILLER_89_1144 ();
 FILLCELL_X2 FILLER_89_1148 ();
 FILLCELL_X1 FILLER_89_1150 ();
 FILLCELL_X2 FILLER_89_1165 ();
 FILLCELL_X4 FILLER_89_1174 ();
 FILLCELL_X1 FILLER_89_1178 ();
 FILLCELL_X8 FILLER_89_1196 ();
 FILLCELL_X1 FILLER_89_1204 ();
 FILLCELL_X8 FILLER_89_1213 ();
 FILLCELL_X1 FILLER_89_1221 ();
 FILLCELL_X8 FILLER_89_1229 ();
 FILLCELL_X1 FILLER_89_1237 ();
 FILLCELL_X1 FILLER_89_1244 ();
 FILLCELL_X1 FILLER_89_1257 ();
 FILLCELL_X2 FILLER_89_1261 ();
 FILLCELL_X1 FILLER_89_1264 ();
 FILLCELL_X4 FILLER_89_1272 ();
 FILLCELL_X2 FILLER_89_1295 ();
 FILLCELL_X4 FILLER_89_1303 ();
 FILLCELL_X2 FILLER_89_1307 ();
 FILLCELL_X8 FILLER_89_1312 ();
 FILLCELL_X2 FILLER_89_1320 ();
 FILLCELL_X1 FILLER_89_1331 ();
 FILLCELL_X1 FILLER_89_1354 ();
 FILLCELL_X2 FILLER_89_1361 ();
 FILLCELL_X2 FILLER_89_1375 ();
 FILLCELL_X1 FILLER_89_1377 ();
 FILLCELL_X1 FILLER_89_1390 ();
 FILLCELL_X1 FILLER_89_1397 ();
 FILLCELL_X1 FILLER_89_1404 ();
 FILLCELL_X2 FILLER_89_1415 ();
 FILLCELL_X32 FILLER_89_1427 ();
 FILLCELL_X1 FILLER_89_1474 ();
 FILLCELL_X4 FILLER_89_1484 ();
 FILLCELL_X4 FILLER_89_1492 ();
 FILLCELL_X2 FILLER_89_1496 ();
 FILLCELL_X1 FILLER_89_1498 ();
 FILLCELL_X8 FILLER_89_1502 ();
 FILLCELL_X1 FILLER_89_1510 ();
 FILLCELL_X32 FILLER_89_1527 ();
 FILLCELL_X2 FILLER_89_1559 ();
 FILLCELL_X1 FILLER_89_1561 ();
 FILLCELL_X1 FILLER_89_1576 ();
 FILLCELL_X1 FILLER_89_1581 ();
 FILLCELL_X2 FILLER_89_1589 ();
 FILLCELL_X1 FILLER_89_1598 ();
 FILLCELL_X2 FILLER_89_1603 ();
 FILLCELL_X32 FILLER_89_1619 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X16 FILLER_90_129 ();
 FILLCELL_X8 FILLER_90_145 ();
 FILLCELL_X16 FILLER_90_182 ();
 FILLCELL_X4 FILLER_90_225 ();
 FILLCELL_X2 FILLER_90_229 ();
 FILLCELL_X4 FILLER_90_265 ();
 FILLCELL_X2 FILLER_90_269 ();
 FILLCELL_X4 FILLER_90_284 ();
 FILLCELL_X1 FILLER_90_288 ();
 FILLCELL_X2 FILLER_90_294 ();
 FILLCELL_X1 FILLER_90_296 ();
 FILLCELL_X8 FILLER_90_322 ();
 FILLCELL_X4 FILLER_90_330 ();
 FILLCELL_X8 FILLER_90_356 ();
 FILLCELL_X2 FILLER_90_364 ();
 FILLCELL_X1 FILLER_90_366 ();
 FILLCELL_X2 FILLER_90_372 ();
 FILLCELL_X2 FILLER_90_381 ();
 FILLCELL_X4 FILLER_90_390 ();
 FILLCELL_X4 FILLER_90_401 ();
 FILLCELL_X4 FILLER_90_412 ();
 FILLCELL_X16 FILLER_90_421 ();
 FILLCELL_X4 FILLER_90_437 ();
 FILLCELL_X1 FILLER_90_441 ();
 FILLCELL_X8 FILLER_90_449 ();
 FILLCELL_X4 FILLER_90_457 ();
 FILLCELL_X2 FILLER_90_461 ();
 FILLCELL_X1 FILLER_90_506 ();
 FILLCELL_X8 FILLER_90_521 ();
 FILLCELL_X1 FILLER_90_529 ();
 FILLCELL_X2 FILLER_90_551 ();
 FILLCELL_X1 FILLER_90_553 ();
 FILLCELL_X4 FILLER_90_562 ();
 FILLCELL_X1 FILLER_90_566 ();
 FILLCELL_X2 FILLER_90_594 ();
 FILLCELL_X1 FILLER_90_596 ();
 FILLCELL_X16 FILLER_90_614 ();
 FILLCELL_X1 FILLER_90_630 ();
 FILLCELL_X4 FILLER_90_632 ();
 FILLCELL_X1 FILLER_90_636 ();
 FILLCELL_X2 FILLER_90_654 ();
 FILLCELL_X1 FILLER_90_656 ();
 FILLCELL_X4 FILLER_90_664 ();
 FILLCELL_X16 FILLER_90_675 ();
 FILLCELL_X2 FILLER_90_711 ();
 FILLCELL_X2 FILLER_90_733 ();
 FILLCELL_X1 FILLER_90_748 ();
 FILLCELL_X4 FILLER_90_772 ();
 FILLCELL_X2 FILLER_90_783 ();
 FILLCELL_X1 FILLER_90_805 ();
 FILLCELL_X8 FILLER_90_826 ();
 FILLCELL_X2 FILLER_90_834 ();
 FILLCELL_X1 FILLER_90_836 ();
 FILLCELL_X1 FILLER_90_844 ();
 FILLCELL_X4 FILLER_90_852 ();
 FILLCELL_X2 FILLER_90_871 ();
 FILLCELL_X1 FILLER_90_873 ();
 FILLCELL_X4 FILLER_90_903 ();
 FILLCELL_X1 FILLER_90_907 ();
 FILLCELL_X2 FILLER_90_915 ();
 FILLCELL_X1 FILLER_90_917 ();
 FILLCELL_X1 FILLER_90_943 ();
 FILLCELL_X2 FILLER_90_946 ();
 FILLCELL_X1 FILLER_90_955 ();
 FILLCELL_X1 FILLER_90_960 ();
 FILLCELL_X1 FILLER_90_965 ();
 FILLCELL_X4 FILLER_90_969 ();
 FILLCELL_X1 FILLER_90_973 ();
 FILLCELL_X4 FILLER_90_984 ();
 FILLCELL_X2 FILLER_90_988 ();
 FILLCELL_X1 FILLER_90_990 ();
 FILLCELL_X16 FILLER_90_1003 ();
 FILLCELL_X8 FILLER_90_1019 ();
 FILLCELL_X4 FILLER_90_1027 ();
 FILLCELL_X2 FILLER_90_1031 ();
 FILLCELL_X1 FILLER_90_1045 ();
 FILLCELL_X1 FILLER_90_1051 ();
 FILLCELL_X8 FILLER_90_1054 ();
 FILLCELL_X4 FILLER_90_1062 ();
 FILLCELL_X2 FILLER_90_1066 ();
 FILLCELL_X4 FILLER_90_1071 ();
 FILLCELL_X2 FILLER_90_1078 ();
 FILLCELL_X4 FILLER_90_1087 ();
 FILLCELL_X2 FILLER_90_1098 ();
 FILLCELL_X4 FILLER_90_1112 ();
 FILLCELL_X2 FILLER_90_1116 ();
 FILLCELL_X1 FILLER_90_1118 ();
 FILLCELL_X8 FILLER_90_1124 ();
 FILLCELL_X4 FILLER_90_1132 ();
 FILLCELL_X1 FILLER_90_1136 ();
 FILLCELL_X1 FILLER_90_1147 ();
 FILLCELL_X2 FILLER_90_1159 ();
 FILLCELL_X1 FILLER_90_1161 ();
 FILLCELL_X4 FILLER_90_1171 ();
 FILLCELL_X2 FILLER_90_1175 ();
 FILLCELL_X4 FILLER_90_1182 ();
 FILLCELL_X1 FILLER_90_1186 ();
 FILLCELL_X8 FILLER_90_1190 ();
 FILLCELL_X4 FILLER_90_1204 ();
 FILLCELL_X16 FILLER_90_1224 ();
 FILLCELL_X4 FILLER_90_1275 ();
 FILLCELL_X2 FILLER_90_1279 ();
 FILLCELL_X1 FILLER_90_1284 ();
 FILLCELL_X8 FILLER_90_1311 ();
 FILLCELL_X4 FILLER_90_1325 ();
 FILLCELL_X1 FILLER_90_1329 ();
 FILLCELL_X4 FILLER_90_1336 ();
 FILLCELL_X2 FILLER_90_1340 ();
 FILLCELL_X1 FILLER_90_1342 ();
 FILLCELL_X2 FILLER_90_1371 ();
 FILLCELL_X1 FILLER_90_1391 ();
 FILLCELL_X2 FILLER_90_1402 ();
 FILLCELL_X2 FILLER_90_1410 ();
 FILLCELL_X32 FILLER_90_1424 ();
 FILLCELL_X1 FILLER_90_1460 ();
 FILLCELL_X4 FILLER_90_1470 ();
 FILLCELL_X1 FILLER_90_1474 ();
 FILLCELL_X8 FILLER_90_1510 ();
 FILLCELL_X4 FILLER_90_1518 ();
 FILLCELL_X2 FILLER_90_1522 ();
 FILLCELL_X8 FILLER_90_1536 ();
 FILLCELL_X2 FILLER_90_1544 ();
 FILLCELL_X1 FILLER_90_1546 ();
 FILLCELL_X8 FILLER_90_1556 ();
 FILLCELL_X4 FILLER_90_1564 ();
 FILLCELL_X1 FILLER_90_1574 ();
 FILLCELL_X1 FILLER_90_1584 ();
 FILLCELL_X1 FILLER_90_1590 ();
 FILLCELL_X1 FILLER_90_1595 ();
 FILLCELL_X2 FILLER_90_1600 ();
 FILLCELL_X2 FILLER_90_1605 ();
 FILLCELL_X2 FILLER_90_1611 ();
 FILLCELL_X32 FILLER_90_1617 ();
 FILLCELL_X2 FILLER_90_1649 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X16 FILLER_91_129 ();
 FILLCELL_X8 FILLER_91_145 ();
 FILLCELL_X4 FILLER_91_153 ();
 FILLCELL_X2 FILLER_91_157 ();
 FILLCELL_X1 FILLER_91_159 ();
 FILLCELL_X8 FILLER_91_196 ();
 FILLCELL_X32 FILLER_91_238 ();
 FILLCELL_X4 FILLER_91_270 ();
 FILLCELL_X8 FILLER_91_287 ();
 FILLCELL_X1 FILLER_91_295 ();
 FILLCELL_X8 FILLER_91_303 ();
 FILLCELL_X8 FILLER_91_340 ();
 FILLCELL_X2 FILLER_91_348 ();
 FILLCELL_X8 FILLER_91_357 ();
 FILLCELL_X4 FILLER_91_365 ();
 FILLCELL_X2 FILLER_91_369 ();
 FILLCELL_X1 FILLER_91_391 ();
 FILLCELL_X4 FILLER_91_417 ();
 FILLCELL_X8 FILLER_91_443 ();
 FILLCELL_X2 FILLER_91_451 ();
 FILLCELL_X1 FILLER_91_453 ();
 FILLCELL_X4 FILLER_91_461 ();
 FILLCELL_X1 FILLER_91_465 ();
 FILLCELL_X16 FILLER_91_471 ();
 FILLCELL_X4 FILLER_91_487 ();
 FILLCELL_X2 FILLER_91_491 ();
 FILLCELL_X1 FILLER_91_493 ();
 FILLCELL_X2 FILLER_91_516 ();
 FILLCELL_X1 FILLER_91_518 ();
 FILLCELL_X4 FILLER_91_541 ();
 FILLCELL_X1 FILLER_91_545 ();
 FILLCELL_X2 FILLER_91_566 ();
 FILLCELL_X4 FILLER_91_575 ();
 FILLCELL_X1 FILLER_91_579 ();
 FILLCELL_X8 FILLER_91_587 ();
 FILLCELL_X1 FILLER_91_595 ();
 FILLCELL_X1 FILLER_91_623 ();
 FILLCELL_X8 FILLER_91_653 ();
 FILLCELL_X1 FILLER_91_661 ();
 FILLCELL_X4 FILLER_91_682 ();
 FILLCELL_X2 FILLER_91_686 ();
 FILLCELL_X2 FILLER_91_695 ();
 FILLCELL_X1 FILLER_91_697 ();
 FILLCELL_X4 FILLER_91_705 ();
 FILLCELL_X2 FILLER_91_709 ();
 FILLCELL_X1 FILLER_91_738 ();
 FILLCELL_X8 FILLER_91_748 ();
 FILLCELL_X4 FILLER_91_783 ();
 FILLCELL_X2 FILLER_91_787 ();
 FILLCELL_X1 FILLER_91_789 ();
 FILLCELL_X16 FILLER_91_797 ();
 FILLCELL_X8 FILLER_91_813 ();
 FILLCELL_X1 FILLER_91_821 ();
 FILLCELL_X2 FILLER_91_844 ();
 FILLCELL_X1 FILLER_91_846 ();
 FILLCELL_X2 FILLER_91_881 ();
 FILLCELL_X16 FILLER_91_890 ();
 FILLCELL_X4 FILLER_91_928 ();
 FILLCELL_X2 FILLER_91_932 ();
 FILLCELL_X2 FILLER_91_938 ();
 FILLCELL_X1 FILLER_91_940 ();
 FILLCELL_X4 FILLER_91_962 ();
 FILLCELL_X2 FILLER_91_966 ();
 FILLCELL_X8 FILLER_91_978 ();
 FILLCELL_X4 FILLER_91_986 ();
 FILLCELL_X1 FILLER_91_990 ();
 FILLCELL_X8 FILLER_91_999 ();
 FILLCELL_X1 FILLER_91_1007 ();
 FILLCELL_X16 FILLER_91_1019 ();
 FILLCELL_X1 FILLER_91_1035 ();
 FILLCELL_X2 FILLER_91_1041 ();
 FILLCELL_X1 FILLER_91_1043 ();
 FILLCELL_X2 FILLER_91_1049 ();
 FILLCELL_X1 FILLER_91_1051 ();
 FILLCELL_X8 FILLER_91_1057 ();
 FILLCELL_X1 FILLER_91_1065 ();
 FILLCELL_X1 FILLER_91_1072 ();
 FILLCELL_X8 FILLER_91_1078 ();
 FILLCELL_X1 FILLER_91_1086 ();
 FILLCELL_X4 FILLER_91_1094 ();
 FILLCELL_X2 FILLER_91_1098 ();
 FILLCELL_X16 FILLER_91_1146 ();
 FILLCELL_X8 FILLER_91_1162 ();
 FILLCELL_X2 FILLER_91_1170 ();
 FILLCELL_X1 FILLER_91_1193 ();
 FILLCELL_X2 FILLER_91_1247 ();
 FILLCELL_X1 FILLER_91_1249 ();
 FILLCELL_X2 FILLER_91_1257 ();
 FILLCELL_X1 FILLER_91_1259 ();
 FILLCELL_X1 FILLER_91_1296 ();
 FILLCELL_X4 FILLER_91_1301 ();
 FILLCELL_X2 FILLER_91_1305 ();
 FILLCELL_X1 FILLER_91_1307 ();
 FILLCELL_X4 FILLER_91_1311 ();
 FILLCELL_X2 FILLER_91_1315 ();
 FILLCELL_X1 FILLER_91_1317 ();
 FILLCELL_X4 FILLER_91_1324 ();
 FILLCELL_X1 FILLER_91_1340 ();
 FILLCELL_X1 FILLER_91_1347 ();
 FILLCELL_X1 FILLER_91_1354 ();
 FILLCELL_X4 FILLER_91_1361 ();
 FILLCELL_X2 FILLER_91_1377 ();
 FILLCELL_X4 FILLER_91_1385 ();
 FILLCELL_X2 FILLER_91_1389 ();
 FILLCELL_X1 FILLER_91_1391 ();
 FILLCELL_X4 FILLER_91_1398 ();
 FILLCELL_X2 FILLER_91_1402 ();
 FILLCELL_X1 FILLER_91_1404 ();
 FILLCELL_X16 FILLER_91_1425 ();
 FILLCELL_X8 FILLER_91_1441 ();
 FILLCELL_X4 FILLER_91_1449 ();
 FILLCELL_X2 FILLER_91_1453 ();
 FILLCELL_X1 FILLER_91_1459 ();
 FILLCELL_X2 FILLER_91_1491 ();
 FILLCELL_X1 FILLER_91_1493 ();
 FILLCELL_X16 FILLER_91_1522 ();
 FILLCELL_X4 FILLER_91_1538 ();
 FILLCELL_X2 FILLER_91_1542 ();
 FILLCELL_X4 FILLER_91_1548 ();
 FILLCELL_X1 FILLER_91_1552 ();
 FILLCELL_X8 FILLER_91_1557 ();
 FILLCELL_X4 FILLER_91_1565 ();
 FILLCELL_X1 FILLER_91_1569 ();
 FILLCELL_X2 FILLER_91_1574 ();
 FILLCELL_X2 FILLER_91_1594 ();
 FILLCELL_X1 FILLER_91_1600 ();
 FILLCELL_X2 FILLER_91_1605 ();
 FILLCELL_X2 FILLER_91_1613 ();
 FILLCELL_X1 FILLER_91_1619 ();
 FILLCELL_X8 FILLER_91_1640 ();
 FILLCELL_X2 FILLER_91_1648 ();
 FILLCELL_X1 FILLER_91_1650 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X16 FILLER_92_129 ();
 FILLCELL_X8 FILLER_92_145 ();
 FILLCELL_X2 FILLER_92_153 ();
 FILLCELL_X1 FILLER_92_155 ();
 FILLCELL_X32 FILLER_92_176 ();
 FILLCELL_X16 FILLER_92_208 ();
 FILLCELL_X2 FILLER_92_224 ();
 FILLCELL_X2 FILLER_92_231 ();
 FILLCELL_X4 FILLER_92_237 ();
 FILLCELL_X2 FILLER_92_241 ();
 FILLCELL_X1 FILLER_92_243 ();
 FILLCELL_X4 FILLER_92_249 ();
 FILLCELL_X1 FILLER_92_253 ();
 FILLCELL_X2 FILLER_92_268 ();
 FILLCELL_X2 FILLER_92_297 ();
 FILLCELL_X4 FILLER_92_304 ();
 FILLCELL_X1 FILLER_92_308 ();
 FILLCELL_X8 FILLER_92_316 ();
 FILLCELL_X1 FILLER_92_324 ();
 FILLCELL_X4 FILLER_92_332 ();
 FILLCELL_X2 FILLER_92_336 ();
 FILLCELL_X1 FILLER_92_338 ();
 FILLCELL_X2 FILLER_92_368 ();
 FILLCELL_X8 FILLER_92_377 ();
 FILLCELL_X2 FILLER_92_385 ();
 FILLCELL_X16 FILLER_92_392 ();
 FILLCELL_X4 FILLER_92_408 ();
 FILLCELL_X4 FILLER_92_419 ();
 FILLCELL_X1 FILLER_92_423 ();
 FILLCELL_X4 FILLER_92_431 ();
 FILLCELL_X1 FILLER_92_435 ();
 FILLCELL_X2 FILLER_92_523 ();
 FILLCELL_X16 FILLER_92_532 ();
 FILLCELL_X2 FILLER_92_602 ();
 FILLCELL_X2 FILLER_92_639 ();
 FILLCELL_X1 FILLER_92_641 ();
 FILLCELL_X1 FILLER_92_662 ();
 FILLCELL_X2 FILLER_92_698 ();
 FILLCELL_X1 FILLER_92_700 ();
 FILLCELL_X2 FILLER_92_723 ();
 FILLCELL_X1 FILLER_92_725 ();
 FILLCELL_X4 FILLER_92_734 ();
 FILLCELL_X1 FILLER_92_738 ();
 FILLCELL_X2 FILLER_92_766 ();
 FILLCELL_X1 FILLER_92_768 ();
 FILLCELL_X16 FILLER_92_772 ();
 FILLCELL_X4 FILLER_92_788 ();
 FILLCELL_X8 FILLER_92_821 ();
 FILLCELL_X4 FILLER_92_829 ();
 FILLCELL_X2 FILLER_92_833 ();
 FILLCELL_X1 FILLER_92_835 ();
 FILLCELL_X2 FILLER_92_850 ();
 FILLCELL_X1 FILLER_92_852 ();
 FILLCELL_X4 FILLER_92_880 ();
 FILLCELL_X2 FILLER_92_884 ();
 FILLCELL_X4 FILLER_92_908 ();
 FILLCELL_X2 FILLER_92_912 ();
 FILLCELL_X1 FILLER_92_914 ();
 FILLCELL_X8 FILLER_92_948 ();
 FILLCELL_X4 FILLER_92_956 ();
 FILLCELL_X2 FILLER_92_960 ();
 FILLCELL_X1 FILLER_92_962 ();
 FILLCELL_X16 FILLER_92_968 ();
 FILLCELL_X2 FILLER_92_984 ();
 FILLCELL_X8 FILLER_92_991 ();
 FILLCELL_X2 FILLER_92_1014 ();
 FILLCELL_X1 FILLER_92_1016 ();
 FILLCELL_X2 FILLER_92_1022 ();
 FILLCELL_X4 FILLER_92_1027 ();
 FILLCELL_X4 FILLER_92_1038 ();
 FILLCELL_X2 FILLER_92_1042 ();
 FILLCELL_X1 FILLER_92_1044 ();
 FILLCELL_X16 FILLER_92_1054 ();
 FILLCELL_X2 FILLER_92_1070 ();
 FILLCELL_X1 FILLER_92_1103 ();
 FILLCELL_X1 FILLER_92_1106 ();
 FILLCELL_X1 FILLER_92_1116 ();
 FILLCELL_X4 FILLER_92_1148 ();
 FILLCELL_X2 FILLER_92_1152 ();
 FILLCELL_X1 FILLER_92_1154 ();
 FILLCELL_X8 FILLER_92_1161 ();
 FILLCELL_X1 FILLER_92_1169 ();
 FILLCELL_X8 FILLER_92_1176 ();
 FILLCELL_X4 FILLER_92_1184 ();
 FILLCELL_X1 FILLER_92_1194 ();
 FILLCELL_X2 FILLER_92_1216 ();
 FILLCELL_X8 FILLER_92_1228 ();
 FILLCELL_X4 FILLER_92_1236 ();
 FILLCELL_X1 FILLER_92_1250 ();
 FILLCELL_X4 FILLER_92_1258 ();
 FILLCELL_X2 FILLER_92_1262 ();
 FILLCELL_X2 FILLER_92_1270 ();
 FILLCELL_X1 FILLER_92_1272 ();
 FILLCELL_X1 FILLER_92_1286 ();
 FILLCELL_X1 FILLER_92_1352 ();
 FILLCELL_X1 FILLER_92_1359 ();
 FILLCELL_X8 FILLER_92_1366 ();
 FILLCELL_X1 FILLER_92_1402 ();
 FILLCELL_X2 FILLER_92_1409 ();
 FILLCELL_X2 FILLER_92_1417 ();
 FILLCELL_X32 FILLER_92_1429 ();
 FILLCELL_X8 FILLER_92_1461 ();
 FILLCELL_X2 FILLER_92_1472 ();
 FILLCELL_X1 FILLER_92_1474 ();
 FILLCELL_X16 FILLER_92_1487 ();
 FILLCELL_X4 FILLER_92_1503 ();
 FILLCELL_X4 FILLER_92_1522 ();
 FILLCELL_X4 FILLER_92_1535 ();
 FILLCELL_X2 FILLER_92_1539 ();
 FILLCELL_X4 FILLER_92_1587 ();
 FILLCELL_X2 FILLER_92_1591 ();
 FILLCELL_X1 FILLER_92_1604 ();
 FILLCELL_X4 FILLER_92_1608 ();
 FILLCELL_X1 FILLER_92_1612 ();
 FILLCELL_X16 FILLER_92_1630 ();
 FILLCELL_X4 FILLER_92_1646 ();
 FILLCELL_X1 FILLER_92_1650 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X16 FILLER_93_161 ();
 FILLCELL_X8 FILLER_93_177 ();
 FILLCELL_X2 FILLER_93_185 ();
 FILLCELL_X1 FILLER_93_187 ();
 FILLCELL_X8 FILLER_93_197 ();
 FILLCELL_X1 FILLER_93_205 ();
 FILLCELL_X2 FILLER_93_235 ();
 FILLCELL_X1 FILLER_93_237 ();
 FILLCELL_X16 FILLER_93_282 ();
 FILLCELL_X2 FILLER_93_298 ();
 FILLCELL_X1 FILLER_93_300 ();
 FILLCELL_X4 FILLER_93_323 ();
 FILLCELL_X8 FILLER_93_349 ();
 FILLCELL_X8 FILLER_93_379 ();
 FILLCELL_X4 FILLER_93_387 ();
 FILLCELL_X4 FILLER_93_442 ();
 FILLCELL_X1 FILLER_93_446 ();
 FILLCELL_X1 FILLER_93_467 ();
 FILLCELL_X1 FILLER_93_494 ();
 FILLCELL_X2 FILLER_93_499 ();
 FILLCELL_X4 FILLER_93_510 ();
 FILLCELL_X4 FILLER_93_543 ();
 FILLCELL_X2 FILLER_93_547 ();
 FILLCELL_X8 FILLER_93_569 ();
 FILLCELL_X2 FILLER_93_577 ();
 FILLCELL_X2 FILLER_93_606 ();
 FILLCELL_X1 FILLER_93_608 ();
 FILLCELL_X2 FILLER_93_614 ();
 FILLCELL_X1 FILLER_93_616 ();
 FILLCELL_X8 FILLER_93_651 ();
 FILLCELL_X4 FILLER_93_659 ();
 FILLCELL_X8 FILLER_93_673 ();
 FILLCELL_X2 FILLER_93_681 ();
 FILLCELL_X1 FILLER_93_710 ();
 FILLCELL_X4 FILLER_93_745 ();
 FILLCELL_X2 FILLER_93_749 ();
 FILLCELL_X16 FILLER_93_758 ();
 FILLCELL_X4 FILLER_93_774 ();
 FILLCELL_X4 FILLER_93_791 ();
 FILLCELL_X16 FILLER_93_817 ();
 FILLCELL_X8 FILLER_93_833 ();
 FILLCELL_X1 FILLER_93_841 ();
 FILLCELL_X4 FILLER_93_871 ();
 FILLCELL_X1 FILLER_93_875 ();
 FILLCELL_X2 FILLER_93_912 ();
 FILLCELL_X1 FILLER_93_914 ();
 FILLCELL_X8 FILLER_93_922 ();
 FILLCELL_X2 FILLER_93_934 ();
 FILLCELL_X1 FILLER_93_942 ();
 FILLCELL_X2 FILLER_93_964 ();
 FILLCELL_X4 FILLER_93_971 ();
 FILLCELL_X2 FILLER_93_975 ();
 FILLCELL_X1 FILLER_93_977 ();
 FILLCELL_X2 FILLER_93_992 ();
 FILLCELL_X2 FILLER_93_1006 ();
 FILLCELL_X1 FILLER_93_1008 ();
 FILLCELL_X4 FILLER_93_1011 ();
 FILLCELL_X2 FILLER_93_1015 ();
 FILLCELL_X8 FILLER_93_1026 ();
 FILLCELL_X1 FILLER_93_1034 ();
 FILLCELL_X2 FILLER_93_1047 ();
 FILLCELL_X1 FILLER_93_1049 ();
 FILLCELL_X16 FILLER_93_1059 ();
 FILLCELL_X4 FILLER_93_1075 ();
 FILLCELL_X1 FILLER_93_1079 ();
 FILLCELL_X4 FILLER_93_1087 ();
 FILLCELL_X2 FILLER_93_1091 ();
 FILLCELL_X1 FILLER_93_1093 ();
 FILLCELL_X8 FILLER_93_1104 ();
 FILLCELL_X1 FILLER_93_1112 ();
 FILLCELL_X4 FILLER_93_1118 ();
 FILLCELL_X1 FILLER_93_1136 ();
 FILLCELL_X2 FILLER_93_1144 ();
 FILLCELL_X8 FILLER_93_1168 ();
 FILLCELL_X2 FILLER_93_1176 ();
 FILLCELL_X8 FILLER_93_1200 ();
 FILLCELL_X2 FILLER_93_1208 ();
 FILLCELL_X4 FILLER_93_1230 ();
 FILLCELL_X1 FILLER_93_1234 ();
 FILLCELL_X2 FILLER_93_1260 ();
 FILLCELL_X1 FILLER_93_1262 ();
 FILLCELL_X4 FILLER_93_1264 ();
 FILLCELL_X2 FILLER_93_1268 ();
 FILLCELL_X2 FILLER_93_1281 ();
 FILLCELL_X1 FILLER_93_1283 ();
 FILLCELL_X16 FILLER_93_1288 ();
 FILLCELL_X8 FILLER_93_1304 ();
 FILLCELL_X4 FILLER_93_1312 ();
 FILLCELL_X2 FILLER_93_1322 ();
 FILLCELL_X2 FILLER_93_1336 ();
 FILLCELL_X1 FILLER_93_1338 ();
 FILLCELL_X1 FILLER_93_1349 ();
 FILLCELL_X2 FILLER_93_1356 ();
 FILLCELL_X1 FILLER_93_1358 ();
 FILLCELL_X1 FILLER_93_1371 ();
 FILLCELL_X4 FILLER_93_1378 ();
 FILLCELL_X8 FILLER_93_1392 ();
 FILLCELL_X4 FILLER_93_1400 ();
 FILLCELL_X1 FILLER_93_1416 ();
 FILLCELL_X32 FILLER_93_1437 ();
 FILLCELL_X8 FILLER_93_1484 ();
 FILLCELL_X1 FILLER_93_1510 ();
 FILLCELL_X2 FILLER_93_1523 ();
 FILLCELL_X1 FILLER_93_1525 ();
 FILLCELL_X4 FILLER_93_1538 ();
 FILLCELL_X2 FILLER_93_1560 ();
 FILLCELL_X1 FILLER_93_1562 ();
 FILLCELL_X16 FILLER_93_1570 ();
 FILLCELL_X4 FILLER_93_1586 ();
 FILLCELL_X1 FILLER_93_1590 ();
 FILLCELL_X2 FILLER_93_1599 ();
 FILLCELL_X4 FILLER_93_1605 ();
 FILLCELL_X2 FILLER_93_1609 ();
 FILLCELL_X2 FILLER_93_1618 ();
 FILLCELL_X1 FILLER_93_1620 ();
 FILLCELL_X16 FILLER_93_1629 ();
 FILLCELL_X4 FILLER_93_1645 ();
 FILLCELL_X2 FILLER_93_1649 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X4 FILLER_94_221 ();
 FILLCELL_X2 FILLER_94_225 ();
 FILLCELL_X1 FILLER_94_256 ();
 FILLCELL_X8 FILLER_94_280 ();
 FILLCELL_X2 FILLER_94_288 ();
 FILLCELL_X2 FILLER_94_300 ();
 FILLCELL_X8 FILLER_94_309 ();
 FILLCELL_X2 FILLER_94_317 ();
 FILLCELL_X1 FILLER_94_319 ();
 FILLCELL_X2 FILLER_94_452 ();
 FILLCELL_X1 FILLER_94_454 ();
 FILLCELL_X1 FILLER_94_480 ();
 FILLCELL_X16 FILLER_94_506 ();
 FILLCELL_X8 FILLER_94_529 ();
 FILLCELL_X4 FILLER_94_537 ();
 FILLCELL_X4 FILLER_94_563 ();
 FILLCELL_X1 FILLER_94_567 ();
 FILLCELL_X8 FILLER_94_584 ();
 FILLCELL_X2 FILLER_94_592 ();
 FILLCELL_X1 FILLER_94_601 ();
 FILLCELL_X16 FILLER_94_632 ();
 FILLCELL_X4 FILLER_94_648 ();
 FILLCELL_X2 FILLER_94_652 ();
 FILLCELL_X1 FILLER_94_654 ();
 FILLCELL_X2 FILLER_94_682 ();
 FILLCELL_X4 FILLER_94_706 ();
 FILLCELL_X2 FILLER_94_710 ();
 FILLCELL_X8 FILLER_94_734 ();
 FILLCELL_X4 FILLER_94_742 ();
 FILLCELL_X2 FILLER_94_746 ();
 FILLCELL_X1 FILLER_94_748 ();
 FILLCELL_X2 FILLER_94_758 ();
 FILLCELL_X1 FILLER_94_760 ();
 FILLCELL_X2 FILLER_94_790 ();
 FILLCELL_X2 FILLER_94_798 ();
 FILLCELL_X1 FILLER_94_800 ();
 FILLCELL_X2 FILLER_94_808 ();
 FILLCELL_X1 FILLER_94_810 ();
 FILLCELL_X2 FILLER_94_833 ();
 FILLCELL_X8 FILLER_94_842 ();
 FILLCELL_X4 FILLER_94_850 ();
 FILLCELL_X2 FILLER_94_854 ();
 FILLCELL_X16 FILLER_94_885 ();
 FILLCELL_X2 FILLER_94_901 ();
 FILLCELL_X4 FILLER_94_925 ();
 FILLCELL_X2 FILLER_94_929 ();
 FILLCELL_X16 FILLER_94_935 ();
 FILLCELL_X8 FILLER_94_951 ();
 FILLCELL_X4 FILLER_94_959 ();
 FILLCELL_X2 FILLER_94_963 ();
 FILLCELL_X1 FILLER_94_965 ();
 FILLCELL_X4 FILLER_94_979 ();
 FILLCELL_X2 FILLER_94_983 ();
 FILLCELL_X2 FILLER_94_989 ();
 FILLCELL_X16 FILLER_94_1004 ();
 FILLCELL_X1 FILLER_94_1020 ();
 FILLCELL_X8 FILLER_94_1025 ();
 FILLCELL_X2 FILLER_94_1033 ();
 FILLCELL_X2 FILLER_94_1049 ();
 FILLCELL_X1 FILLER_94_1051 ();
 FILLCELL_X16 FILLER_94_1070 ();
 FILLCELL_X8 FILLER_94_1086 ();
 FILLCELL_X4 FILLER_94_1094 ();
 FILLCELL_X8 FILLER_94_1108 ();
 FILLCELL_X1 FILLER_94_1116 ();
 FILLCELL_X2 FILLER_94_1127 ();
 FILLCELL_X4 FILLER_94_1140 ();
 FILLCELL_X1 FILLER_94_1144 ();
 FILLCELL_X4 FILLER_94_1151 ();
 FILLCELL_X2 FILLER_94_1155 ();
 FILLCELL_X8 FILLER_94_1163 ();
 FILLCELL_X2 FILLER_94_1171 ();
 FILLCELL_X1 FILLER_94_1173 ();
 FILLCELL_X16 FILLER_94_1180 ();
 FILLCELL_X8 FILLER_94_1196 ();
 FILLCELL_X2 FILLER_94_1204 ();
 FILLCELL_X1 FILLER_94_1206 ();
 FILLCELL_X4 FILLER_94_1232 ();
 FILLCELL_X2 FILLER_94_1236 ();
 FILLCELL_X1 FILLER_94_1247 ();
 FILLCELL_X1 FILLER_94_1252 ();
 FILLCELL_X2 FILLER_94_1331 ();
 FILLCELL_X1 FILLER_94_1333 ();
 FILLCELL_X4 FILLER_94_1350 ();
 FILLCELL_X1 FILLER_94_1364 ();
 FILLCELL_X4 FILLER_94_1377 ();
 FILLCELL_X2 FILLER_94_1381 ();
 FILLCELL_X1 FILLER_94_1383 ();
 FILLCELL_X4 FILLER_94_1394 ();
 FILLCELL_X32 FILLER_94_1418 ();
 FILLCELL_X8 FILLER_94_1450 ();
 FILLCELL_X1 FILLER_94_1477 ();
 FILLCELL_X1 FILLER_94_1482 ();
 FILLCELL_X4 FILLER_94_1485 ();
 FILLCELL_X1 FILLER_94_1530 ();
 FILLCELL_X2 FILLER_94_1540 ();
 FILLCELL_X1 FILLER_94_1547 ();
 FILLCELL_X2 FILLER_94_1553 ();
 FILLCELL_X1 FILLER_94_1562 ();
 FILLCELL_X8 FILLER_94_1566 ();
 FILLCELL_X1 FILLER_94_1574 ();
 FILLCELL_X2 FILLER_94_1595 ();
 FILLCELL_X32 FILLER_94_1609 ();
 FILLCELL_X8 FILLER_94_1641 ();
 FILLCELL_X2 FILLER_94_1649 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X8 FILLER_95_161 ();
 FILLCELL_X4 FILLER_95_169 ();
 FILLCELL_X1 FILLER_95_173 ();
 FILLCELL_X2 FILLER_95_182 ();
 FILLCELL_X2 FILLER_95_211 ();
 FILLCELL_X1 FILLER_95_213 ();
 FILLCELL_X8 FILLER_95_217 ();
 FILLCELL_X2 FILLER_95_225 ();
 FILLCELL_X1 FILLER_95_227 ();
 FILLCELL_X4 FILLER_95_252 ();
 FILLCELL_X2 FILLER_95_256 ();
 FILLCELL_X8 FILLER_95_265 ();
 FILLCELL_X1 FILLER_95_273 ();
 FILLCELL_X2 FILLER_95_312 ();
 FILLCELL_X8 FILLER_95_321 ();
 FILLCELL_X4 FILLER_95_329 ();
 FILLCELL_X2 FILLER_95_333 ();
 FILLCELL_X1 FILLER_95_345 ();
 FILLCELL_X4 FILLER_95_366 ();
 FILLCELL_X1 FILLER_95_370 ();
 FILLCELL_X2 FILLER_95_386 ();
 FILLCELL_X1 FILLER_95_388 ();
 FILLCELL_X2 FILLER_95_396 ();
 FILLCELL_X16 FILLER_95_407 ();
 FILLCELL_X2 FILLER_95_439 ();
 FILLCELL_X4 FILLER_95_444 ();
 FILLCELL_X2 FILLER_95_448 ();
 FILLCELL_X1 FILLER_95_456 ();
 FILLCELL_X8 FILLER_95_466 ();
 FILLCELL_X1 FILLER_95_474 ();
 FILLCELL_X16 FILLER_95_484 ();
 FILLCELL_X1 FILLER_95_500 ();
 FILLCELL_X1 FILLER_95_557 ();
 FILLCELL_X8 FILLER_95_588 ();
 FILLCELL_X2 FILLER_95_603 ();
 FILLCELL_X1 FILLER_95_605 ();
 FILLCELL_X8 FILLER_95_611 ();
 FILLCELL_X2 FILLER_95_619 ();
 FILLCELL_X1 FILLER_95_621 ();
 FILLCELL_X2 FILLER_95_629 ();
 FILLCELL_X1 FILLER_95_631 ();
 FILLCELL_X4 FILLER_95_679 ();
 FILLCELL_X2 FILLER_95_683 ();
 FILLCELL_X1 FILLER_95_685 ();
 FILLCELL_X2 FILLER_95_693 ();
 FILLCELL_X1 FILLER_95_695 ();
 FILLCELL_X8 FILLER_95_703 ();
 FILLCELL_X4 FILLER_95_711 ();
 FILLCELL_X2 FILLER_95_715 ();
 FILLCELL_X1 FILLER_95_717 ();
 FILLCELL_X1 FILLER_95_723 ();
 FILLCELL_X16 FILLER_95_763 ();
 FILLCELL_X2 FILLER_95_779 ();
 FILLCELL_X8 FILLER_95_877 ();
 FILLCELL_X4 FILLER_95_885 ();
 FILLCELL_X16 FILLER_95_901 ();
 FILLCELL_X8 FILLER_95_917 ();
 FILLCELL_X4 FILLER_95_934 ();
 FILLCELL_X4 FILLER_95_953 ();
 FILLCELL_X2 FILLER_95_957 ();
 FILLCELL_X8 FILLER_95_970 ();
 FILLCELL_X4 FILLER_95_978 ();
 FILLCELL_X1 FILLER_95_982 ();
 FILLCELL_X2 FILLER_95_985 ();
 FILLCELL_X4 FILLER_95_992 ();
 FILLCELL_X16 FILLER_95_1006 ();
 FILLCELL_X4 FILLER_95_1022 ();
 FILLCELL_X2 FILLER_95_1032 ();
 FILLCELL_X16 FILLER_95_1038 ();
 FILLCELL_X8 FILLER_95_1058 ();
 FILLCELL_X1 FILLER_95_1066 ();
 FILLCELL_X4 FILLER_95_1069 ();
 FILLCELL_X2 FILLER_95_1073 ();
 FILLCELL_X1 FILLER_95_1075 ();
 FILLCELL_X1 FILLER_95_1086 ();
 FILLCELL_X2 FILLER_95_1089 ();
 FILLCELL_X1 FILLER_95_1096 ();
 FILLCELL_X1 FILLER_95_1107 ();
 FILLCELL_X2 FILLER_95_1112 ();
 FILLCELL_X2 FILLER_95_1129 ();
 FILLCELL_X2 FILLER_95_1193 ();
 FILLCELL_X32 FILLER_95_1227 ();
 FILLCELL_X4 FILLER_95_1259 ();
 FILLCELL_X16 FILLER_95_1282 ();
 FILLCELL_X1 FILLER_95_1298 ();
 FILLCELL_X2 FILLER_95_1303 ();
 FILLCELL_X1 FILLER_95_1305 ();
 FILLCELL_X1 FILLER_95_1310 ();
 FILLCELL_X8 FILLER_95_1314 ();
 FILLCELL_X1 FILLER_95_1322 ();
 FILLCELL_X1 FILLER_95_1365 ();
 FILLCELL_X4 FILLER_95_1372 ();
 FILLCELL_X2 FILLER_95_1376 ();
 FILLCELL_X1 FILLER_95_1378 ();
 FILLCELL_X1 FILLER_95_1401 ();
 FILLCELL_X8 FILLER_95_1414 ();
 FILLCELL_X4 FILLER_95_1422 ();
 FILLCELL_X1 FILLER_95_1426 ();
 FILLCELL_X4 FILLER_95_1433 ();
 FILLCELL_X8 FILLER_95_1447 ();
 FILLCELL_X4 FILLER_95_1462 ();
 FILLCELL_X2 FILLER_95_1475 ();
 FILLCELL_X1 FILLER_95_1477 ();
 FILLCELL_X1 FILLER_95_1482 ();
 FILLCELL_X1 FILLER_95_1488 ();
 FILLCELL_X1 FILLER_95_1493 ();
 FILLCELL_X1 FILLER_95_1497 ();
 FILLCELL_X2 FILLER_95_1503 ();
 FILLCELL_X1 FILLER_95_1562 ();
 FILLCELL_X2 FILLER_95_1567 ();
 FILLCELL_X1 FILLER_95_1569 ();
 FILLCELL_X4 FILLER_95_1575 ();
 FILLCELL_X2 FILLER_95_1579 ();
 FILLCELL_X1 FILLER_95_1581 ();
 FILLCELL_X1 FILLER_95_1585 ();
 FILLCELL_X2 FILLER_95_1597 ();
 FILLCELL_X2 FILLER_95_1602 ();
 FILLCELL_X32 FILLER_95_1607 ();
 FILLCELL_X8 FILLER_95_1639 ();
 FILLCELL_X4 FILLER_95_1647 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X8 FILLER_96_129 ();
 FILLCELL_X4 FILLER_96_137 ();
 FILLCELL_X2 FILLER_96_141 ();
 FILLCELL_X1 FILLER_96_202 ();
 FILLCELL_X2 FILLER_96_211 ();
 FILLCELL_X1 FILLER_96_213 ();
 FILLCELL_X4 FILLER_96_223 ();
 FILLCELL_X1 FILLER_96_227 ();
 FILLCELL_X2 FILLER_96_247 ();
 FILLCELL_X4 FILLER_96_255 ();
 FILLCELL_X2 FILLER_96_259 ();
 FILLCELL_X4 FILLER_96_283 ();
 FILLCELL_X1 FILLER_96_291 ();
 FILLCELL_X8 FILLER_96_327 ();
 FILLCELL_X4 FILLER_96_335 ();
 FILLCELL_X1 FILLER_96_342 ();
 FILLCELL_X8 FILLER_96_356 ();
 FILLCELL_X2 FILLER_96_364 ();
 FILLCELL_X1 FILLER_96_366 ();
 FILLCELL_X4 FILLER_96_380 ();
 FILLCELL_X2 FILLER_96_384 ();
 FILLCELL_X1 FILLER_96_435 ();
 FILLCELL_X2 FILLER_96_453 ();
 FILLCELL_X4 FILLER_96_465 ();
 FILLCELL_X1 FILLER_96_469 ();
 FILLCELL_X2 FILLER_96_493 ();
 FILLCELL_X1 FILLER_96_508 ();
 FILLCELL_X8 FILLER_96_531 ();
 FILLCELL_X2 FILLER_96_539 ();
 FILLCELL_X8 FILLER_96_546 ();
 FILLCELL_X4 FILLER_96_554 ();
 FILLCELL_X2 FILLER_96_558 ();
 FILLCELL_X1 FILLER_96_560 ();
 FILLCELL_X4 FILLER_96_590 ();
 FILLCELL_X8 FILLER_96_616 ();
 FILLCELL_X4 FILLER_96_624 ();
 FILLCELL_X2 FILLER_96_628 ();
 FILLCELL_X1 FILLER_96_630 ();
 FILLCELL_X2 FILLER_96_632 ();
 FILLCELL_X1 FILLER_96_634 ();
 FILLCELL_X1 FILLER_96_647 ();
 FILLCELL_X16 FILLER_96_727 ();
 FILLCELL_X2 FILLER_96_761 ();
 FILLCELL_X1 FILLER_96_763 ();
 FILLCELL_X2 FILLER_96_791 ();
 FILLCELL_X2 FILLER_96_815 ();
 FILLCELL_X2 FILLER_96_829 ();
 FILLCELL_X32 FILLER_96_838 ();
 FILLCELL_X1 FILLER_96_870 ();
 FILLCELL_X1 FILLER_96_896 ();
 FILLCELL_X8 FILLER_96_919 ();
 FILLCELL_X1 FILLER_96_947 ();
 FILLCELL_X2 FILLER_96_952 ();
 FILLCELL_X1 FILLER_96_963 ();
 FILLCELL_X2 FILLER_96_968 ();
 FILLCELL_X1 FILLER_96_970 ();
 FILLCELL_X2 FILLER_96_976 ();
 FILLCELL_X1 FILLER_96_978 ();
 FILLCELL_X8 FILLER_96_994 ();
 FILLCELL_X4 FILLER_96_1002 ();
 FILLCELL_X1 FILLER_96_1017 ();
 FILLCELL_X16 FILLER_96_1052 ();
 FILLCELL_X8 FILLER_96_1068 ();
 FILLCELL_X2 FILLER_96_1081 ();
 FILLCELL_X1 FILLER_96_1083 ();
 FILLCELL_X2 FILLER_96_1110 ();
 FILLCELL_X2 FILLER_96_1122 ();
 FILLCELL_X8 FILLER_96_1130 ();
 FILLCELL_X2 FILLER_96_1153 ();
 FILLCELL_X2 FILLER_96_1158 ();
 FILLCELL_X2 FILLER_96_1170 ();
 FILLCELL_X8 FILLER_96_1177 ();
 FILLCELL_X4 FILLER_96_1185 ();
 FILLCELL_X2 FILLER_96_1189 ();
 FILLCELL_X1 FILLER_96_1199 ();
 FILLCELL_X8 FILLER_96_1255 ();
 FILLCELL_X2 FILLER_96_1263 ();
 FILLCELL_X1 FILLER_96_1268 ();
 FILLCELL_X4 FILLER_96_1278 ();
 FILLCELL_X2 FILLER_96_1282 ();
 FILLCELL_X1 FILLER_96_1297 ();
 FILLCELL_X2 FILLER_96_1308 ();
 FILLCELL_X4 FILLER_96_1338 ();
 FILLCELL_X8 FILLER_96_1362 ();
 FILLCELL_X1 FILLER_96_1370 ();
 FILLCELL_X4 FILLER_96_1420 ();
 FILLCELL_X2 FILLER_96_1424 ();
 FILLCELL_X1 FILLER_96_1426 ();
 FILLCELL_X16 FILLER_96_1437 ();
 FILLCELL_X4 FILLER_96_1453 ();
 FILLCELL_X1 FILLER_96_1457 ();
 FILLCELL_X4 FILLER_96_1469 ();
 FILLCELL_X1 FILLER_96_1473 ();
 FILLCELL_X1 FILLER_96_1485 ();
 FILLCELL_X1 FILLER_96_1490 ();
 FILLCELL_X1 FILLER_96_1498 ();
 FILLCELL_X1 FILLER_96_1504 ();
 FILLCELL_X8 FILLER_96_1514 ();
 FILLCELL_X2 FILLER_96_1522 ();
 FILLCELL_X8 FILLER_96_1553 ();
 FILLCELL_X2 FILLER_96_1561 ();
 FILLCELL_X4 FILLER_96_1567 ();
 FILLCELL_X1 FILLER_96_1571 ();
 FILLCELL_X2 FILLER_96_1580 ();
 FILLCELL_X1 FILLER_96_1582 ();
 FILLCELL_X2 FILLER_96_1595 ();
 FILLCELL_X2 FILLER_96_1601 ();
 FILLCELL_X1 FILLER_96_1603 ();
 FILLCELL_X4 FILLER_96_1612 ();
 FILLCELL_X2 FILLER_96_1616 ();
 FILLCELL_X1 FILLER_96_1618 ();
 FILLCELL_X16 FILLER_96_1625 ();
 FILLCELL_X8 FILLER_96_1641 ();
 FILLCELL_X2 FILLER_96_1649 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X16 FILLER_97_97 ();
 FILLCELL_X8 FILLER_97_113 ();
 FILLCELL_X2 FILLER_97_121 ();
 FILLCELL_X4 FILLER_97_143 ();
 FILLCELL_X2 FILLER_97_147 ();
 FILLCELL_X1 FILLER_97_149 ();
 FILLCELL_X4 FILLER_97_190 ();
 FILLCELL_X1 FILLER_97_194 ();
 FILLCELL_X16 FILLER_97_217 ();
 FILLCELL_X1 FILLER_97_233 ();
 FILLCELL_X16 FILLER_97_256 ();
 FILLCELL_X4 FILLER_97_272 ();
 FILLCELL_X1 FILLER_97_276 ();
 FILLCELL_X4 FILLER_97_290 ();
 FILLCELL_X1 FILLER_97_294 ();
 FILLCELL_X4 FILLER_97_308 ();
 FILLCELL_X2 FILLER_97_409 ();
 FILLCELL_X8 FILLER_97_414 ();
 FILLCELL_X4 FILLER_97_422 ();
 FILLCELL_X4 FILLER_97_450 ();
 FILLCELL_X1 FILLER_97_454 ();
 FILLCELL_X1 FILLER_97_486 ();
 FILLCELL_X8 FILLER_97_514 ();
 FILLCELL_X4 FILLER_97_522 ();
 FILLCELL_X8 FILLER_97_533 ();
 FILLCELL_X4 FILLER_97_541 ();
 FILLCELL_X1 FILLER_97_545 ();
 FILLCELL_X8 FILLER_97_553 ();
 FILLCELL_X1 FILLER_97_561 ();
 FILLCELL_X1 FILLER_97_582 ();
 FILLCELL_X16 FILLER_97_585 ();
 FILLCELL_X4 FILLER_97_601 ();
 FILLCELL_X2 FILLER_97_605 ();
 FILLCELL_X2 FILLER_97_614 ();
 FILLCELL_X1 FILLER_97_616 ();
 FILLCELL_X2 FILLER_97_646 ();
 FILLCELL_X1 FILLER_97_648 ();
 FILLCELL_X8 FILLER_97_676 ();
 FILLCELL_X4 FILLER_97_684 ();
 FILLCELL_X2 FILLER_97_688 ();
 FILLCELL_X1 FILLER_97_690 ();
 FILLCELL_X4 FILLER_97_710 ();
 FILLCELL_X1 FILLER_97_721 ();
 FILLCELL_X1 FILLER_97_744 ();
 FILLCELL_X32 FILLER_97_765 ();
 FILLCELL_X16 FILLER_97_797 ();
 FILLCELL_X2 FILLER_97_813 ();
 FILLCELL_X1 FILLER_97_815 ();
 FILLCELL_X16 FILLER_97_838 ();
 FILLCELL_X2 FILLER_97_854 ();
 FILLCELL_X8 FILLER_97_914 ();
 FILLCELL_X4 FILLER_97_922 ();
 FILLCELL_X2 FILLER_97_926 ();
 FILLCELL_X1 FILLER_97_928 ();
 FILLCELL_X4 FILLER_97_932 ();
 FILLCELL_X1 FILLER_97_952 ();
 FILLCELL_X1 FILLER_97_964 ();
 FILLCELL_X1 FILLER_97_972 ();
 FILLCELL_X2 FILLER_97_977 ();
 FILLCELL_X8 FILLER_97_987 ();
 FILLCELL_X4 FILLER_97_995 ();
 FILLCELL_X8 FILLER_97_1008 ();
 FILLCELL_X1 FILLER_97_1016 ();
 FILLCELL_X2 FILLER_97_1026 ();
 FILLCELL_X2 FILLER_97_1030 ();
 FILLCELL_X1 FILLER_97_1032 ();
 FILLCELL_X1 FILLER_97_1037 ();
 FILLCELL_X1 FILLER_97_1041 ();
 FILLCELL_X1 FILLER_97_1047 ();
 FILLCELL_X4 FILLER_97_1053 ();
 FILLCELL_X2 FILLER_97_1057 ();
 FILLCELL_X1 FILLER_97_1059 ();
 FILLCELL_X2 FILLER_97_1065 ();
 FILLCELL_X1 FILLER_97_1067 ();
 FILLCELL_X1 FILLER_97_1071 ();
 FILLCELL_X4 FILLER_97_1082 ();
 FILLCELL_X1 FILLER_97_1086 ();
 FILLCELL_X1 FILLER_97_1128 ();
 FILLCELL_X2 FILLER_97_1139 ();
 FILLCELL_X4 FILLER_97_1147 ();
 FILLCELL_X2 FILLER_97_1181 ();
 FILLCELL_X1 FILLER_97_1183 ();
 FILLCELL_X1 FILLER_97_1196 ();
 FILLCELL_X1 FILLER_97_1200 ();
 FILLCELL_X8 FILLER_97_1208 ();
 FILLCELL_X1 FILLER_97_1216 ();
 FILLCELL_X4 FILLER_97_1221 ();
 FILLCELL_X4 FILLER_97_1230 ();
 FILLCELL_X4 FILLER_97_1244 ();
 FILLCELL_X2 FILLER_97_1258 ();
 FILLCELL_X8 FILLER_97_1286 ();
 FILLCELL_X1 FILLER_97_1294 ();
 FILLCELL_X4 FILLER_97_1301 ();
 FILLCELL_X4 FILLER_97_1333 ();
 FILLCELL_X1 FILLER_97_1359 ();
 FILLCELL_X4 FILLER_97_1370 ();
 FILLCELL_X4 FILLER_97_1390 ();
 FILLCELL_X1 FILLER_97_1394 ();
 FILLCELL_X4 FILLER_97_1401 ();
 FILLCELL_X1 FILLER_97_1405 ();
 FILLCELL_X2 FILLER_97_1412 ();
 FILLCELL_X1 FILLER_97_1414 ();
 FILLCELL_X32 FILLER_97_1425 ();
 FILLCELL_X4 FILLER_97_1457 ();
 FILLCELL_X2 FILLER_97_1474 ();
 FILLCELL_X4 FILLER_97_1487 ();
 FILLCELL_X1 FILLER_97_1497 ();
 FILLCELL_X8 FILLER_97_1509 ();
 FILLCELL_X2 FILLER_97_1525 ();
 FILLCELL_X2 FILLER_97_1530 ();
 FILLCELL_X1 FILLER_97_1541 ();
 FILLCELL_X16 FILLER_97_1551 ();
 FILLCELL_X2 FILLER_97_1567 ();
 FILLCELL_X1 FILLER_97_1588 ();
 FILLCELL_X2 FILLER_97_1592 ();
 FILLCELL_X16 FILLER_97_1606 ();
 FILLCELL_X8 FILLER_97_1622 ();
 FILLCELL_X4 FILLER_97_1630 ();
 FILLCELL_X8 FILLER_97_1637 ();
 FILLCELL_X2 FILLER_97_1648 ();
 FILLCELL_X1 FILLER_97_1650 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X16 FILLER_98_33 ();
 FILLCELL_X8 FILLER_98_49 ();
 FILLCELL_X2 FILLER_98_57 ();
 FILLCELL_X16 FILLER_98_66 ();
 FILLCELL_X4 FILLER_98_82 ();
 FILLCELL_X2 FILLER_98_86 ();
 FILLCELL_X1 FILLER_98_88 ();
 FILLCELL_X4 FILLER_98_96 ();
 FILLCELL_X2 FILLER_98_100 ();
 FILLCELL_X1 FILLER_98_102 ();
 FILLCELL_X8 FILLER_98_130 ();
 FILLCELL_X1 FILLER_98_150 ();
 FILLCELL_X4 FILLER_98_195 ();
 FILLCELL_X2 FILLER_98_199 ();
 FILLCELL_X1 FILLER_98_201 ();
 FILLCELL_X2 FILLER_98_249 ();
 FILLCELL_X8 FILLER_98_253 ();
 FILLCELL_X4 FILLER_98_261 ();
 FILLCELL_X2 FILLER_98_265 ();
 FILLCELL_X8 FILLER_98_272 ();
 FILLCELL_X2 FILLER_98_280 ();
 FILLCELL_X8 FILLER_98_289 ();
 FILLCELL_X4 FILLER_98_297 ();
 FILLCELL_X1 FILLER_98_301 ();
 FILLCELL_X4 FILLER_98_325 ();
 FILLCELL_X2 FILLER_98_329 ();
 FILLCELL_X1 FILLER_98_331 ();
 FILLCELL_X1 FILLER_98_352 ();
 FILLCELL_X4 FILLER_98_383 ();
 FILLCELL_X2 FILLER_98_387 ();
 FILLCELL_X8 FILLER_98_396 ();
 FILLCELL_X2 FILLER_98_404 ();
 FILLCELL_X2 FILLER_98_413 ();
 FILLCELL_X1 FILLER_98_415 ();
 FILLCELL_X4 FILLER_98_491 ();
 FILLCELL_X2 FILLER_98_495 ();
 FILLCELL_X1 FILLER_98_497 ();
 FILLCELL_X2 FILLER_98_622 ();
 FILLCELL_X8 FILLER_98_632 ();
 FILLCELL_X8 FILLER_98_676 ();
 FILLCELL_X1 FILLER_98_684 ();
 FILLCELL_X4 FILLER_98_732 ();
 FILLCELL_X1 FILLER_98_736 ();
 FILLCELL_X1 FILLER_98_740 ();
 FILLCELL_X1 FILLER_98_748 ();
 FILLCELL_X1 FILLER_98_756 ();
 FILLCELL_X1 FILLER_98_779 ();
 FILLCELL_X2 FILLER_98_783 ();
 FILLCELL_X2 FILLER_98_788 ();
 FILLCELL_X2 FILLER_98_810 ();
 FILLCELL_X2 FILLER_98_841 ();
 FILLCELL_X1 FILLER_98_843 ();
 FILLCELL_X1 FILLER_98_864 ();
 FILLCELL_X4 FILLER_98_879 ();
 FILLCELL_X2 FILLER_98_883 ();
 FILLCELL_X4 FILLER_98_892 ();
 FILLCELL_X16 FILLER_98_925 ();
 FILLCELL_X8 FILLER_98_941 ();
 FILLCELL_X1 FILLER_98_954 ();
 FILLCELL_X8 FILLER_98_962 ();
 FILLCELL_X2 FILLER_98_970 ();
 FILLCELL_X1 FILLER_98_972 ();
 FILLCELL_X4 FILLER_98_983 ();
 FILLCELL_X2 FILLER_98_987 ();
 FILLCELL_X1 FILLER_98_989 ();
 FILLCELL_X8 FILLER_98_997 ();
 FILLCELL_X4 FILLER_98_1005 ();
 FILLCELL_X2 FILLER_98_1009 ();
 FILLCELL_X16 FILLER_98_1026 ();
 FILLCELL_X4 FILLER_98_1042 ();
 FILLCELL_X2 FILLER_98_1056 ();
 FILLCELL_X16 FILLER_98_1076 ();
 FILLCELL_X4 FILLER_98_1092 ();
 FILLCELL_X2 FILLER_98_1096 ();
 FILLCELL_X4 FILLER_98_1101 ();
 FILLCELL_X1 FILLER_98_1105 ();
 FILLCELL_X2 FILLER_98_1119 ();
 FILLCELL_X1 FILLER_98_1127 ();
 FILLCELL_X2 FILLER_98_1139 ();
 FILLCELL_X1 FILLER_98_1141 ();
 FILLCELL_X8 FILLER_98_1146 ();
 FILLCELL_X1 FILLER_98_1156 ();
 FILLCELL_X16 FILLER_98_1163 ();
 FILLCELL_X1 FILLER_98_1179 ();
 FILLCELL_X2 FILLER_98_1186 ();
 FILLCELL_X1 FILLER_98_1188 ();
 FILLCELL_X4 FILLER_98_1216 ();
 FILLCELL_X2 FILLER_98_1220 ();
 FILLCELL_X1 FILLER_98_1222 ();
 FILLCELL_X8 FILLER_98_1239 ();
 FILLCELL_X2 FILLER_98_1256 ();
 FILLCELL_X1 FILLER_98_1258 ();
 FILLCELL_X1 FILLER_98_1266 ();
 FILLCELL_X2 FILLER_98_1277 ();
 FILLCELL_X1 FILLER_98_1279 ();
 FILLCELL_X8 FILLER_98_1284 ();
 FILLCELL_X2 FILLER_98_1292 ();
 FILLCELL_X1 FILLER_98_1311 ();
 FILLCELL_X4 FILLER_98_1315 ();
 FILLCELL_X1 FILLER_98_1319 ();
 FILLCELL_X4 FILLER_98_1335 ();
 FILLCELL_X4 FILLER_98_1355 ();
 FILLCELL_X1 FILLER_98_1359 ();
 FILLCELL_X4 FILLER_98_1372 ();
 FILLCELL_X16 FILLER_98_1434 ();
 FILLCELL_X8 FILLER_98_1450 ();
 FILLCELL_X4 FILLER_98_1458 ();
 FILLCELL_X2 FILLER_98_1462 ();
 FILLCELL_X1 FILLER_98_1464 ();
 FILLCELL_X4 FILLER_98_1487 ();
 FILLCELL_X2 FILLER_98_1491 ();
 FILLCELL_X2 FILLER_98_1496 ();
 FILLCELL_X2 FILLER_98_1512 ();
 FILLCELL_X2 FILLER_98_1545 ();
 FILLCELL_X4 FILLER_98_1554 ();
 FILLCELL_X2 FILLER_98_1558 ();
 FILLCELL_X1 FILLER_98_1560 ();
 FILLCELL_X1 FILLER_98_1567 ();
 FILLCELL_X2 FILLER_98_1575 ();
 FILLCELL_X1 FILLER_98_1582 ();
 FILLCELL_X2 FILLER_98_1594 ();
 FILLCELL_X2 FILLER_98_1600 ();
 FILLCELL_X2 FILLER_98_1605 ();
 FILLCELL_X1 FILLER_98_1607 ();
 FILLCELL_X8 FILLER_98_1616 ();
 FILLCELL_X16 FILLER_98_1633 ();
 FILLCELL_X2 FILLER_98_1649 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X16 FILLER_99_33 ();
 FILLCELL_X2 FILLER_99_49 ();
 FILLCELL_X1 FILLER_99_51 ();
 FILLCELL_X4 FILLER_99_72 ();
 FILLCELL_X4 FILLER_99_96 ();
 FILLCELL_X1 FILLER_99_100 ();
 FILLCELL_X8 FILLER_99_121 ();
 FILLCELL_X1 FILLER_99_129 ();
 FILLCELL_X1 FILLER_99_171 ();
 FILLCELL_X8 FILLER_99_202 ();
 FILLCELL_X1 FILLER_99_210 ();
 FILLCELL_X4 FILLER_99_231 ();
 FILLCELL_X2 FILLER_99_235 ();
 FILLCELL_X1 FILLER_99_244 ();
 FILLCELL_X1 FILLER_99_285 ();
 FILLCELL_X8 FILLER_99_313 ();
 FILLCELL_X4 FILLER_99_321 ();
 FILLCELL_X2 FILLER_99_325 ();
 FILLCELL_X1 FILLER_99_327 ();
 FILLCELL_X8 FILLER_99_331 ();
 FILLCELL_X2 FILLER_99_339 ();
 FILLCELL_X1 FILLER_99_341 ();
 FILLCELL_X2 FILLER_99_352 ();
 FILLCELL_X4 FILLER_99_368 ();
 FILLCELL_X4 FILLER_99_418 ();
 FILLCELL_X2 FILLER_99_422 ();
 FILLCELL_X1 FILLER_99_424 ();
 FILLCELL_X4 FILLER_99_507 ();
 FILLCELL_X2 FILLER_99_521 ();
 FILLCELL_X2 FILLER_99_543 ();
 FILLCELL_X1 FILLER_99_545 ();
 FILLCELL_X4 FILLER_99_551 ();
 FILLCELL_X2 FILLER_99_555 ();
 FILLCELL_X8 FILLER_99_573 ();
 FILLCELL_X2 FILLER_99_581 ();
 FILLCELL_X8 FILLER_99_590 ();
 FILLCELL_X2 FILLER_99_598 ();
 FILLCELL_X1 FILLER_99_600 ();
 FILLCELL_X8 FILLER_99_657 ();
 FILLCELL_X4 FILLER_99_665 ();
 FILLCELL_X2 FILLER_99_669 ();
 FILLCELL_X1 FILLER_99_671 ();
 FILLCELL_X4 FILLER_99_702 ();
 FILLCELL_X2 FILLER_99_706 ();
 FILLCELL_X8 FILLER_99_744 ();
 FILLCELL_X4 FILLER_99_752 ();
 FILLCELL_X2 FILLER_99_762 ();
 FILLCELL_X32 FILLER_99_798 ();
 FILLCELL_X4 FILLER_99_830 ();
 FILLCELL_X1 FILLER_99_834 ();
 FILLCELL_X2 FILLER_99_865 ();
 FILLCELL_X8 FILLER_99_874 ();
 FILLCELL_X4 FILLER_99_882 ();
 FILLCELL_X4 FILLER_99_913 ();
 FILLCELL_X2 FILLER_99_917 ();
 FILLCELL_X16 FILLER_99_954 ();
 FILLCELL_X4 FILLER_99_970 ();
 FILLCELL_X2 FILLER_99_974 ();
 FILLCELL_X4 FILLER_99_986 ();
 FILLCELL_X4 FILLER_99_1001 ();
 FILLCELL_X2 FILLER_99_1005 ();
 FILLCELL_X16 FILLER_99_1025 ();
 FILLCELL_X8 FILLER_99_1041 ();
 FILLCELL_X1 FILLER_99_1049 ();
 FILLCELL_X1 FILLER_99_1060 ();
 FILLCELL_X16 FILLER_99_1066 ();
 FILLCELL_X4 FILLER_99_1082 ();
 FILLCELL_X2 FILLER_99_1086 ();
 FILLCELL_X1 FILLER_99_1088 ();
 FILLCELL_X16 FILLER_99_1118 ();
 FILLCELL_X8 FILLER_99_1134 ();
 FILLCELL_X16 FILLER_99_1151 ();
 FILLCELL_X1 FILLER_99_1167 ();
 FILLCELL_X2 FILLER_99_1190 ();
 FILLCELL_X1 FILLER_99_1192 ();
 FILLCELL_X1 FILLER_99_1209 ();
 FILLCELL_X1 FILLER_99_1232 ();
 FILLCELL_X8 FILLER_99_1255 ();
 FILLCELL_X4 FILLER_99_1293 ();
 FILLCELL_X2 FILLER_99_1302 ();
 FILLCELL_X16 FILLER_99_1310 ();
 FILLCELL_X2 FILLER_99_1326 ();
 FILLCELL_X4 FILLER_99_1334 ();
 FILLCELL_X2 FILLER_99_1338 ();
 FILLCELL_X1 FILLER_99_1346 ();
 FILLCELL_X1 FILLER_99_1353 ();
 FILLCELL_X16 FILLER_99_1366 ();
 FILLCELL_X2 FILLER_99_1382 ();
 FILLCELL_X1 FILLER_99_1384 ();
 FILLCELL_X2 FILLER_99_1403 ();
 FILLCELL_X1 FILLER_99_1405 ();
 FILLCELL_X16 FILLER_99_1435 ();
 FILLCELL_X4 FILLER_99_1451 ();
 FILLCELL_X2 FILLER_99_1455 ();
 FILLCELL_X4 FILLER_99_1461 ();
 FILLCELL_X2 FILLER_99_1465 ();
 FILLCELL_X1 FILLER_99_1467 ();
 FILLCELL_X16 FILLER_99_1505 ();
 FILLCELL_X1 FILLER_99_1521 ();
 FILLCELL_X1 FILLER_99_1546 ();
 FILLCELL_X16 FILLER_99_1551 ();
 FILLCELL_X1 FILLER_99_1578 ();
 FILLCELL_X1 FILLER_99_1584 ();
 FILLCELL_X2 FILLER_99_1589 ();
 FILLCELL_X2 FILLER_99_1595 ();
 FILLCELL_X4 FILLER_99_1602 ();
 FILLCELL_X1 FILLER_99_1606 ();
 FILLCELL_X1 FILLER_99_1613 ();
 FILLCELL_X4 FILLER_99_1621 ();
 FILLCELL_X1 FILLER_99_1625 ();
 FILLCELL_X16 FILLER_99_1629 ();
 FILLCELL_X4 FILLER_99_1645 ();
 FILLCELL_X2 FILLER_99_1649 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X8 FILLER_100_33 ();
 FILLCELL_X4 FILLER_100_41 ();
 FILLCELL_X2 FILLER_100_45 ();
 FILLCELL_X1 FILLER_100_47 ();
 FILLCELL_X16 FILLER_100_53 ();
 FILLCELL_X16 FILLER_100_89 ();
 FILLCELL_X2 FILLER_100_112 ();
 FILLCELL_X1 FILLER_100_121 ();
 FILLCELL_X4 FILLER_100_156 ();
 FILLCELL_X2 FILLER_100_160 ();
 FILLCELL_X16 FILLER_100_169 ();
 FILLCELL_X1 FILLER_100_185 ();
 FILLCELL_X2 FILLER_100_193 ();
 FILLCELL_X1 FILLER_100_195 ();
 FILLCELL_X4 FILLER_100_216 ();
 FILLCELL_X2 FILLER_100_220 ();
 FILLCELL_X1 FILLER_100_229 ();
 FILLCELL_X2 FILLER_100_241 ();
 FILLCELL_X1 FILLER_100_243 ();
 FILLCELL_X2 FILLER_100_264 ();
 FILLCELL_X4 FILLER_100_286 ();
 FILLCELL_X32 FILLER_100_294 ();
 FILLCELL_X16 FILLER_100_326 ();
 FILLCELL_X2 FILLER_100_358 ();
 FILLCELL_X4 FILLER_100_367 ();
 FILLCELL_X2 FILLER_100_371 ();
 FILLCELL_X8 FILLER_100_383 ();
 FILLCELL_X1 FILLER_100_391 ();
 FILLCELL_X4 FILLER_100_405 ();
 FILLCELL_X8 FILLER_100_416 ();
 FILLCELL_X1 FILLER_100_424 ();
 FILLCELL_X8 FILLER_100_469 ();
 FILLCELL_X2 FILLER_100_477 ();
 FILLCELL_X4 FILLER_100_484 ();
 FILLCELL_X2 FILLER_100_488 ();
 FILLCELL_X1 FILLER_100_490 ();
 FILLCELL_X2 FILLER_100_527 ();
 FILLCELL_X1 FILLER_100_529 ();
 FILLCELL_X2 FILLER_100_550 ();
 FILLCELL_X1 FILLER_100_552 ();
 FILLCELL_X1 FILLER_100_578 ();
 FILLCELL_X4 FILLER_100_601 ();
 FILLCELL_X2 FILLER_100_605 ();
 FILLCELL_X1 FILLER_100_616 ();
 FILLCELL_X4 FILLER_100_627 ();
 FILLCELL_X2 FILLER_100_632 ();
 FILLCELL_X1 FILLER_100_634 ();
 FILLCELL_X16 FILLER_100_638 ();
 FILLCELL_X4 FILLER_100_654 ();
 FILLCELL_X2 FILLER_100_658 ();
 FILLCELL_X4 FILLER_100_711 ();
 FILLCELL_X8 FILLER_100_724 ();
 FILLCELL_X4 FILLER_100_732 ();
 FILLCELL_X2 FILLER_100_736 ();
 FILLCELL_X1 FILLER_100_738 ();
 FILLCELL_X8 FILLER_100_766 ();
 FILLCELL_X2 FILLER_100_774 ();
 FILLCELL_X16 FILLER_100_816 ();
 FILLCELL_X2 FILLER_100_846 ();
 FILLCELL_X1 FILLER_100_848 ();
 FILLCELL_X8 FILLER_100_900 ();
 FILLCELL_X1 FILLER_100_908 ();
 FILLCELL_X4 FILLER_100_936 ();
 FILLCELL_X2 FILLER_100_940 ();
 FILLCELL_X1 FILLER_100_942 ();
 FILLCELL_X4 FILLER_100_949 ();
 FILLCELL_X2 FILLER_100_953 ();
 FILLCELL_X1 FILLER_100_955 ();
 FILLCELL_X8 FILLER_100_959 ();
 FILLCELL_X4 FILLER_100_967 ();
 FILLCELL_X1 FILLER_100_971 ();
 FILLCELL_X1 FILLER_100_978 ();
 FILLCELL_X16 FILLER_100_982 ();
 FILLCELL_X8 FILLER_100_1013 ();
 FILLCELL_X1 FILLER_100_1021 ();
 FILLCELL_X2 FILLER_100_1034 ();
 FILLCELL_X4 FILLER_100_1039 ();
 FILLCELL_X2 FILLER_100_1048 ();
 FILLCELL_X4 FILLER_100_1055 ();
 FILLCELL_X4 FILLER_100_1062 ();
 FILLCELL_X2 FILLER_100_1066 ();
 FILLCELL_X16 FILLER_100_1080 ();
 FILLCELL_X8 FILLER_100_1096 ();
 FILLCELL_X1 FILLER_100_1104 ();
 FILLCELL_X4 FILLER_100_1114 ();
 FILLCELL_X2 FILLER_100_1118 ();
 FILLCELL_X2 FILLER_100_1147 ();
 FILLCELL_X1 FILLER_100_1159 ();
 FILLCELL_X2 FILLER_100_1165 ();
 FILLCELL_X1 FILLER_100_1186 ();
 FILLCELL_X8 FILLER_100_1192 ();
 FILLCELL_X2 FILLER_100_1200 ();
 FILLCELL_X1 FILLER_100_1218 ();
 FILLCELL_X4 FILLER_100_1229 ();
 FILLCELL_X2 FILLER_100_1233 ();
 FILLCELL_X1 FILLER_100_1247 ();
 FILLCELL_X2 FILLER_100_1255 ();
 FILLCELL_X1 FILLER_100_1257 ();
 FILLCELL_X2 FILLER_100_1262 ();
 FILLCELL_X1 FILLER_100_1270 ();
 FILLCELL_X1 FILLER_100_1277 ();
 FILLCELL_X4 FILLER_100_1311 ();
 FILLCELL_X2 FILLER_100_1337 ();
 FILLCELL_X1 FILLER_100_1339 ();
 FILLCELL_X4 FILLER_100_1362 ();
 FILLCELL_X4 FILLER_100_1376 ();
 FILLCELL_X1 FILLER_100_1380 ();
 FILLCELL_X1 FILLER_100_1433 ();
 FILLCELL_X4 FILLER_100_1440 ();
 FILLCELL_X4 FILLER_100_1451 ();
 FILLCELL_X2 FILLER_100_1455 ();
 FILLCELL_X2 FILLER_100_1468 ();
 FILLCELL_X2 FILLER_100_1477 ();
 FILLCELL_X1 FILLER_100_1479 ();
 FILLCELL_X1 FILLER_100_1485 ();
 FILLCELL_X2 FILLER_100_1493 ();
 FILLCELL_X1 FILLER_100_1495 ();
 FILLCELL_X1 FILLER_100_1507 ();
 FILLCELL_X1 FILLER_100_1513 ();
 FILLCELL_X8 FILLER_100_1527 ();
 FILLCELL_X4 FILLER_100_1535 ();
 FILLCELL_X1 FILLER_100_1539 ();
 FILLCELL_X16 FILLER_100_1549 ();
 FILLCELL_X2 FILLER_100_1574 ();
 FILLCELL_X1 FILLER_100_1576 ();
 FILLCELL_X8 FILLER_100_1588 ();
 FILLCELL_X2 FILLER_100_1596 ();
 FILLCELL_X1 FILLER_100_1598 ();
 FILLCELL_X2 FILLER_100_1603 ();
 FILLCELL_X32 FILLER_100_1610 ();
 FILLCELL_X8 FILLER_100_1642 ();
 FILLCELL_X1 FILLER_100_1650 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X2 FILLER_101_33 ();
 FILLCELL_X1 FILLER_101_35 ();
 FILLCELL_X2 FILLER_101_63 ();
 FILLCELL_X8 FILLER_101_76 ();
 FILLCELL_X4 FILLER_101_84 ();
 FILLCELL_X1 FILLER_101_88 ();
 FILLCELL_X2 FILLER_101_102 ();
 FILLCELL_X2 FILLER_101_124 ();
 FILLCELL_X1 FILLER_101_166 ();
 FILLCELL_X8 FILLER_101_187 ();
 FILLCELL_X1 FILLER_101_222 ();
 FILLCELL_X1 FILLER_101_243 ();
 FILLCELL_X4 FILLER_101_248 ();
 FILLCELL_X1 FILLER_101_266 ();
 FILLCELL_X2 FILLER_101_274 ();
 FILLCELL_X2 FILLER_101_285 ();
 FILLCELL_X1 FILLER_101_287 ();
 FILLCELL_X2 FILLER_101_308 ();
 FILLCELL_X1 FILLER_101_310 ();
 FILLCELL_X2 FILLER_101_349 ();
 FILLCELL_X4 FILLER_101_371 ();
 FILLCELL_X8 FILLER_101_395 ();
 FILLCELL_X4 FILLER_101_423 ();
 FILLCELL_X4 FILLER_101_431 ();
 FILLCELL_X4 FILLER_101_448 ();
 FILLCELL_X2 FILLER_101_455 ();
 FILLCELL_X1 FILLER_101_457 ();
 FILLCELL_X4 FILLER_101_460 ();
 FILLCELL_X2 FILLER_101_464 ();
 FILLCELL_X8 FILLER_101_475 ();
 FILLCELL_X1 FILLER_101_489 ();
 FILLCELL_X1 FILLER_101_495 ();
 FILLCELL_X16 FILLER_101_500 ();
 FILLCELL_X2 FILLER_101_516 ();
 FILLCELL_X1 FILLER_101_518 ();
 FILLCELL_X4 FILLER_101_534 ();
 FILLCELL_X2 FILLER_101_538 ();
 FILLCELL_X1 FILLER_101_540 ();
 FILLCELL_X8 FILLER_101_548 ();
 FILLCELL_X4 FILLER_101_556 ();
 FILLCELL_X2 FILLER_101_560 ();
 FILLCELL_X2 FILLER_101_591 ();
 FILLCELL_X1 FILLER_101_600 ();
 FILLCELL_X2 FILLER_101_630 ();
 FILLCELL_X1 FILLER_101_632 ();
 FILLCELL_X2 FILLER_101_732 ();
 FILLCELL_X1 FILLER_101_734 ();
 FILLCELL_X1 FILLER_101_737 ();
 FILLCELL_X2 FILLER_101_747 ();
 FILLCELL_X1 FILLER_101_749 ();
 FILLCELL_X4 FILLER_101_753 ();
 FILLCELL_X1 FILLER_101_790 ();
 FILLCELL_X16 FILLER_101_799 ();
 FILLCELL_X2 FILLER_101_815 ();
 FILLCELL_X4 FILLER_101_824 ();
 FILLCELL_X2 FILLER_101_828 ();
 FILLCELL_X8 FILLER_101_852 ();
 FILLCELL_X4 FILLER_101_867 ();
 FILLCELL_X2 FILLER_101_878 ();
 FILLCELL_X1 FILLER_101_887 ();
 FILLCELL_X2 FILLER_101_893 ();
 FILLCELL_X8 FILLER_101_917 ();
 FILLCELL_X4 FILLER_101_932 ();
 FILLCELL_X2 FILLER_101_936 ();
 FILLCELL_X2 FILLER_101_943 ();
 FILLCELL_X1 FILLER_101_945 ();
 FILLCELL_X4 FILLER_101_965 ();
 FILLCELL_X2 FILLER_101_969 ();
 FILLCELL_X1 FILLER_101_971 ();
 FILLCELL_X4 FILLER_101_984 ();
 FILLCELL_X32 FILLER_101_994 ();
 FILLCELL_X4 FILLER_101_1026 ();
 FILLCELL_X4 FILLER_101_1039 ();
 FILLCELL_X2 FILLER_101_1043 ();
 FILLCELL_X4 FILLER_101_1061 ();
 FILLCELL_X2 FILLER_101_1065 ();
 FILLCELL_X16 FILLER_101_1072 ();
 FILLCELL_X1 FILLER_101_1088 ();
 FILLCELL_X2 FILLER_101_1095 ();
 FILLCELL_X4 FILLER_101_1102 ();
 FILLCELL_X8 FILLER_101_1133 ();
 FILLCELL_X2 FILLER_101_1186 ();
 FILLCELL_X1 FILLER_101_1188 ();
 FILLCELL_X4 FILLER_101_1199 ();
 FILLCELL_X2 FILLER_101_1203 ();
 FILLCELL_X4 FILLER_101_1222 ();
 FILLCELL_X4 FILLER_101_1232 ();
 FILLCELL_X2 FILLER_101_1238 ();
 FILLCELL_X1 FILLER_101_1240 ();
 FILLCELL_X2 FILLER_101_1261 ();
 FILLCELL_X8 FILLER_101_1264 ();
 FILLCELL_X1 FILLER_101_1272 ();
 FILLCELL_X1 FILLER_101_1277 ();
 FILLCELL_X2 FILLER_101_1303 ();
 FILLCELL_X1 FILLER_101_1305 ();
 FILLCELL_X1 FILLER_101_1326 ();
 FILLCELL_X8 FILLER_101_1329 ();
 FILLCELL_X4 FILLER_101_1337 ();
 FILLCELL_X2 FILLER_101_1341 ();
 FILLCELL_X1 FILLER_101_1343 ();
 FILLCELL_X4 FILLER_101_1362 ();
 FILLCELL_X2 FILLER_101_1369 ();
 FILLCELL_X1 FILLER_101_1371 ();
 FILLCELL_X2 FILLER_101_1382 ();
 FILLCELL_X1 FILLER_101_1384 ();
 FILLCELL_X2 FILLER_101_1391 ();
 FILLCELL_X4 FILLER_101_1399 ();
 FILLCELL_X1 FILLER_101_1409 ();
 FILLCELL_X2 FILLER_101_1416 ();
 FILLCELL_X16 FILLER_101_1440 ();
 FILLCELL_X4 FILLER_101_1456 ();
 FILLCELL_X2 FILLER_101_1460 ();
 FILLCELL_X4 FILLER_101_1465 ();
 FILLCELL_X2 FILLER_101_1469 ();
 FILLCELL_X2 FILLER_101_1482 ();
 FILLCELL_X2 FILLER_101_1501 ();
 FILLCELL_X2 FILLER_101_1507 ();
 FILLCELL_X2 FILLER_101_1523 ();
 FILLCELL_X1 FILLER_101_1542 ();
 FILLCELL_X1 FILLER_101_1554 ();
 FILLCELL_X2 FILLER_101_1572 ();
 FILLCELL_X4 FILLER_101_1586 ();
 FILLCELL_X1 FILLER_101_1590 ();
 FILLCELL_X2 FILLER_101_1599 ();
 FILLCELL_X32 FILLER_101_1612 ();
 FILLCELL_X4 FILLER_101_1644 ();
 FILLCELL_X2 FILLER_101_1648 ();
 FILLCELL_X1 FILLER_101_1650 ();
 FILLCELL_X16 FILLER_102_1 ();
 FILLCELL_X2 FILLER_102_17 ();
 FILLCELL_X1 FILLER_102_19 ();
 FILLCELL_X2 FILLER_102_47 ();
 FILLCELL_X4 FILLER_102_106 ();
 FILLCELL_X1 FILLER_102_110 ();
 FILLCELL_X2 FILLER_102_116 ();
 FILLCELL_X1 FILLER_102_118 ();
 FILLCELL_X2 FILLER_102_127 ();
 FILLCELL_X8 FILLER_102_136 ();
 FILLCELL_X1 FILLER_102_144 ();
 FILLCELL_X8 FILLER_102_150 ();
 FILLCELL_X4 FILLER_102_158 ();
 FILLCELL_X2 FILLER_102_162 ();
 FILLCELL_X1 FILLER_102_164 ();
 FILLCELL_X4 FILLER_102_170 ();
 FILLCELL_X1 FILLER_102_174 ();
 FILLCELL_X1 FILLER_102_182 ();
 FILLCELL_X16 FILLER_102_188 ();
 FILLCELL_X2 FILLER_102_204 ();
 FILLCELL_X4 FILLER_102_213 ();
 FILLCELL_X16 FILLER_102_242 ();
 FILLCELL_X2 FILLER_102_258 ();
 FILLCELL_X2 FILLER_102_269 ();
 FILLCELL_X1 FILLER_102_271 ();
 FILLCELL_X2 FILLER_102_277 ();
 FILLCELL_X1 FILLER_102_286 ();
 FILLCELL_X4 FILLER_102_294 ();
 FILLCELL_X2 FILLER_102_298 ();
 FILLCELL_X1 FILLER_102_300 ();
 FILLCELL_X16 FILLER_102_364 ();
 FILLCELL_X2 FILLER_102_380 ();
 FILLCELL_X2 FILLER_102_391 ();
 FILLCELL_X8 FILLER_102_419 ();
 FILLCELL_X2 FILLER_102_427 ();
 FILLCELL_X1 FILLER_102_429 ();
 FILLCELL_X4 FILLER_102_439 ();
 FILLCELL_X2 FILLER_102_448 ();
 FILLCELL_X1 FILLER_102_450 ();
 FILLCELL_X2 FILLER_102_464 ();
 FILLCELL_X1 FILLER_102_475 ();
 FILLCELL_X1 FILLER_102_522 ();
 FILLCELL_X2 FILLER_102_527 ();
 FILLCELL_X8 FILLER_102_531 ();
 FILLCELL_X2 FILLER_102_539 ();
 FILLCELL_X8 FILLER_102_545 ();
 FILLCELL_X2 FILLER_102_553 ();
 FILLCELL_X16 FILLER_102_562 ();
 FILLCELL_X4 FILLER_102_578 ();
 FILLCELL_X1 FILLER_102_582 ();
 FILLCELL_X1 FILLER_102_587 ();
 FILLCELL_X16 FILLER_102_608 ();
 FILLCELL_X4 FILLER_102_624 ();
 FILLCELL_X2 FILLER_102_628 ();
 FILLCELL_X1 FILLER_102_630 ();
 FILLCELL_X8 FILLER_102_632 ();
 FILLCELL_X4 FILLER_102_711 ();
 FILLCELL_X1 FILLER_102_715 ();
 FILLCELL_X8 FILLER_102_751 ();
 FILLCELL_X4 FILLER_102_767 ();
 FILLCELL_X2 FILLER_102_775 ();
 FILLCELL_X1 FILLER_102_777 ();
 FILLCELL_X2 FILLER_102_780 ();
 FILLCELL_X1 FILLER_102_782 ();
 FILLCELL_X8 FILLER_102_796 ();
 FILLCELL_X2 FILLER_102_808 ();
 FILLCELL_X1 FILLER_102_810 ();
 FILLCELL_X16 FILLER_102_833 ();
 FILLCELL_X2 FILLER_102_849 ();
 FILLCELL_X2 FILLER_102_858 ();
 FILLCELL_X8 FILLER_102_902 ();
 FILLCELL_X2 FILLER_102_917 ();
 FILLCELL_X1 FILLER_102_924 ();
 FILLCELL_X8 FILLER_102_957 ();
 FILLCELL_X4 FILLER_102_965 ();
 FILLCELL_X2 FILLER_102_969 ();
 FILLCELL_X1 FILLER_102_971 ();
 FILLCELL_X2 FILLER_102_982 ();
 FILLCELL_X1 FILLER_102_984 ();
 FILLCELL_X2 FILLER_102_996 ();
 FILLCELL_X4 FILLER_102_1003 ();
 FILLCELL_X2 FILLER_102_1007 ();
 FILLCELL_X4 FILLER_102_1016 ();
 FILLCELL_X1 FILLER_102_1020 ();
 FILLCELL_X8 FILLER_102_1039 ();
 FILLCELL_X4 FILLER_102_1047 ();
 FILLCELL_X1 FILLER_102_1051 ();
 FILLCELL_X4 FILLER_102_1121 ();
 FILLCELL_X2 FILLER_102_1125 ();
 FILLCELL_X8 FILLER_102_1137 ();
 FILLCELL_X8 FILLER_102_1162 ();
 FILLCELL_X2 FILLER_102_1170 ();
 FILLCELL_X1 FILLER_102_1172 ();
 FILLCELL_X1 FILLER_102_1207 ();
 FILLCELL_X2 FILLER_102_1230 ();
 FILLCELL_X1 FILLER_102_1232 ();
 FILLCELL_X4 FILLER_102_1264 ();
 FILLCELL_X2 FILLER_102_1268 ();
 FILLCELL_X4 FILLER_102_1284 ();
 FILLCELL_X2 FILLER_102_1288 ();
 FILLCELL_X2 FILLER_102_1300 ();
 FILLCELL_X4 FILLER_102_1312 ();
 FILLCELL_X1 FILLER_102_1320 ();
 FILLCELL_X8 FILLER_102_1343 ();
 FILLCELL_X4 FILLER_102_1351 ();
 FILLCELL_X2 FILLER_102_1397 ();
 FILLCELL_X2 FILLER_102_1405 ();
 FILLCELL_X1 FILLER_102_1417 ();
 FILLCELL_X2 FILLER_102_1424 ();
 FILLCELL_X32 FILLER_102_1432 ();
 FILLCELL_X32 FILLER_102_1464 ();
 FILLCELL_X4 FILLER_102_1496 ();
 FILLCELL_X8 FILLER_102_1503 ();
 FILLCELL_X2 FILLER_102_1511 ();
 FILLCELL_X1 FILLER_102_1513 ();
 FILLCELL_X1 FILLER_102_1518 ();
 FILLCELL_X8 FILLER_102_1528 ();
 FILLCELL_X4 FILLER_102_1536 ();
 FILLCELL_X2 FILLER_102_1540 ();
 FILLCELL_X1 FILLER_102_1542 ();
 FILLCELL_X1 FILLER_102_1547 ();
 FILLCELL_X4 FILLER_102_1553 ();
 FILLCELL_X4 FILLER_102_1572 ();
 FILLCELL_X4 FILLER_102_1580 ();
 FILLCELL_X2 FILLER_102_1584 ();
 FILLCELL_X32 FILLER_102_1593 ();
 FILLCELL_X16 FILLER_102_1625 ();
 FILLCELL_X8 FILLER_102_1641 ();
 FILLCELL_X2 FILLER_102_1649 ();
 FILLCELL_X16 FILLER_103_1 ();
 FILLCELL_X8 FILLER_103_17 ();
 FILLCELL_X2 FILLER_103_25 ();
 FILLCELL_X4 FILLER_103_79 ();
 FILLCELL_X2 FILLER_103_83 ();
 FILLCELL_X1 FILLER_103_85 ();
 FILLCELL_X1 FILLER_103_95 ();
 FILLCELL_X4 FILLER_103_105 ();
 FILLCELL_X2 FILLER_103_109 ();
 FILLCELL_X1 FILLER_103_143 ();
 FILLCELL_X8 FILLER_103_148 ();
 FILLCELL_X1 FILLER_103_156 ();
 FILLCELL_X8 FILLER_103_164 ();
 FILLCELL_X4 FILLER_103_172 ();
 FILLCELL_X2 FILLER_103_179 ();
 FILLCELL_X2 FILLER_103_190 ();
 FILLCELL_X1 FILLER_103_192 ();
 FILLCELL_X4 FILLER_103_200 ();
 FILLCELL_X4 FILLER_103_229 ();
 FILLCELL_X2 FILLER_103_233 ();
 FILLCELL_X8 FILLER_103_240 ();
 FILLCELL_X4 FILLER_103_248 ();
 FILLCELL_X1 FILLER_103_295 ();
 FILLCELL_X2 FILLER_103_300 ();
 FILLCELL_X1 FILLER_103_302 ();
 FILLCELL_X1 FILLER_103_322 ();
 FILLCELL_X16 FILLER_103_340 ();
 FILLCELL_X8 FILLER_103_356 ();
 FILLCELL_X1 FILLER_103_364 ();
 FILLCELL_X1 FILLER_103_368 ();
 FILLCELL_X1 FILLER_103_385 ();
 FILLCELL_X2 FILLER_103_394 ();
 FILLCELL_X1 FILLER_103_396 ();
 FILLCELL_X4 FILLER_103_399 ();
 FILLCELL_X2 FILLER_103_403 ();
 FILLCELL_X1 FILLER_103_405 ();
 FILLCELL_X1 FILLER_103_450 ();
 FILLCELL_X8 FILLER_103_455 ();
 FILLCELL_X1 FILLER_103_472 ();
 FILLCELL_X2 FILLER_103_502 ();
 FILLCELL_X2 FILLER_103_508 ();
 FILLCELL_X2 FILLER_103_515 ();
 FILLCELL_X4 FILLER_103_537 ();
 FILLCELL_X1 FILLER_103_541 ();
 FILLCELL_X4 FILLER_103_544 ();
 FILLCELL_X4 FILLER_103_575 ();
 FILLCELL_X2 FILLER_103_579 ();
 FILLCELL_X8 FILLER_103_586 ();
 FILLCELL_X4 FILLER_103_598 ();
 FILLCELL_X2 FILLER_103_602 ();
 FILLCELL_X1 FILLER_103_604 ();
 FILLCELL_X1 FILLER_103_610 ();
 FILLCELL_X8 FILLER_103_616 ();
 FILLCELL_X2 FILLER_103_624 ();
 FILLCELL_X8 FILLER_103_633 ();
 FILLCELL_X8 FILLER_103_648 ();
 FILLCELL_X4 FILLER_103_661 ();
 FILLCELL_X2 FILLER_103_669 ();
 FILLCELL_X4 FILLER_103_702 ();
 FILLCELL_X1 FILLER_103_706 ();
 FILLCELL_X8 FILLER_103_718 ();
 FILLCELL_X4 FILLER_103_797 ();
 FILLCELL_X2 FILLER_103_801 ();
 FILLCELL_X1 FILLER_103_823 ();
 FILLCELL_X1 FILLER_103_871 ();
 FILLCELL_X8 FILLER_103_879 ();
 FILLCELL_X16 FILLER_103_916 ();
 FILLCELL_X8 FILLER_103_932 ();
 FILLCELL_X4 FILLER_103_940 ();
 FILLCELL_X2 FILLER_103_944 ();
 FILLCELL_X2 FILLER_103_952 ();
 FILLCELL_X16 FILLER_103_959 ();
 FILLCELL_X1 FILLER_103_975 ();
 FILLCELL_X4 FILLER_103_986 ();
 FILLCELL_X2 FILLER_103_1001 ();
 FILLCELL_X1 FILLER_103_1003 ();
 FILLCELL_X1 FILLER_103_1033 ();
 FILLCELL_X4 FILLER_103_1041 ();
 FILLCELL_X2 FILLER_103_1050 ();
 FILLCELL_X2 FILLER_103_1057 ();
 FILLCELL_X1 FILLER_103_1059 ();
 FILLCELL_X4 FILLER_103_1088 ();
 FILLCELL_X2 FILLER_103_1092 ();
 FILLCELL_X2 FILLER_103_1103 ();
 FILLCELL_X1 FILLER_103_1105 ();
 FILLCELL_X8 FILLER_103_1128 ();
 FILLCELL_X4 FILLER_103_1136 ();
 FILLCELL_X2 FILLER_103_1140 ();
 FILLCELL_X16 FILLER_103_1164 ();
 FILLCELL_X1 FILLER_103_1180 ();
 FILLCELL_X4 FILLER_103_1217 ();
 FILLCELL_X2 FILLER_103_1221 ();
 FILLCELL_X4 FILLER_103_1243 ();
 FILLCELL_X1 FILLER_103_1247 ();
 FILLCELL_X1 FILLER_103_1264 ();
 FILLCELL_X8 FILLER_103_1271 ();
 FILLCELL_X8 FILLER_103_1290 ();
 FILLCELL_X4 FILLER_103_1298 ();
 FILLCELL_X1 FILLER_103_1302 ();
 FILLCELL_X2 FILLER_103_1328 ();
 FILLCELL_X1 FILLER_103_1359 ();
 FILLCELL_X1 FILLER_103_1382 ();
 FILLCELL_X1 FILLER_103_1395 ();
 FILLCELL_X1 FILLER_103_1402 ();
 FILLCELL_X2 FILLER_103_1413 ();
 FILLCELL_X32 FILLER_103_1425 ();
 FILLCELL_X8 FILLER_103_1457 ();
 FILLCELL_X2 FILLER_103_1465 ();
 FILLCELL_X1 FILLER_103_1467 ();
 FILLCELL_X32 FILLER_103_1471 ();
 FILLCELL_X8 FILLER_103_1503 ();
 FILLCELL_X4 FILLER_103_1511 ();
 FILLCELL_X2 FILLER_103_1518 ();
 FILLCELL_X1 FILLER_103_1520 ();
 FILLCELL_X4 FILLER_103_1525 ();
 FILLCELL_X8 FILLER_103_1533 ();
 FILLCELL_X2 FILLER_103_1541 ();
 FILLCELL_X4 FILLER_103_1546 ();
 FILLCELL_X2 FILLER_103_1550 ();
 FILLCELL_X1 FILLER_103_1552 ();
 FILLCELL_X4 FILLER_103_1560 ();
 FILLCELL_X2 FILLER_103_1564 ();
 FILLCELL_X1 FILLER_103_1566 ();
 FILLCELL_X8 FILLER_103_1574 ();
 FILLCELL_X1 FILLER_103_1594 ();
 FILLCELL_X4 FILLER_103_1599 ();
 FILLCELL_X1 FILLER_103_1603 ();
 FILLCELL_X32 FILLER_103_1615 ();
 FILLCELL_X4 FILLER_103_1647 ();
 FILLCELL_X16 FILLER_104_1 ();
 FILLCELL_X8 FILLER_104_17 ();
 FILLCELL_X4 FILLER_104_25 ();
 FILLCELL_X1 FILLER_104_29 ();
 FILLCELL_X8 FILLER_104_37 ();
 FILLCELL_X2 FILLER_104_45 ();
 FILLCELL_X4 FILLER_104_54 ();
 FILLCELL_X2 FILLER_104_58 ();
 FILLCELL_X1 FILLER_104_60 ();
 FILLCELL_X16 FILLER_104_70 ();
 FILLCELL_X4 FILLER_104_86 ();
 FILLCELL_X4 FILLER_104_94 ();
 FILLCELL_X2 FILLER_104_98 ();
 FILLCELL_X1 FILLER_104_100 ();
 FILLCELL_X2 FILLER_104_108 ();
 FILLCELL_X1 FILLER_104_110 ();
 FILLCELL_X1 FILLER_104_118 ();
 FILLCELL_X1 FILLER_104_124 ();
 FILLCELL_X8 FILLER_104_150 ();
 FILLCELL_X2 FILLER_104_158 ();
 FILLCELL_X1 FILLER_104_160 ();
 FILLCELL_X2 FILLER_104_211 ();
 FILLCELL_X2 FILLER_104_225 ();
 FILLCELL_X1 FILLER_104_274 ();
 FILLCELL_X1 FILLER_104_295 ();
 FILLCELL_X2 FILLER_104_333 ();
 FILLCELL_X2 FILLER_104_344 ();
 FILLCELL_X1 FILLER_104_346 ();
 FILLCELL_X4 FILLER_104_397 ();
 FILLCELL_X1 FILLER_104_401 ();
 FILLCELL_X2 FILLER_104_406 ();
 FILLCELL_X1 FILLER_104_408 ();
 FILLCELL_X8 FILLER_104_414 ();
 FILLCELL_X4 FILLER_104_422 ();
 FILLCELL_X1 FILLER_104_426 ();
 FILLCELL_X1 FILLER_104_439 ();
 FILLCELL_X1 FILLER_104_462 ();
 FILLCELL_X2 FILLER_104_469 ();
 FILLCELL_X16 FILLER_104_475 ();
 FILLCELL_X4 FILLER_104_491 ();
 FILLCELL_X1 FILLER_104_495 ();
 FILLCELL_X4 FILLER_104_499 ();
 FILLCELL_X2 FILLER_104_503 ();
 FILLCELL_X4 FILLER_104_509 ();
 FILLCELL_X1 FILLER_104_513 ();
 FILLCELL_X2 FILLER_104_547 ();
 FILLCELL_X1 FILLER_104_549 ();
 FILLCELL_X2 FILLER_104_563 ();
 FILLCELL_X4 FILLER_104_578 ();
 FILLCELL_X1 FILLER_104_582 ();
 FILLCELL_X2 FILLER_104_590 ();
 FILLCELL_X4 FILLER_104_606 ();
 FILLCELL_X1 FILLER_104_610 ();
 FILLCELL_X4 FILLER_104_620 ();
 FILLCELL_X1 FILLER_104_632 ();
 FILLCELL_X1 FILLER_104_675 ();
 FILLCELL_X2 FILLER_104_691 ();
 FILLCELL_X1 FILLER_104_706 ();
 FILLCELL_X32 FILLER_104_729 ();
 FILLCELL_X2 FILLER_104_774 ();
 FILLCELL_X4 FILLER_104_789 ();
 FILLCELL_X4 FILLER_104_797 ();
 FILLCELL_X8 FILLER_104_806 ();
 FILLCELL_X1 FILLER_104_814 ();
 FILLCELL_X4 FILLER_104_819 ();
 FILLCELL_X16 FILLER_104_834 ();
 FILLCELL_X4 FILLER_104_850 ();
 FILLCELL_X2 FILLER_104_854 ();
 FILLCELL_X8 FILLER_104_863 ();
 FILLCELL_X2 FILLER_104_871 ();
 FILLCELL_X1 FILLER_104_873 ();
 FILLCELL_X16 FILLER_104_896 ();
 FILLCELL_X32 FILLER_104_917 ();
 FILLCELL_X8 FILLER_104_949 ();
 FILLCELL_X4 FILLER_104_957 ();
 FILLCELL_X2 FILLER_104_961 ();
 FILLCELL_X1 FILLER_104_963 ();
 FILLCELL_X8 FILLER_104_971 ();
 FILLCELL_X2 FILLER_104_979 ();
 FILLCELL_X4 FILLER_104_988 ();
 FILLCELL_X8 FILLER_104_1001 ();
 FILLCELL_X4 FILLER_104_1009 ();
 FILLCELL_X1 FILLER_104_1038 ();
 FILLCELL_X1 FILLER_104_1064 ();
 FILLCELL_X4 FILLER_104_1069 ();
 FILLCELL_X8 FILLER_104_1102 ();
 FILLCELL_X2 FILLER_104_1110 ();
 FILLCELL_X1 FILLER_104_1112 ();
 FILLCELL_X16 FILLER_104_1123 ();
 FILLCELL_X4 FILLER_104_1139 ();
 FILLCELL_X1 FILLER_104_1143 ();
 FILLCELL_X4 FILLER_104_1177 ();
 FILLCELL_X1 FILLER_104_1181 ();
 FILLCELL_X4 FILLER_104_1187 ();
 FILLCELL_X4 FILLER_104_1201 ();
 FILLCELL_X1 FILLER_104_1205 ();
 FILLCELL_X2 FILLER_104_1225 ();
 FILLCELL_X4 FILLER_104_1235 ();
 FILLCELL_X8 FILLER_104_1244 ();
 FILLCELL_X2 FILLER_104_1269 ();
 FILLCELL_X8 FILLER_104_1278 ();
 FILLCELL_X4 FILLER_104_1286 ();
 FILLCELL_X1 FILLER_104_1296 ();
 FILLCELL_X2 FILLER_104_1307 ();
 FILLCELL_X4 FILLER_104_1313 ();
 FILLCELL_X1 FILLER_104_1317 ();
 FILLCELL_X2 FILLER_104_1323 ();
 FILLCELL_X4 FILLER_104_1351 ();
 FILLCELL_X2 FILLER_104_1355 ();
 FILLCELL_X1 FILLER_104_1357 ();
 FILLCELL_X2 FILLER_104_1362 ();
 FILLCELL_X8 FILLER_104_1371 ();
 FILLCELL_X4 FILLER_104_1389 ();
 FILLCELL_X1 FILLER_104_1399 ();
 FILLCELL_X2 FILLER_104_1406 ();
 FILLCELL_X1 FILLER_104_1418 ();
 FILLCELL_X32 FILLER_104_1425 ();
 FILLCELL_X16 FILLER_104_1457 ();
 FILLCELL_X4 FILLER_104_1473 ();
 FILLCELL_X4 FILLER_104_1487 ();
 FILLCELL_X1 FILLER_104_1495 ();
 FILLCELL_X2 FILLER_104_1500 ();
 FILLCELL_X2 FILLER_104_1506 ();
 FILLCELL_X2 FILLER_104_1512 ();
 FILLCELL_X1 FILLER_104_1514 ();
 FILLCELL_X2 FILLER_104_1540 ();
 FILLCELL_X8 FILLER_104_1546 ();
 FILLCELL_X8 FILLER_104_1559 ();
 FILLCELL_X2 FILLER_104_1567 ();
 FILLCELL_X1 FILLER_104_1569 ();
 FILLCELL_X32 FILLER_104_1576 ();
 FILLCELL_X32 FILLER_104_1608 ();
 FILLCELL_X8 FILLER_104_1640 ();
 FILLCELL_X2 FILLER_104_1648 ();
 FILLCELL_X1 FILLER_104_1650 ();
 FILLCELL_X8 FILLER_105_1 ();
 FILLCELL_X4 FILLER_105_9 ();
 FILLCELL_X1 FILLER_105_13 ();
 FILLCELL_X4 FILLER_105_48 ();
 FILLCELL_X4 FILLER_105_59 ();
 FILLCELL_X2 FILLER_105_63 ();
 FILLCELL_X1 FILLER_105_105 ();
 FILLCELL_X8 FILLER_105_133 ();
 FILLCELL_X4 FILLER_105_141 ();
 FILLCELL_X2 FILLER_105_145 ();
 FILLCELL_X1 FILLER_105_160 ();
 FILLCELL_X2 FILLER_105_168 ();
 FILLCELL_X8 FILLER_105_197 ();
 FILLCELL_X1 FILLER_105_205 ();
 FILLCELL_X4 FILLER_105_231 ();
 FILLCELL_X16 FILLER_105_242 ();
 FILLCELL_X16 FILLER_105_263 ();
 FILLCELL_X2 FILLER_105_279 ();
 FILLCELL_X1 FILLER_105_359 ();
 FILLCELL_X8 FILLER_105_393 ();
 FILLCELL_X1 FILLER_105_401 ();
 FILLCELL_X1 FILLER_105_421 ();
 FILLCELL_X1 FILLER_105_467 ();
 FILLCELL_X1 FILLER_105_482 ();
 FILLCELL_X1 FILLER_105_496 ();
 FILLCELL_X1 FILLER_105_524 ();
 FILLCELL_X2 FILLER_105_529 ();
 FILLCELL_X1 FILLER_105_531 ();
 FILLCELL_X8 FILLER_105_534 ();
 FILLCELL_X2 FILLER_105_542 ();
 FILLCELL_X1 FILLER_105_544 ();
 FILLCELL_X1 FILLER_105_548 ();
 FILLCELL_X2 FILLER_105_553 ();
 FILLCELL_X1 FILLER_105_555 ();
 FILLCELL_X1 FILLER_105_569 ();
 FILLCELL_X2 FILLER_105_574 ();
 FILLCELL_X1 FILLER_105_593 ();
 FILLCELL_X8 FILLER_105_597 ();
 FILLCELL_X1 FILLER_105_605 ();
 FILLCELL_X2 FILLER_105_609 ();
 FILLCELL_X8 FILLER_105_639 ();
 FILLCELL_X2 FILLER_105_647 ();
 FILLCELL_X2 FILLER_105_662 ();
 FILLCELL_X4 FILLER_105_669 ();
 FILLCELL_X1 FILLER_105_673 ();
 FILLCELL_X16 FILLER_105_687 ();
 FILLCELL_X8 FILLER_105_703 ();
 FILLCELL_X1 FILLER_105_711 ();
 FILLCELL_X2 FILLER_105_746 ();
 FILLCELL_X4 FILLER_105_750 ();
 FILLCELL_X1 FILLER_105_754 ();
 FILLCELL_X4 FILLER_105_789 ();
 FILLCELL_X1 FILLER_105_841 ();
 FILLCELL_X1 FILLER_105_844 ();
 FILLCELL_X1 FILLER_105_848 ();
 FILLCELL_X2 FILLER_105_856 ();
 FILLCELL_X1 FILLER_105_880 ();
 FILLCELL_X2 FILLER_105_888 ();
 FILLCELL_X1 FILLER_105_905 ();
 FILLCELL_X8 FILLER_105_942 ();
 FILLCELL_X4 FILLER_105_950 ();
 FILLCELL_X2 FILLER_105_954 ();
 FILLCELL_X1 FILLER_105_956 ();
 FILLCELL_X1 FILLER_105_979 ();
 FILLCELL_X8 FILLER_105_987 ();
 FILLCELL_X4 FILLER_105_995 ();
 FILLCELL_X8 FILLER_105_1001 ();
 FILLCELL_X4 FILLER_105_1009 ();
 FILLCELL_X2 FILLER_105_1013 ();
 FILLCELL_X8 FILLER_105_1023 ();
 FILLCELL_X4 FILLER_105_1031 ();
 FILLCELL_X2 FILLER_105_1035 ();
 FILLCELL_X4 FILLER_105_1045 ();
 FILLCELL_X2 FILLER_105_1049 ();
 FILLCELL_X1 FILLER_105_1056 ();
 FILLCELL_X1 FILLER_105_1060 ();
 FILLCELL_X1 FILLER_105_1065 ();
 FILLCELL_X1 FILLER_105_1073 ();
 FILLCELL_X16 FILLER_105_1079 ();
 FILLCELL_X2 FILLER_105_1095 ();
 FILLCELL_X1 FILLER_105_1097 ();
 FILLCELL_X1 FILLER_105_1140 ();
 FILLCELL_X1 FILLER_105_1160 ();
 FILLCELL_X4 FILLER_105_1216 ();
 FILLCELL_X1 FILLER_105_1226 ();
 FILLCELL_X4 FILLER_105_1252 ();
 FILLCELL_X1 FILLER_105_1262 ();
 FILLCELL_X2 FILLER_105_1264 ();
 FILLCELL_X2 FILLER_105_1295 ();
 FILLCELL_X1 FILLER_105_1297 ();
 FILLCELL_X4 FILLER_105_1303 ();
 FILLCELL_X1 FILLER_105_1307 ();
 FILLCELL_X16 FILLER_105_1319 ();
 FILLCELL_X4 FILLER_105_1335 ();
 FILLCELL_X8 FILLER_105_1354 ();
 FILLCELL_X2 FILLER_105_1362 ();
 FILLCELL_X1 FILLER_105_1364 ();
 FILLCELL_X8 FILLER_105_1387 ();
 FILLCELL_X4 FILLER_105_1395 ();
 FILLCELL_X2 FILLER_105_1399 ();
 FILLCELL_X2 FILLER_105_1411 ();
 FILLCELL_X1 FILLER_105_1413 ();
 FILLCELL_X32 FILLER_105_1440 ();
 FILLCELL_X8 FILLER_105_1472 ();
 FILLCELL_X4 FILLER_105_1480 ();
 FILLCELL_X2 FILLER_105_1484 ();
 FILLCELL_X1 FILLER_105_1486 ();
 FILLCELL_X16 FILLER_105_1498 ();
 FILLCELL_X4 FILLER_105_1514 ();
 FILLCELL_X16 FILLER_105_1523 ();
 FILLCELL_X4 FILLER_105_1539 ();
 FILLCELL_X1 FILLER_105_1543 ();
 FILLCELL_X8 FILLER_105_1547 ();
 FILLCELL_X4 FILLER_105_1555 ();
 FILLCELL_X1 FILLER_105_1559 ();
 FILLCELL_X32 FILLER_105_1570 ();
 FILLCELL_X32 FILLER_105_1602 ();
 FILLCELL_X16 FILLER_105_1634 ();
 FILLCELL_X1 FILLER_105_1650 ();
 FILLCELL_X8 FILLER_106_1 ();
 FILLCELL_X2 FILLER_106_9 ();
 FILLCELL_X1 FILLER_106_11 ();
 FILLCELL_X1 FILLER_106_32 ();
 FILLCELL_X2 FILLER_106_40 ();
 FILLCELL_X2 FILLER_106_49 ();
 FILLCELL_X2 FILLER_106_60 ();
 FILLCELL_X1 FILLER_106_62 ();
 FILLCELL_X8 FILLER_106_110 ();
 FILLCELL_X2 FILLER_106_123 ();
 FILLCELL_X1 FILLER_106_125 ();
 FILLCELL_X2 FILLER_106_149 ();
 FILLCELL_X1 FILLER_106_151 ();
 FILLCELL_X4 FILLER_106_209 ();
 FILLCELL_X2 FILLER_106_213 ();
 FILLCELL_X1 FILLER_106_215 ();
 FILLCELL_X8 FILLER_106_223 ();
 FILLCELL_X2 FILLER_106_231 ();
 FILLCELL_X4 FILLER_106_241 ();
 FILLCELL_X2 FILLER_106_245 ();
 FILLCELL_X1 FILLER_106_247 ();
 FILLCELL_X4 FILLER_106_275 ();
 FILLCELL_X1 FILLER_106_279 ();
 FILLCELL_X8 FILLER_106_300 ();
 FILLCELL_X4 FILLER_106_308 ();
 FILLCELL_X1 FILLER_106_312 ();
 FILLCELL_X16 FILLER_106_320 ();
 FILLCELL_X4 FILLER_106_336 ();
 FILLCELL_X16 FILLER_106_349 ();
 FILLCELL_X8 FILLER_106_365 ();
 FILLCELL_X2 FILLER_106_373 ();
 FILLCELL_X1 FILLER_106_375 ();
 FILLCELL_X4 FILLER_106_409 ();
 FILLCELL_X2 FILLER_106_413 ();
 FILLCELL_X1 FILLER_106_449 ();
 FILLCELL_X1 FILLER_106_454 ();
 FILLCELL_X4 FILLER_106_460 ();
 FILLCELL_X4 FILLER_106_471 ();
 FILLCELL_X1 FILLER_106_475 ();
 FILLCELL_X16 FILLER_106_503 ();
 FILLCELL_X1 FILLER_106_519 ();
 FILLCELL_X1 FILLER_106_540 ();
 FILLCELL_X4 FILLER_106_563 ();
 FILLCELL_X1 FILLER_106_567 ();
 FILLCELL_X1 FILLER_106_595 ();
 FILLCELL_X8 FILLER_106_600 ();
 FILLCELL_X2 FILLER_106_608 ();
 FILLCELL_X8 FILLER_106_614 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X16 FILLER_106_652 ();
 FILLCELL_X4 FILLER_106_677 ();
 FILLCELL_X1 FILLER_106_681 ();
 FILLCELL_X1 FILLER_106_689 ();
 FILLCELL_X8 FILLER_106_717 ();
 FILLCELL_X4 FILLER_106_725 ();
 FILLCELL_X2 FILLER_106_729 ();
 FILLCELL_X1 FILLER_106_731 ();
 FILLCELL_X4 FILLER_106_735 ();
 FILLCELL_X2 FILLER_106_739 ();
 FILLCELL_X16 FILLER_106_761 ();
 FILLCELL_X1 FILLER_106_777 ();
 FILLCELL_X2 FILLER_106_781 ();
 FILLCELL_X1 FILLER_106_783 ();
 FILLCELL_X4 FILLER_106_797 ();
 FILLCELL_X2 FILLER_106_801 ();
 FILLCELL_X4 FILLER_106_854 ();
 FILLCELL_X4 FILLER_106_887 ();
 FILLCELL_X8 FILLER_106_911 ();
 FILLCELL_X4 FILLER_106_919 ();
 FILLCELL_X2 FILLER_106_923 ();
 FILLCELL_X1 FILLER_106_925 ();
 FILLCELL_X8 FILLER_106_933 ();
 FILLCELL_X4 FILLER_106_941 ();
 FILLCELL_X1 FILLER_106_945 ();
 FILLCELL_X4 FILLER_106_950 ();
 FILLCELL_X1 FILLER_106_954 ();
 FILLCELL_X1 FILLER_106_965 ();
 FILLCELL_X1 FILLER_106_973 ();
 FILLCELL_X2 FILLER_106_985 ();
 FILLCELL_X2 FILLER_106_1008 ();
 FILLCELL_X2 FILLER_106_1017 ();
 FILLCELL_X2 FILLER_106_1032 ();
 FILLCELL_X8 FILLER_106_1037 ();
 FILLCELL_X2 FILLER_106_1045 ();
 FILLCELL_X16 FILLER_106_1050 ();
 FILLCELL_X8 FILLER_106_1071 ();
 FILLCELL_X1 FILLER_106_1079 ();
 FILLCELL_X8 FILLER_106_1090 ();
 FILLCELL_X4 FILLER_106_1098 ();
 FILLCELL_X2 FILLER_106_1138 ();
 FILLCELL_X1 FILLER_106_1140 ();
 FILLCELL_X4 FILLER_106_1149 ();
 FILLCELL_X8 FILLER_106_1156 ();
 FILLCELL_X4 FILLER_106_1164 ();
 FILLCELL_X2 FILLER_106_1168 ();
 FILLCELL_X1 FILLER_106_1170 ();
 FILLCELL_X1 FILLER_106_1177 ();
 FILLCELL_X2 FILLER_106_1188 ();
 FILLCELL_X4 FILLER_106_1195 ();
 FILLCELL_X1 FILLER_106_1199 ();
 FILLCELL_X1 FILLER_106_1237 ();
 FILLCELL_X8 FILLER_106_1250 ();
 FILLCELL_X1 FILLER_106_1258 ();
 FILLCELL_X2 FILLER_106_1269 ();
 FILLCELL_X4 FILLER_106_1275 ();
 FILLCELL_X2 FILLER_106_1279 ();
 FILLCELL_X1 FILLER_106_1281 ();
 FILLCELL_X8 FILLER_106_1312 ();
 FILLCELL_X4 FILLER_106_1320 ();
 FILLCELL_X2 FILLER_106_1324 ();
 FILLCELL_X8 FILLER_106_1344 ();
 FILLCELL_X4 FILLER_106_1352 ();
 FILLCELL_X1 FILLER_106_1356 ();
 FILLCELL_X1 FILLER_106_1361 ();
 FILLCELL_X2 FILLER_106_1388 ();
 FILLCELL_X1 FILLER_106_1390 ();
 FILLCELL_X1 FILLER_106_1397 ();
 FILLCELL_X1 FILLER_106_1424 ();
 FILLCELL_X32 FILLER_106_1435 ();
 FILLCELL_X32 FILLER_106_1467 ();
 FILLCELL_X32 FILLER_106_1499 ();
 FILLCELL_X32 FILLER_106_1531 ();
 FILLCELL_X32 FILLER_106_1563 ();
 FILLCELL_X32 FILLER_106_1595 ();
 FILLCELL_X16 FILLER_106_1627 ();
 FILLCELL_X8 FILLER_106_1643 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X4 FILLER_107_33 ();
 FILLCELL_X1 FILLER_107_37 ();
 FILLCELL_X1 FILLER_107_58 ();
 FILLCELL_X4 FILLER_107_73 ();
 FILLCELL_X1 FILLER_107_77 ();
 FILLCELL_X8 FILLER_107_92 ();
 FILLCELL_X1 FILLER_107_100 ();
 FILLCELL_X2 FILLER_107_110 ();
 FILLCELL_X1 FILLER_107_112 ();
 FILLCELL_X2 FILLER_107_118 ();
 FILLCELL_X2 FILLER_107_134 ();
 FILLCELL_X4 FILLER_107_141 ();
 FILLCELL_X4 FILLER_107_154 ();
 FILLCELL_X4 FILLER_107_178 ();
 FILLCELL_X4 FILLER_107_202 ();
 FILLCELL_X2 FILLER_107_206 ();
 FILLCELL_X16 FILLER_107_248 ();
 FILLCELL_X1 FILLER_107_264 ();
 FILLCELL_X2 FILLER_107_281 ();
 FILLCELL_X8 FILLER_107_301 ();
 FILLCELL_X2 FILLER_107_309 ();
 FILLCELL_X4 FILLER_107_316 ();
 FILLCELL_X4 FILLER_107_347 ();
 FILLCELL_X1 FILLER_107_354 ();
 FILLCELL_X2 FILLER_107_386 ();
 FILLCELL_X8 FILLER_107_401 ();
 FILLCELL_X8 FILLER_107_442 ();
 FILLCELL_X1 FILLER_107_450 ();
 FILLCELL_X4 FILLER_107_454 ();
 FILLCELL_X1 FILLER_107_458 ();
 FILLCELL_X16 FILLER_107_468 ();
 FILLCELL_X2 FILLER_107_484 ();
 FILLCELL_X1 FILLER_107_497 ();
 FILLCELL_X2 FILLER_107_525 ();
 FILLCELL_X1 FILLER_107_527 ();
 FILLCELL_X2 FILLER_107_541 ();
 FILLCELL_X8 FILLER_107_568 ();
 FILLCELL_X2 FILLER_107_584 ();
 FILLCELL_X1 FILLER_107_586 ();
 FILLCELL_X2 FILLER_107_594 ();
 FILLCELL_X2 FILLER_107_618 ();
 FILLCELL_X2 FILLER_107_640 ();
 FILLCELL_X1 FILLER_107_642 ();
 FILLCELL_X16 FILLER_107_681 ();
 FILLCELL_X8 FILLER_107_697 ();
 FILLCELL_X2 FILLER_107_705 ();
 FILLCELL_X1 FILLER_107_707 ();
 FILLCELL_X4 FILLER_107_713 ();
 FILLCELL_X1 FILLER_107_747 ();
 FILLCELL_X2 FILLER_107_781 ();
 FILLCELL_X8 FILLER_107_796 ();
 FILLCELL_X2 FILLER_107_804 ();
 FILLCELL_X16 FILLER_107_830 ();
 FILLCELL_X4 FILLER_107_846 ();
 FILLCELL_X1 FILLER_107_850 ();
 FILLCELL_X4 FILLER_107_860 ();
 FILLCELL_X8 FILLER_107_876 ();
 FILLCELL_X4 FILLER_107_955 ();
 FILLCELL_X1 FILLER_107_959 ();
 FILLCELL_X1 FILLER_107_974 ();
 FILLCELL_X1 FILLER_107_982 ();
 FILLCELL_X1 FILLER_107_990 ();
 FILLCELL_X16 FILLER_107_998 ();
 FILLCELL_X8 FILLER_107_1020 ();
 FILLCELL_X1 FILLER_107_1028 ();
 FILLCELL_X8 FILLER_107_1055 ();
 FILLCELL_X2 FILLER_107_1087 ();
 FILLCELL_X1 FILLER_107_1089 ();
 FILLCELL_X1 FILLER_107_1096 ();
 FILLCELL_X4 FILLER_107_1103 ();
 FILLCELL_X1 FILLER_107_1107 ();
 FILLCELL_X1 FILLER_107_1120 ();
 FILLCELL_X4 FILLER_107_1141 ();
 FILLCELL_X1 FILLER_107_1145 ();
 FILLCELL_X8 FILLER_107_1150 ();
 FILLCELL_X4 FILLER_107_1158 ();
 FILLCELL_X2 FILLER_107_1162 ();
 FILLCELL_X4 FILLER_107_1180 ();
 FILLCELL_X2 FILLER_107_1184 ();
 FILLCELL_X8 FILLER_107_1207 ();
 FILLCELL_X2 FILLER_107_1215 ();
 FILLCELL_X2 FILLER_107_1245 ();
 FILLCELL_X4 FILLER_107_1258 ();
 FILLCELL_X1 FILLER_107_1262 ();
 FILLCELL_X4 FILLER_107_1264 ();
 FILLCELL_X2 FILLER_107_1268 ();
 FILLCELL_X4 FILLER_107_1296 ();
 FILLCELL_X2 FILLER_107_1300 ();
 FILLCELL_X1 FILLER_107_1302 ();
 FILLCELL_X1 FILLER_107_1305 ();
 FILLCELL_X1 FILLER_107_1330 ();
 FILLCELL_X1 FILLER_107_1337 ();
 FILLCELL_X1 FILLER_107_1360 ();
 FILLCELL_X1 FILLER_107_1368 ();
 FILLCELL_X1 FILLER_107_1373 ();
 FILLCELL_X16 FILLER_107_1377 ();
 FILLCELL_X32 FILLER_107_1422 ();
 FILLCELL_X32 FILLER_107_1454 ();
 FILLCELL_X32 FILLER_107_1486 ();
 FILLCELL_X32 FILLER_107_1518 ();
 FILLCELL_X32 FILLER_107_1550 ();
 FILLCELL_X32 FILLER_107_1582 ();
 FILLCELL_X32 FILLER_107_1614 ();
 FILLCELL_X4 FILLER_107_1646 ();
 FILLCELL_X1 FILLER_107_1650 ();
 FILLCELL_X16 FILLER_108_1 ();
 FILLCELL_X4 FILLER_108_17 ();
 FILLCELL_X1 FILLER_108_36 ();
 FILLCELL_X8 FILLER_108_64 ();
 FILLCELL_X4 FILLER_108_72 ();
 FILLCELL_X2 FILLER_108_76 ();
 FILLCELL_X1 FILLER_108_78 ();
 FILLCELL_X2 FILLER_108_119 ();
 FILLCELL_X1 FILLER_108_121 ();
 FILLCELL_X2 FILLER_108_145 ();
 FILLCELL_X2 FILLER_108_152 ();
 FILLCELL_X2 FILLER_108_161 ();
 FILLCELL_X1 FILLER_108_163 ();
 FILLCELL_X2 FILLER_108_171 ();
 FILLCELL_X2 FILLER_108_178 ();
 FILLCELL_X1 FILLER_108_180 ();
 FILLCELL_X2 FILLER_108_185 ();
 FILLCELL_X1 FILLER_108_187 ();
 FILLCELL_X2 FILLER_108_195 ();
 FILLCELL_X4 FILLER_108_209 ();
 FILLCELL_X2 FILLER_108_244 ();
 FILLCELL_X2 FILLER_108_250 ();
 FILLCELL_X1 FILLER_108_252 ();
 FILLCELL_X4 FILLER_108_273 ();
 FILLCELL_X2 FILLER_108_277 ();
 FILLCELL_X8 FILLER_108_308 ();
 FILLCELL_X8 FILLER_108_333 ();
 FILLCELL_X4 FILLER_108_364 ();
 FILLCELL_X2 FILLER_108_368 ();
 FILLCELL_X1 FILLER_108_370 ();
 FILLCELL_X1 FILLER_108_388 ();
 FILLCELL_X2 FILLER_108_398 ();
 FILLCELL_X1 FILLER_108_400 ();
 FILLCELL_X8 FILLER_108_410 ();
 FILLCELL_X1 FILLER_108_426 ();
 FILLCELL_X8 FILLER_108_499 ();
 FILLCELL_X4 FILLER_108_507 ();
 FILLCELL_X2 FILLER_108_511 ();
 FILLCELL_X1 FILLER_108_513 ();
 FILLCELL_X4 FILLER_108_516 ();
 FILLCELL_X16 FILLER_108_523 ();
 FILLCELL_X2 FILLER_108_552 ();
 FILLCELL_X1 FILLER_108_554 ();
 FILLCELL_X16 FILLER_108_575 ();
 FILLCELL_X8 FILLER_108_598 ();
 FILLCELL_X8 FILLER_108_613 ();
 FILLCELL_X1 FILLER_108_621 ();
 FILLCELL_X4 FILLER_108_626 ();
 FILLCELL_X1 FILLER_108_630 ();
 FILLCELL_X1 FILLER_108_632 ();
 FILLCELL_X1 FILLER_108_636 ();
 FILLCELL_X1 FILLER_108_650 ();
 FILLCELL_X2 FILLER_108_653 ();
 FILLCELL_X2 FILLER_108_659 ();
 FILLCELL_X4 FILLER_108_663 ();
 FILLCELL_X1 FILLER_108_670 ();
 FILLCELL_X4 FILLER_108_698 ();
 FILLCELL_X1 FILLER_108_702 ();
 FILLCELL_X4 FILLER_108_715 ();
 FILLCELL_X1 FILLER_108_732 ();
 FILLCELL_X2 FILLER_108_753 ();
 FILLCELL_X1 FILLER_108_759 ();
 FILLCELL_X2 FILLER_108_782 ();
 FILLCELL_X1 FILLER_108_784 ();
 FILLCELL_X2 FILLER_108_795 ();
 FILLCELL_X2 FILLER_108_806 ();
 FILLCELL_X4 FILLER_108_816 ();
 FILLCELL_X8 FILLER_108_824 ();
 FILLCELL_X1 FILLER_108_832 ();
 FILLCELL_X2 FILLER_108_850 ();
 FILLCELL_X1 FILLER_108_852 ();
 FILLCELL_X2 FILLER_108_866 ();
 FILLCELL_X1 FILLER_108_868 ();
 FILLCELL_X16 FILLER_108_891 ();
 FILLCELL_X4 FILLER_108_907 ();
 FILLCELL_X2 FILLER_108_911 ();
 FILLCELL_X1 FILLER_108_913 ();
 FILLCELL_X2 FILLER_108_943 ();
 FILLCELL_X8 FILLER_108_947 ();
 FILLCELL_X2 FILLER_108_955 ();
 FILLCELL_X4 FILLER_108_982 ();
 FILLCELL_X2 FILLER_108_986 ();
 FILLCELL_X1 FILLER_108_988 ();
 FILLCELL_X4 FILLER_108_1002 ();
 FILLCELL_X2 FILLER_108_1006 ();
 FILLCELL_X1 FILLER_108_1008 ();
 FILLCELL_X1 FILLER_108_1012 ();
 FILLCELL_X8 FILLER_108_1017 ();
 FILLCELL_X2 FILLER_108_1025 ();
 FILLCELL_X32 FILLER_108_1033 ();
 FILLCELL_X16 FILLER_108_1065 ();
 FILLCELL_X2 FILLER_108_1081 ();
 FILLCELL_X1 FILLER_108_1083 ();
 FILLCELL_X16 FILLER_108_1094 ();
 FILLCELL_X1 FILLER_108_1120 ();
 FILLCELL_X2 FILLER_108_1131 ();
 FILLCELL_X1 FILLER_108_1133 ();
 FILLCELL_X1 FILLER_108_1160 ();
 FILLCELL_X16 FILLER_108_1188 ();
 FILLCELL_X8 FILLER_108_1204 ();
 FILLCELL_X4 FILLER_108_1212 ();
 FILLCELL_X2 FILLER_108_1237 ();
 FILLCELL_X2 FILLER_108_1252 ();
 FILLCELL_X1 FILLER_108_1254 ();
 FILLCELL_X8 FILLER_108_1276 ();
 FILLCELL_X2 FILLER_108_1294 ();
 FILLCELL_X1 FILLER_108_1304 ();
 FILLCELL_X4 FILLER_108_1327 ();
 FILLCELL_X2 FILLER_108_1341 ();
 FILLCELL_X1 FILLER_108_1343 ();
 FILLCELL_X8 FILLER_108_1354 ();
 FILLCELL_X1 FILLER_108_1362 ();
 FILLCELL_X8 FILLER_108_1370 ();
 FILLCELL_X4 FILLER_108_1378 ();
 FILLCELL_X2 FILLER_108_1382 ();
 FILLCELL_X1 FILLER_108_1384 ();
 FILLCELL_X1 FILLER_108_1396 ();
 FILLCELL_X16 FILLER_108_1423 ();
 FILLCELL_X8 FILLER_108_1439 ();
 FILLCELL_X4 FILLER_108_1447 ();
 FILLCELL_X1 FILLER_108_1451 ();
 FILLCELL_X32 FILLER_108_1462 ();
 FILLCELL_X32 FILLER_108_1494 ();
 FILLCELL_X32 FILLER_108_1526 ();
 FILLCELL_X32 FILLER_108_1558 ();
 FILLCELL_X32 FILLER_108_1590 ();
 FILLCELL_X16 FILLER_108_1622 ();
 FILLCELL_X8 FILLER_108_1638 ();
 FILLCELL_X4 FILLER_108_1646 ();
 FILLCELL_X1 FILLER_108_1650 ();
 FILLCELL_X16 FILLER_109_1 ();
 FILLCELL_X4 FILLER_109_17 ();
 FILLCELL_X1 FILLER_109_21 ();
 FILLCELL_X1 FILLER_109_97 ();
 FILLCELL_X1 FILLER_109_103 ();
 FILLCELL_X2 FILLER_109_117 ();
 FILLCELL_X4 FILLER_109_128 ();
 FILLCELL_X2 FILLER_109_132 ();
 FILLCELL_X4 FILLER_109_186 ();
 FILLCELL_X2 FILLER_109_214 ();
 FILLCELL_X1 FILLER_109_216 ();
 FILLCELL_X2 FILLER_109_267 ();
 FILLCELL_X2 FILLER_109_298 ();
 FILLCELL_X8 FILLER_109_337 ();
 FILLCELL_X4 FILLER_109_345 ();
 FILLCELL_X2 FILLER_109_349 ();
 FILLCELL_X1 FILLER_109_354 ();
 FILLCELL_X8 FILLER_109_368 ();
 FILLCELL_X4 FILLER_109_376 ();
 FILLCELL_X2 FILLER_109_380 ();
 FILLCELL_X4 FILLER_109_386 ();
 FILLCELL_X2 FILLER_109_390 ();
 FILLCELL_X1 FILLER_109_392 ();
 FILLCELL_X2 FILLER_109_395 ();
 FILLCELL_X8 FILLER_109_432 ();
 FILLCELL_X8 FILLER_109_455 ();
 FILLCELL_X4 FILLER_109_463 ();
 FILLCELL_X2 FILLER_109_467 ();
 FILLCELL_X1 FILLER_109_489 ();
 FILLCELL_X2 FILLER_109_519 ();
 FILLCELL_X4 FILLER_109_534 ();
 FILLCELL_X2 FILLER_109_571 ();
 FILLCELL_X1 FILLER_109_573 ();
 FILLCELL_X2 FILLER_109_597 ();
 FILLCELL_X8 FILLER_109_624 ();
 FILLCELL_X2 FILLER_109_632 ();
 FILLCELL_X1 FILLER_109_634 ();
 FILLCELL_X16 FILLER_109_680 ();
 FILLCELL_X2 FILLER_109_705 ();
 FILLCELL_X4 FILLER_109_734 ();
 FILLCELL_X2 FILLER_109_738 ();
 FILLCELL_X1 FILLER_109_740 ();
 FILLCELL_X8 FILLER_109_748 ();
 FILLCELL_X2 FILLER_109_756 ();
 FILLCELL_X1 FILLER_109_758 ();
 FILLCELL_X1 FILLER_109_762 ();
 FILLCELL_X8 FILLER_109_779 ();
 FILLCELL_X4 FILLER_109_787 ();
 FILLCELL_X1 FILLER_109_791 ();
 FILLCELL_X2 FILLER_109_812 ();
 FILLCELL_X4 FILLER_109_819 ();
 FILLCELL_X2 FILLER_109_823 ();
 FILLCELL_X2 FILLER_109_828 ();
 FILLCELL_X2 FILLER_109_840 ();
 FILLCELL_X1 FILLER_109_842 ();
 FILLCELL_X4 FILLER_109_871 ();
 FILLCELL_X16 FILLER_109_888 ();
 FILLCELL_X2 FILLER_109_904 ();
 FILLCELL_X1 FILLER_109_913 ();
 FILLCELL_X4 FILLER_109_921 ();
 FILLCELL_X2 FILLER_109_925 ();
 FILLCELL_X4 FILLER_109_932 ();
 FILLCELL_X4 FILLER_109_977 ();
 FILLCELL_X4 FILLER_109_983 ();
 FILLCELL_X2 FILLER_109_987 ();
 FILLCELL_X16 FILLER_109_992 ();
 FILLCELL_X1 FILLER_109_1008 ();
 FILLCELL_X1 FILLER_109_1023 ();
 FILLCELL_X8 FILLER_109_1031 ();
 FILLCELL_X4 FILLER_109_1039 ();
 FILLCELL_X4 FILLER_109_1059 ();
 FILLCELL_X1 FILLER_109_1065 ();
 FILLCELL_X1 FILLER_109_1075 ();
 FILLCELL_X2 FILLER_109_1079 ();
 FILLCELL_X1 FILLER_109_1081 ();
 FILLCELL_X1 FILLER_109_1085 ();
 FILLCELL_X16 FILLER_109_1092 ();
 FILLCELL_X4 FILLER_109_1108 ();
 FILLCELL_X1 FILLER_109_1112 ();
 FILLCELL_X4 FILLER_109_1130 ();
 FILLCELL_X1 FILLER_109_1149 ();
 FILLCELL_X8 FILLER_109_1153 ();
 FILLCELL_X4 FILLER_109_1161 ();
 FILLCELL_X1 FILLER_109_1165 ();
 FILLCELL_X2 FILLER_109_1182 ();
 FILLCELL_X1 FILLER_109_1184 ();
 FILLCELL_X1 FILLER_109_1214 ();
 FILLCELL_X1 FILLER_109_1219 ();
 FILLCELL_X2 FILLER_109_1227 ();
 FILLCELL_X2 FILLER_109_1232 ();
 FILLCELL_X2 FILLER_109_1244 ();
 FILLCELL_X4 FILLER_109_1309 ();
 FILLCELL_X2 FILLER_109_1313 ();
 FILLCELL_X1 FILLER_109_1315 ();
 FILLCELL_X2 FILLER_109_1321 ();
 FILLCELL_X2 FILLER_109_1329 ();
 FILLCELL_X1 FILLER_109_1331 ();
 FILLCELL_X1 FILLER_109_1341 ();
 FILLCELL_X2 FILLER_109_1348 ();
 FILLCELL_X1 FILLER_109_1350 ();
 FILLCELL_X1 FILLER_109_1358 ();
 FILLCELL_X1 FILLER_109_1363 ();
 FILLCELL_X16 FILLER_109_1403 ();
 FILLCELL_X4 FILLER_109_1431 ();
 FILLCELL_X32 FILLER_109_1473 ();
 FILLCELL_X32 FILLER_109_1505 ();
 FILLCELL_X32 FILLER_109_1537 ();
 FILLCELL_X32 FILLER_109_1569 ();
 FILLCELL_X32 FILLER_109_1601 ();
 FILLCELL_X16 FILLER_109_1633 ();
 FILLCELL_X2 FILLER_109_1649 ();
 FILLCELL_X8 FILLER_110_1 ();
 FILLCELL_X4 FILLER_110_9 ();
 FILLCELL_X2 FILLER_110_13 ();
 FILLCELL_X1 FILLER_110_15 ();
 FILLCELL_X4 FILLER_110_73 ();
 FILLCELL_X2 FILLER_110_77 ();
 FILLCELL_X1 FILLER_110_79 ();
 FILLCELL_X4 FILLER_110_87 ();
 FILLCELL_X2 FILLER_110_91 ();
 FILLCELL_X1 FILLER_110_93 ();
 FILLCELL_X4 FILLER_110_101 ();
 FILLCELL_X1 FILLER_110_105 ();
 FILLCELL_X4 FILLER_110_126 ();
 FILLCELL_X2 FILLER_110_130 ();
 FILLCELL_X2 FILLER_110_159 ();
 FILLCELL_X1 FILLER_110_161 ();
 FILLCELL_X8 FILLER_110_171 ();
 FILLCELL_X4 FILLER_110_179 ();
 FILLCELL_X1 FILLER_110_183 ();
 FILLCELL_X2 FILLER_110_204 ();
 FILLCELL_X8 FILLER_110_226 ();
 FILLCELL_X4 FILLER_110_234 ();
 FILLCELL_X8 FILLER_110_241 ();
 FILLCELL_X8 FILLER_110_252 ();
 FILLCELL_X2 FILLER_110_260 ();
 FILLCELL_X1 FILLER_110_262 ();
 FILLCELL_X4 FILLER_110_268 ();
 FILLCELL_X1 FILLER_110_272 ();
 FILLCELL_X4 FILLER_110_300 ();
 FILLCELL_X2 FILLER_110_327 ();
 FILLCELL_X1 FILLER_110_342 ();
 FILLCELL_X1 FILLER_110_350 ();
 FILLCELL_X1 FILLER_110_364 ();
 FILLCELL_X8 FILLER_110_372 ();
 FILLCELL_X4 FILLER_110_402 ();
 FILLCELL_X2 FILLER_110_410 ();
 FILLCELL_X2 FILLER_110_432 ();
 FILLCELL_X1 FILLER_110_434 ();
 FILLCELL_X8 FILLER_110_442 ();
 FILLCELL_X4 FILLER_110_450 ();
 FILLCELL_X1 FILLER_110_454 ();
 FILLCELL_X4 FILLER_110_462 ();
 FILLCELL_X2 FILLER_110_466 ();
 FILLCELL_X1 FILLER_110_472 ();
 FILLCELL_X1 FILLER_110_479 ();
 FILLCELL_X2 FILLER_110_484 ();
 FILLCELL_X2 FILLER_110_496 ();
 FILLCELL_X8 FILLER_110_535 ();
 FILLCELL_X1 FILLER_110_543 ();
 FILLCELL_X16 FILLER_110_550 ();
 FILLCELL_X8 FILLER_110_566 ();
 FILLCELL_X4 FILLER_110_601 ();
 FILLCELL_X1 FILLER_110_605 ();
 FILLCELL_X4 FILLER_110_619 ();
 FILLCELL_X2 FILLER_110_623 ();
 FILLCELL_X1 FILLER_110_625 ();
 FILLCELL_X4 FILLER_110_632 ();
 FILLCELL_X8 FILLER_110_656 ();
 FILLCELL_X4 FILLER_110_664 ();
 FILLCELL_X16 FILLER_110_681 ();
 FILLCELL_X2 FILLER_110_697 ();
 FILLCELL_X4 FILLER_110_719 ();
 FILLCELL_X1 FILLER_110_727 ();
 FILLCELL_X8 FILLER_110_736 ();
 FILLCELL_X1 FILLER_110_744 ();
 FILLCELL_X2 FILLER_110_776 ();
 FILLCELL_X8 FILLER_110_791 ();
 FILLCELL_X2 FILLER_110_799 ();
 FILLCELL_X1 FILLER_110_801 ();
 FILLCELL_X8 FILLER_110_819 ();
 FILLCELL_X4 FILLER_110_827 ();
 FILLCELL_X1 FILLER_110_831 ();
 FILLCELL_X2 FILLER_110_839 ();
 FILLCELL_X8 FILLER_110_854 ();
 FILLCELL_X2 FILLER_110_862 ();
 FILLCELL_X1 FILLER_110_864 ();
 FILLCELL_X1 FILLER_110_887 ();
 FILLCELL_X16 FILLER_110_937 ();
 FILLCELL_X8 FILLER_110_953 ();
 FILLCELL_X4 FILLER_110_961 ();
 FILLCELL_X2 FILLER_110_965 ();
 FILLCELL_X1 FILLER_110_967 ();
 FILLCELL_X2 FILLER_110_982 ();
 FILLCELL_X1 FILLER_110_984 ();
 FILLCELL_X1 FILLER_110_989 ();
 FILLCELL_X16 FILLER_110_997 ();
 FILLCELL_X8 FILLER_110_1013 ();
 FILLCELL_X4 FILLER_110_1021 ();
 FILLCELL_X1 FILLER_110_1025 ();
 FILLCELL_X1 FILLER_110_1054 ();
 FILLCELL_X2 FILLER_110_1060 ();
 FILLCELL_X2 FILLER_110_1069 ();
 FILLCELL_X1 FILLER_110_1071 ();
 FILLCELL_X1 FILLER_110_1078 ();
 FILLCELL_X8 FILLER_110_1084 ();
 FILLCELL_X4 FILLER_110_1092 ();
 FILLCELL_X1 FILLER_110_1096 ();
 FILLCELL_X8 FILLER_110_1107 ();
 FILLCELL_X2 FILLER_110_1115 ();
 FILLCELL_X8 FILLER_110_1127 ();
 FILLCELL_X4 FILLER_110_1135 ();
 FILLCELL_X8 FILLER_110_1144 ();
 FILLCELL_X1 FILLER_110_1152 ();
 FILLCELL_X8 FILLER_110_1160 ();
 FILLCELL_X2 FILLER_110_1168 ();
 FILLCELL_X1 FILLER_110_1170 ();
 FILLCELL_X2 FILLER_110_1174 ();
 FILLCELL_X1 FILLER_110_1186 ();
 FILLCELL_X8 FILLER_110_1202 ();
 FILLCELL_X1 FILLER_110_1239 ();
 FILLCELL_X4 FILLER_110_1247 ();
 FILLCELL_X2 FILLER_110_1263 ();
 FILLCELL_X8 FILLER_110_1272 ();
 FILLCELL_X4 FILLER_110_1280 ();
 FILLCELL_X1 FILLER_110_1315 ();
 FILLCELL_X2 FILLER_110_1342 ();
 FILLCELL_X2 FILLER_110_1348 ();
 FILLCELL_X2 FILLER_110_1372 ();
 FILLCELL_X1 FILLER_110_1374 ();
 FILLCELL_X4 FILLER_110_1379 ();
 FILLCELL_X1 FILLER_110_1389 ();
 FILLCELL_X4 FILLER_110_1402 ();
 FILLCELL_X2 FILLER_110_1406 ();
 FILLCELL_X1 FILLER_110_1408 ();
 FILLCELL_X2 FILLER_110_1419 ();
 FILLCELL_X2 FILLER_110_1427 ();
 FILLCELL_X2 FILLER_110_1439 ();
 FILLCELL_X1 FILLER_110_1441 ();
 FILLCELL_X4 FILLER_110_1448 ();
 FILLCELL_X2 FILLER_110_1452 ();
 FILLCELL_X32 FILLER_110_1472 ();
 FILLCELL_X32 FILLER_110_1504 ();
 FILLCELL_X32 FILLER_110_1536 ();
 FILLCELL_X32 FILLER_110_1568 ();
 FILLCELL_X32 FILLER_110_1600 ();
 FILLCELL_X16 FILLER_110_1632 ();
 FILLCELL_X2 FILLER_110_1648 ();
 FILLCELL_X1 FILLER_110_1650 ();
 FILLCELL_X16 FILLER_111_1 ();
 FILLCELL_X1 FILLER_111_17 ();
 FILLCELL_X4 FILLER_111_66 ();
 FILLCELL_X1 FILLER_111_70 ();
 FILLCELL_X4 FILLER_111_80 ();
 FILLCELL_X2 FILLER_111_84 ();
 FILLCELL_X4 FILLER_111_149 ();
 FILLCELL_X2 FILLER_111_153 ();
 FILLCELL_X16 FILLER_111_160 ();
 FILLCELL_X4 FILLER_111_176 ();
 FILLCELL_X1 FILLER_111_180 ();
 FILLCELL_X1 FILLER_111_207 ();
 FILLCELL_X4 FILLER_111_215 ();
 FILLCELL_X2 FILLER_111_219 ();
 FILLCELL_X1 FILLER_111_221 ();
 FILLCELL_X4 FILLER_111_229 ();
 FILLCELL_X2 FILLER_111_233 ();
 FILLCELL_X8 FILLER_111_249 ();
 FILLCELL_X2 FILLER_111_257 ();
 FILLCELL_X1 FILLER_111_259 ();
 FILLCELL_X4 FILLER_111_264 ();
 FILLCELL_X2 FILLER_111_268 ();
 FILLCELL_X1 FILLER_111_270 ();
 FILLCELL_X8 FILLER_111_300 ();
 FILLCELL_X4 FILLER_111_328 ();
 FILLCELL_X2 FILLER_111_332 ();
 FILLCELL_X2 FILLER_111_354 ();
 FILLCELL_X16 FILLER_111_396 ();
 FILLCELL_X4 FILLER_111_412 ();
 FILLCELL_X2 FILLER_111_416 ();
 FILLCELL_X8 FILLER_111_431 ();
 FILLCELL_X2 FILLER_111_439 ();
 FILLCELL_X2 FILLER_111_448 ();
 FILLCELL_X1 FILLER_111_450 ();
 FILLCELL_X2 FILLER_111_458 ();
 FILLCELL_X1 FILLER_111_460 ();
 FILLCELL_X1 FILLER_111_481 ();
 FILLCELL_X8 FILLER_111_502 ();
 FILLCELL_X2 FILLER_111_510 ();
 FILLCELL_X4 FILLER_111_516 ();
 FILLCELL_X2 FILLER_111_520 ();
 FILLCELL_X1 FILLER_111_522 ();
 FILLCELL_X1 FILLER_111_526 ();
 FILLCELL_X2 FILLER_111_536 ();
 FILLCELL_X1 FILLER_111_538 ();
 FILLCELL_X8 FILLER_111_559 ();
 FILLCELL_X4 FILLER_111_567 ();
 FILLCELL_X2 FILLER_111_571 ();
 FILLCELL_X1 FILLER_111_573 ();
 FILLCELL_X1 FILLER_111_578 ();
 FILLCELL_X1 FILLER_111_596 ();
 FILLCELL_X1 FILLER_111_617 ();
 FILLCELL_X2 FILLER_111_647 ();
 FILLCELL_X1 FILLER_111_649 ();
 FILLCELL_X16 FILLER_111_654 ();
 FILLCELL_X1 FILLER_111_670 ();
 FILLCELL_X4 FILLER_111_678 ();
 FILLCELL_X4 FILLER_111_686 ();
 FILLCELL_X2 FILLER_111_720 ();
 FILLCELL_X4 FILLER_111_753 ();
 FILLCELL_X1 FILLER_111_757 ();
 FILLCELL_X1 FILLER_111_771 ();
 FILLCELL_X2 FILLER_111_799 ();
 FILLCELL_X1 FILLER_111_801 ();
 FILLCELL_X8 FILLER_111_824 ();
 FILLCELL_X4 FILLER_111_832 ();
 FILLCELL_X1 FILLER_111_836 ();
 FILLCELL_X4 FILLER_111_857 ();
 FILLCELL_X1 FILLER_111_861 ();
 FILLCELL_X4 FILLER_111_869 ();
 FILLCELL_X8 FILLER_111_880 ();
 FILLCELL_X2 FILLER_111_888 ();
 FILLCELL_X2 FILLER_111_926 ();
 FILLCELL_X4 FILLER_111_935 ();
 FILLCELL_X8 FILLER_111_959 ();
 FILLCELL_X2 FILLER_111_967 ();
 FILLCELL_X1 FILLER_111_969 ();
 FILLCELL_X4 FILLER_111_990 ();
 FILLCELL_X1 FILLER_111_994 ();
 FILLCELL_X1 FILLER_111_1007 ();
 FILLCELL_X1 FILLER_111_1017 ();
 FILLCELL_X8 FILLER_111_1028 ();
 FILLCELL_X4 FILLER_111_1036 ();
 FILLCELL_X2 FILLER_111_1040 ();
 FILLCELL_X4 FILLER_111_1050 ();
 FILLCELL_X1 FILLER_111_1054 ();
 FILLCELL_X8 FILLER_111_1060 ();
 FILLCELL_X4 FILLER_111_1068 ();
 FILLCELL_X2 FILLER_111_1072 ();
 FILLCELL_X1 FILLER_111_1074 ();
 FILLCELL_X8 FILLER_111_1082 ();
 FILLCELL_X2 FILLER_111_1090 ();
 FILLCELL_X8 FILLER_111_1098 ();
 FILLCELL_X4 FILLER_111_1106 ();
 FILLCELL_X2 FILLER_111_1110 ();
 FILLCELL_X8 FILLER_111_1135 ();
 FILLCELL_X1 FILLER_111_1143 ();
 FILLCELL_X4 FILLER_111_1149 ();
 FILLCELL_X8 FILLER_111_1160 ();
 FILLCELL_X16 FILLER_111_1204 ();
 FILLCELL_X8 FILLER_111_1220 ();
 FILLCELL_X2 FILLER_111_1232 ();
 FILLCELL_X4 FILLER_111_1256 ();
 FILLCELL_X2 FILLER_111_1260 ();
 FILLCELL_X1 FILLER_111_1262 ();
 FILLCELL_X8 FILLER_111_1284 ();
 FILLCELL_X8 FILLER_111_1294 ();
 FILLCELL_X2 FILLER_111_1302 ();
 FILLCELL_X1 FILLER_111_1304 ();
 FILLCELL_X4 FILLER_111_1315 ();
 FILLCELL_X2 FILLER_111_1319 ();
 FILLCELL_X1 FILLER_111_1321 ();
 FILLCELL_X16 FILLER_111_1326 ();
 FILLCELL_X8 FILLER_111_1342 ();
 FILLCELL_X4 FILLER_111_1350 ();
 FILLCELL_X1 FILLER_111_1354 ();
 FILLCELL_X16 FILLER_111_1377 ();
 FILLCELL_X2 FILLER_111_1393 ();
 FILLCELL_X1 FILLER_111_1405 ();
 FILLCELL_X1 FILLER_111_1416 ();
 FILLCELL_X1 FILLER_111_1423 ();
 FILLCELL_X1 FILLER_111_1434 ();
 FILLCELL_X1 FILLER_111_1441 ();
 FILLCELL_X8 FILLER_111_1452 ();
 FILLCELL_X4 FILLER_111_1460 ();
 FILLCELL_X1 FILLER_111_1464 ();
 FILLCELL_X32 FILLER_111_1471 ();
 FILLCELL_X32 FILLER_111_1503 ();
 FILLCELL_X32 FILLER_111_1535 ();
 FILLCELL_X32 FILLER_111_1567 ();
 FILLCELL_X32 FILLER_111_1599 ();
 FILLCELL_X16 FILLER_111_1631 ();
 FILLCELL_X4 FILLER_111_1647 ();
 FILLCELL_X16 FILLER_112_1 ();
 FILLCELL_X8 FILLER_112_17 ();
 FILLCELL_X4 FILLER_112_25 ();
 FILLCELL_X2 FILLER_112_36 ();
 FILLCELL_X1 FILLER_112_38 ();
 FILLCELL_X8 FILLER_112_44 ();
 FILLCELL_X2 FILLER_112_52 ();
 FILLCELL_X1 FILLER_112_54 ();
 FILLCELL_X1 FILLER_112_75 ();
 FILLCELL_X4 FILLER_112_83 ();
 FILLCELL_X2 FILLER_112_87 ();
 FILLCELL_X1 FILLER_112_109 ();
 FILLCELL_X2 FILLER_112_115 ();
 FILLCELL_X2 FILLER_112_130 ();
 FILLCELL_X1 FILLER_112_132 ();
 FILLCELL_X1 FILLER_112_153 ();
 FILLCELL_X2 FILLER_112_161 ();
 FILLCELL_X1 FILLER_112_163 ();
 FILLCELL_X4 FILLER_112_191 ();
 FILLCELL_X8 FILLER_112_202 ();
 FILLCELL_X4 FILLER_112_210 ();
 FILLCELL_X1 FILLER_112_214 ();
 FILLCELL_X2 FILLER_112_235 ();
 FILLCELL_X1 FILLER_112_237 ();
 FILLCELL_X4 FILLER_112_242 ();
 FILLCELL_X1 FILLER_112_246 ();
 FILLCELL_X2 FILLER_112_254 ();
 FILLCELL_X4 FILLER_112_276 ();
 FILLCELL_X1 FILLER_112_280 ();
 FILLCELL_X16 FILLER_112_291 ();
 FILLCELL_X4 FILLER_112_307 ();
 FILLCELL_X8 FILLER_112_318 ();
 FILLCELL_X8 FILLER_112_333 ();
 FILLCELL_X4 FILLER_112_341 ();
 FILLCELL_X1 FILLER_112_345 ();
 FILLCELL_X2 FILLER_112_349 ();
 FILLCELL_X4 FILLER_112_364 ();
 FILLCELL_X4 FILLER_112_412 ();
 FILLCELL_X1 FILLER_112_416 ();
 FILLCELL_X4 FILLER_112_461 ();
 FILLCELL_X2 FILLER_112_465 ();
 FILLCELL_X1 FILLER_112_467 ();
 FILLCELL_X2 FILLER_112_510 ();
 FILLCELL_X1 FILLER_112_512 ();
 FILLCELL_X4 FILLER_112_516 ();
 FILLCELL_X2 FILLER_112_520 ();
 FILLCELL_X1 FILLER_112_522 ();
 FILLCELL_X2 FILLER_112_556 ();
 FILLCELL_X1 FILLER_112_558 ();
 FILLCELL_X4 FILLER_112_563 ();
 FILLCELL_X2 FILLER_112_596 ();
 FILLCELL_X8 FILLER_112_605 ();
 FILLCELL_X1 FILLER_112_613 ();
 FILLCELL_X4 FILLER_112_632 ();
 FILLCELL_X2 FILLER_112_640 ();
 FILLCELL_X2 FILLER_112_662 ();
 FILLCELL_X1 FILLER_112_664 ();
 FILLCELL_X2 FILLER_112_685 ();
 FILLCELL_X1 FILLER_112_687 ();
 FILLCELL_X4 FILLER_112_695 ();
 FILLCELL_X1 FILLER_112_699 ();
 FILLCELL_X2 FILLER_112_731 ();
 FILLCELL_X1 FILLER_112_733 ();
 FILLCELL_X2 FILLER_112_737 ();
 FILLCELL_X1 FILLER_112_739 ();
 FILLCELL_X2 FILLER_112_760 ();
 FILLCELL_X1 FILLER_112_762 ();
 FILLCELL_X2 FILLER_112_783 ();
 FILLCELL_X8 FILLER_112_825 ();
 FILLCELL_X4 FILLER_112_833 ();
 FILLCELL_X8 FILLER_112_842 ();
 FILLCELL_X2 FILLER_112_850 ();
 FILLCELL_X1 FILLER_112_852 ();
 FILLCELL_X2 FILLER_112_869 ();
 FILLCELL_X1 FILLER_112_871 ();
 FILLCELL_X16 FILLER_112_894 ();
 FILLCELL_X8 FILLER_112_910 ();
 FILLCELL_X4 FILLER_112_918 ();
 FILLCELL_X16 FILLER_112_944 ();
 FILLCELL_X8 FILLER_112_960 ();
 FILLCELL_X4 FILLER_112_968 ();
 FILLCELL_X1 FILLER_112_972 ();
 FILLCELL_X8 FILLER_112_994 ();
 FILLCELL_X1 FILLER_112_1002 ();
 FILLCELL_X4 FILLER_112_1010 ();
 FILLCELL_X1 FILLER_112_1014 ();
 FILLCELL_X8 FILLER_112_1028 ();
 FILLCELL_X4 FILLER_112_1036 ();
 FILLCELL_X32 FILLER_112_1063 ();
 FILLCELL_X8 FILLER_112_1095 ();
 FILLCELL_X4 FILLER_112_1103 ();
 FILLCELL_X1 FILLER_112_1107 ();
 FILLCELL_X4 FILLER_112_1124 ();
 FILLCELL_X1 FILLER_112_1128 ();
 FILLCELL_X4 FILLER_112_1136 ();
 FILLCELL_X4 FILLER_112_1192 ();
 FILLCELL_X8 FILLER_112_1218 ();
 FILLCELL_X2 FILLER_112_1226 ();
 FILLCELL_X2 FILLER_112_1235 ();
 FILLCELL_X1 FILLER_112_1237 ();
 FILLCELL_X4 FILLER_112_1243 ();
 FILLCELL_X4 FILLER_112_1257 ();
 FILLCELL_X2 FILLER_112_1261 ();
 FILLCELL_X2 FILLER_112_1285 ();
 FILLCELL_X4 FILLER_112_1344 ();
 FILLCELL_X4 FILLER_112_1362 ();
 FILLCELL_X2 FILLER_112_1366 ();
 FILLCELL_X1 FILLER_112_1368 ();
 FILLCELL_X8 FILLER_112_1375 ();
 FILLCELL_X4 FILLER_112_1383 ();
 FILLCELL_X4 FILLER_112_1399 ();
 FILLCELL_X8 FILLER_112_1413 ();
 FILLCELL_X1 FILLER_112_1421 ();
 FILLCELL_X2 FILLER_112_1437 ();
 FILLCELL_X1 FILLER_112_1449 ();
 FILLCELL_X4 FILLER_112_1460 ();
 FILLCELL_X2 FILLER_112_1464 ();
 FILLCELL_X2 FILLER_112_1472 ();
 FILLCELL_X32 FILLER_112_1484 ();
 FILLCELL_X32 FILLER_112_1516 ();
 FILLCELL_X32 FILLER_112_1548 ();
 FILLCELL_X32 FILLER_112_1580 ();
 FILLCELL_X32 FILLER_112_1612 ();
 FILLCELL_X4 FILLER_112_1644 ();
 FILLCELL_X2 FILLER_112_1648 ();
 FILLCELL_X1 FILLER_112_1650 ();
 FILLCELL_X8 FILLER_113_1 ();
 FILLCELL_X2 FILLER_113_9 ();
 FILLCELL_X1 FILLER_113_11 ();
 FILLCELL_X1 FILLER_113_32 ();
 FILLCELL_X2 FILLER_113_63 ();
 FILLCELL_X1 FILLER_113_65 ();
 FILLCELL_X4 FILLER_113_113 ();
 FILLCELL_X1 FILLER_113_117 ();
 FILLCELL_X4 FILLER_113_154 ();
 FILLCELL_X2 FILLER_113_158 ();
 FILLCELL_X4 FILLER_113_178 ();
 FILLCELL_X2 FILLER_113_182 ();
 FILLCELL_X1 FILLER_113_184 ();
 FILLCELL_X1 FILLER_113_190 ();
 FILLCELL_X1 FILLER_113_211 ();
 FILLCELL_X1 FILLER_113_232 ();
 FILLCELL_X1 FILLER_113_253 ();
 FILLCELL_X2 FILLER_113_259 ();
 FILLCELL_X4 FILLER_113_263 ();
 FILLCELL_X1 FILLER_113_267 ();
 FILLCELL_X2 FILLER_113_288 ();
 FILLCELL_X1 FILLER_113_290 ();
 FILLCELL_X4 FILLER_113_318 ();
 FILLCELL_X2 FILLER_113_322 ();
 FILLCELL_X16 FILLER_113_344 ();
 FILLCELL_X8 FILLER_113_360 ();
 FILLCELL_X4 FILLER_113_368 ();
 FILLCELL_X2 FILLER_113_392 ();
 FILLCELL_X4 FILLER_113_410 ();
 FILLCELL_X1 FILLER_113_414 ();
 FILLCELL_X2 FILLER_113_441 ();
 FILLCELL_X1 FILLER_113_443 ();
 FILLCELL_X2 FILLER_113_469 ();
 FILLCELL_X1 FILLER_113_478 ();
 FILLCELL_X8 FILLER_113_484 ();
 FILLCELL_X4 FILLER_113_492 ();
 FILLCELL_X1 FILLER_113_551 ();
 FILLCELL_X2 FILLER_113_561 ();
 FILLCELL_X1 FILLER_113_563 ();
 FILLCELL_X2 FILLER_113_589 ();
 FILLCELL_X1 FILLER_113_591 ();
 FILLCELL_X4 FILLER_113_615 ();
 FILLCELL_X1 FILLER_113_619 ();
 FILLCELL_X8 FILLER_113_647 ();
 FILLCELL_X4 FILLER_113_655 ();
 FILLCELL_X1 FILLER_113_659 ();
 FILLCELL_X4 FILLER_113_676 ();
 FILLCELL_X1 FILLER_113_680 ();
 FILLCELL_X4 FILLER_113_727 ();
 FILLCELL_X2 FILLER_113_735 ();
 FILLCELL_X8 FILLER_113_758 ();
 FILLCELL_X4 FILLER_113_766 ();
 FILLCELL_X2 FILLER_113_770 ();
 FILLCELL_X1 FILLER_113_788 ();
 FILLCELL_X8 FILLER_113_796 ();
 FILLCELL_X1 FILLER_113_804 ();
 FILLCELL_X4 FILLER_113_812 ();
 FILLCELL_X1 FILLER_113_816 ();
 FILLCELL_X4 FILLER_113_870 ();
 FILLCELL_X2 FILLER_113_874 ();
 FILLCELL_X16 FILLER_113_889 ();
 FILLCELL_X8 FILLER_113_919 ();
 FILLCELL_X2 FILLER_113_927 ();
 FILLCELL_X1 FILLER_113_929 ();
 FILLCELL_X16 FILLER_113_944 ();
 FILLCELL_X4 FILLER_113_960 ();
 FILLCELL_X8 FILLER_113_978 ();
 FILLCELL_X4 FILLER_113_986 ();
 FILLCELL_X2 FILLER_113_1000 ();
 FILLCELL_X4 FILLER_113_1011 ();
 FILLCELL_X16 FILLER_113_1022 ();
 FILLCELL_X1 FILLER_113_1038 ();
 FILLCELL_X2 FILLER_113_1045 ();
 FILLCELL_X4 FILLER_113_1068 ();
 FILLCELL_X1 FILLER_113_1101 ();
 FILLCELL_X1 FILLER_113_1124 ();
 FILLCELL_X16 FILLER_113_1147 ();
 FILLCELL_X2 FILLER_113_1163 ();
 FILLCELL_X4 FILLER_113_1190 ();
 FILLCELL_X1 FILLER_113_1194 ();
 FILLCELL_X1 FILLER_113_1206 ();
 FILLCELL_X2 FILLER_113_1229 ();
 FILLCELL_X2 FILLER_113_1261 ();
 FILLCELL_X2 FILLER_113_1264 ();
 FILLCELL_X4 FILLER_113_1275 ();
 FILLCELL_X2 FILLER_113_1279 ();
 FILLCELL_X1 FILLER_113_1301 ();
 FILLCELL_X1 FILLER_113_1312 ();
 FILLCELL_X2 FILLER_113_1323 ();
 FILLCELL_X1 FILLER_113_1328 ();
 FILLCELL_X2 FILLER_113_1338 ();
 FILLCELL_X16 FILLER_113_1350 ();
 FILLCELL_X8 FILLER_113_1366 ();
 FILLCELL_X4 FILLER_113_1374 ();
 FILLCELL_X2 FILLER_113_1378 ();
 FILLCELL_X16 FILLER_113_1404 ();
 FILLCELL_X1 FILLER_113_1420 ();
 FILLCELL_X4 FILLER_113_1439 ();
 FILLCELL_X2 FILLER_113_1480 ();
 FILLCELL_X32 FILLER_113_1492 ();
 FILLCELL_X32 FILLER_113_1524 ();
 FILLCELL_X32 FILLER_113_1556 ();
 FILLCELL_X32 FILLER_113_1588 ();
 FILLCELL_X16 FILLER_113_1620 ();
 FILLCELL_X8 FILLER_113_1636 ();
 FILLCELL_X4 FILLER_113_1644 ();
 FILLCELL_X2 FILLER_113_1648 ();
 FILLCELL_X1 FILLER_113_1650 ();
 FILLCELL_X8 FILLER_114_28 ();
 FILLCELL_X2 FILLER_114_36 ();
 FILLCELL_X1 FILLER_114_38 ();
 FILLCELL_X16 FILLER_114_82 ();
 FILLCELL_X2 FILLER_114_98 ();
 FILLCELL_X1 FILLER_114_100 ();
 FILLCELL_X8 FILLER_114_160 ();
 FILLCELL_X4 FILLER_114_168 ();
 FILLCELL_X1 FILLER_114_172 ();
 FILLCELL_X4 FILLER_114_193 ();
 FILLCELL_X4 FILLER_114_202 ();
 FILLCELL_X1 FILLER_114_206 ();
 FILLCELL_X2 FILLER_114_222 ();
 FILLCELL_X1 FILLER_114_231 ();
 FILLCELL_X8 FILLER_114_237 ();
 FILLCELL_X1 FILLER_114_245 ();
 FILLCELL_X8 FILLER_114_279 ();
 FILLCELL_X2 FILLER_114_287 ();
 FILLCELL_X2 FILLER_114_321 ();
 FILLCELL_X1 FILLER_114_323 ();
 FILLCELL_X2 FILLER_114_342 ();
 FILLCELL_X1 FILLER_114_371 ();
 FILLCELL_X8 FILLER_114_385 ();
 FILLCELL_X4 FILLER_114_393 ();
 FILLCELL_X2 FILLER_114_397 ();
 FILLCELL_X1 FILLER_114_399 ();
 FILLCELL_X1 FILLER_114_418 ();
 FILLCELL_X1 FILLER_114_426 ();
 FILLCELL_X1 FILLER_114_430 ();
 FILLCELL_X2 FILLER_114_435 ();
 FILLCELL_X4 FILLER_114_444 ();
 FILLCELL_X2 FILLER_114_448 ();
 FILLCELL_X4 FILLER_114_457 ();
 FILLCELL_X2 FILLER_114_461 ();
 FILLCELL_X8 FILLER_114_483 ();
 FILLCELL_X1 FILLER_114_491 ();
 FILLCELL_X1 FILLER_114_512 ();
 FILLCELL_X16 FILLER_114_521 ();
 FILLCELL_X8 FILLER_114_537 ();
 FILLCELL_X1 FILLER_114_545 ();
 FILLCELL_X8 FILLER_114_553 ();
 FILLCELL_X2 FILLER_114_561 ();
 FILLCELL_X2 FILLER_114_583 ();
 FILLCELL_X8 FILLER_114_596 ();
 FILLCELL_X4 FILLER_114_604 ();
 FILLCELL_X1 FILLER_114_608 ();
 FILLCELL_X4 FILLER_114_614 ();
 FILLCELL_X2 FILLER_114_618 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X16 FILLER_114_632 ();
 FILLCELL_X2 FILLER_114_648 ();
 FILLCELL_X1 FILLER_114_650 ();
 FILLCELL_X8 FILLER_114_671 ();
 FILLCELL_X2 FILLER_114_679 ();
 FILLCELL_X1 FILLER_114_681 ();
 FILLCELL_X1 FILLER_114_708 ();
 FILLCELL_X2 FILLER_114_729 ();
 FILLCELL_X2 FILLER_114_736 ();
 FILLCELL_X2 FILLER_114_758 ();
 FILLCELL_X1 FILLER_114_760 ();
 FILLCELL_X2 FILLER_114_813 ();
 FILLCELL_X4 FILLER_114_821 ();
 FILLCELL_X8 FILLER_114_837 ();
 FILLCELL_X2 FILLER_114_845 ();
 FILLCELL_X4 FILLER_114_851 ();
 FILLCELL_X1 FILLER_114_855 ();
 FILLCELL_X8 FILLER_114_859 ();
 FILLCELL_X4 FILLER_114_867 ();
 FILLCELL_X1 FILLER_114_871 ();
 FILLCELL_X1 FILLER_114_893 ();
 FILLCELL_X2 FILLER_114_904 ();
 FILLCELL_X4 FILLER_114_928 ();
 FILLCELL_X4 FILLER_114_954 ();
 FILLCELL_X4 FILLER_114_980 ();
 FILLCELL_X1 FILLER_114_991 ();
 FILLCELL_X8 FILLER_114_1002 ();
 FILLCELL_X2 FILLER_114_1068 ();
 FILLCELL_X1 FILLER_114_1077 ();
 FILLCELL_X4 FILLER_114_1085 ();
 FILLCELL_X2 FILLER_114_1089 ();
 FILLCELL_X1 FILLER_114_1097 ();
 FILLCELL_X16 FILLER_114_1104 ();
 FILLCELL_X2 FILLER_114_1120 ();
 FILLCELL_X1 FILLER_114_1122 ();
 FILLCELL_X4 FILLER_114_1135 ();
 FILLCELL_X8 FILLER_114_1169 ();
 FILLCELL_X2 FILLER_114_1177 ();
 FILLCELL_X1 FILLER_114_1189 ();
 FILLCELL_X2 FILLER_114_1198 ();
 FILLCELL_X2 FILLER_114_1264 ();
 FILLCELL_X1 FILLER_114_1266 ();
 FILLCELL_X1 FILLER_114_1269 ();
 FILLCELL_X1 FILLER_114_1292 ();
 FILLCELL_X16 FILLER_114_1319 ();
 FILLCELL_X4 FILLER_114_1337 ();
 FILLCELL_X2 FILLER_114_1341 ();
 FILLCELL_X8 FILLER_114_1365 ();
 FILLCELL_X1 FILLER_114_1373 ();
 FILLCELL_X4 FILLER_114_1384 ();
 FILLCELL_X2 FILLER_114_1388 ();
 FILLCELL_X2 FILLER_114_1402 ();
 FILLCELL_X1 FILLER_114_1404 ();
 FILLCELL_X2 FILLER_114_1411 ();
 FILLCELL_X1 FILLER_114_1413 ();
 FILLCELL_X2 FILLER_114_1420 ();
 FILLCELL_X4 FILLER_114_1428 ();
 FILLCELL_X1 FILLER_114_1432 ();
 FILLCELL_X2 FILLER_114_1479 ();
 FILLCELL_X32 FILLER_114_1487 ();
 FILLCELL_X32 FILLER_114_1519 ();
 FILLCELL_X32 FILLER_114_1551 ();
 FILLCELL_X32 FILLER_114_1583 ();
 FILLCELL_X32 FILLER_114_1615 ();
 FILLCELL_X4 FILLER_114_1647 ();
 FILLCELL_X16 FILLER_115_1 ();
 FILLCELL_X8 FILLER_115_17 ();
 FILLCELL_X1 FILLER_115_25 ();
 FILLCELL_X2 FILLER_115_33 ();
 FILLCELL_X16 FILLER_115_39 ();
 FILLCELL_X8 FILLER_115_55 ();
 FILLCELL_X2 FILLER_115_83 ();
 FILLCELL_X8 FILLER_115_132 ();
 FILLCELL_X2 FILLER_115_140 ();
 FILLCELL_X2 FILLER_115_151 ();
 FILLCELL_X4 FILLER_115_173 ();
 FILLCELL_X2 FILLER_115_184 ();
 FILLCELL_X4 FILLER_115_216 ();
 FILLCELL_X2 FILLER_115_220 ();
 FILLCELL_X8 FILLER_115_242 ();
 FILLCELL_X1 FILLER_115_254 ();
 FILLCELL_X8 FILLER_115_283 ();
 FILLCELL_X4 FILLER_115_291 ();
 FILLCELL_X2 FILLER_115_295 ();
 FILLCELL_X1 FILLER_115_300 ();
 FILLCELL_X4 FILLER_115_348 ();
 FILLCELL_X4 FILLER_115_359 ();
 FILLCELL_X2 FILLER_115_363 ();
 FILLCELL_X1 FILLER_115_365 ();
 FILLCELL_X1 FILLER_115_371 ();
 FILLCELL_X4 FILLER_115_398 ();
 FILLCELL_X2 FILLER_115_402 ();
 FILLCELL_X4 FILLER_115_413 ();
 FILLCELL_X2 FILLER_115_417 ();
 FILLCELL_X1 FILLER_115_419 ();
 FILLCELL_X4 FILLER_115_422 ();
 FILLCELL_X2 FILLER_115_434 ();
 FILLCELL_X16 FILLER_115_456 ();
 FILLCELL_X2 FILLER_115_472 ();
 FILLCELL_X1 FILLER_115_474 ();
 FILLCELL_X8 FILLER_115_485 ();
 FILLCELL_X8 FILLER_115_497 ();
 FILLCELL_X2 FILLER_115_505 ();
 FILLCELL_X2 FILLER_115_510 ();
 FILLCELL_X16 FILLER_115_555 ();
 FILLCELL_X1 FILLER_115_591 ();
 FILLCELL_X4 FILLER_115_612 ();
 FILLCELL_X2 FILLER_115_616 ();
 FILLCELL_X1 FILLER_115_618 ();
 FILLCELL_X4 FILLER_115_622 ();
 FILLCELL_X2 FILLER_115_633 ();
 FILLCELL_X1 FILLER_115_635 ();
 FILLCELL_X4 FILLER_115_656 ();
 FILLCELL_X2 FILLER_115_660 ();
 FILLCELL_X2 FILLER_115_702 ();
 FILLCELL_X2 FILLER_115_724 ();
 FILLCELL_X4 FILLER_115_731 ();
 FILLCELL_X16 FILLER_115_742 ();
 FILLCELL_X2 FILLER_115_758 ();
 FILLCELL_X1 FILLER_115_760 ();
 FILLCELL_X8 FILLER_115_768 ();
 FILLCELL_X4 FILLER_115_776 ();
 FILLCELL_X2 FILLER_115_784 ();
 FILLCELL_X2 FILLER_115_793 ();
 FILLCELL_X1 FILLER_115_795 ();
 FILLCELL_X8 FILLER_115_824 ();
 FILLCELL_X4 FILLER_115_832 ();
 FILLCELL_X1 FILLER_115_836 ();
 FILLCELL_X4 FILLER_115_864 ();
 FILLCELL_X2 FILLER_115_868 ();
 FILLCELL_X4 FILLER_115_906 ();
 FILLCELL_X2 FILLER_115_910 ();
 FILLCELL_X8 FILLER_115_956 ();
 FILLCELL_X1 FILLER_115_964 ();
 FILLCELL_X4 FILLER_115_993 ();
 FILLCELL_X2 FILLER_115_1031 ();
 FILLCELL_X2 FILLER_115_1040 ();
 FILLCELL_X2 FILLER_115_1047 ();
 FILLCELL_X1 FILLER_115_1049 ();
 FILLCELL_X1 FILLER_115_1057 ();
 FILLCELL_X2 FILLER_115_1060 ();
 FILLCELL_X2 FILLER_115_1064 ();
 FILLCELL_X4 FILLER_115_1071 ();
 FILLCELL_X8 FILLER_115_1082 ();
 FILLCELL_X4 FILLER_115_1090 ();
 FILLCELL_X2 FILLER_115_1094 ();
 FILLCELL_X4 FILLER_115_1106 ();
 FILLCELL_X2 FILLER_115_1110 ();
 FILLCELL_X1 FILLER_115_1112 ();
 FILLCELL_X4 FILLER_115_1122 ();
 FILLCELL_X1 FILLER_115_1126 ();
 FILLCELL_X2 FILLER_115_1131 ();
 FILLCELL_X4 FILLER_115_1139 ();
 FILLCELL_X2 FILLER_115_1143 ();
 FILLCELL_X1 FILLER_115_1145 ();
 FILLCELL_X1 FILLER_115_1163 ();
 FILLCELL_X8 FILLER_115_1169 ();
 FILLCELL_X4 FILLER_115_1177 ();
 FILLCELL_X4 FILLER_115_1185 ();
 FILLCELL_X1 FILLER_115_1195 ();
 FILLCELL_X4 FILLER_115_1200 ();
 FILLCELL_X2 FILLER_115_1204 ();
 FILLCELL_X1 FILLER_115_1206 ();
 FILLCELL_X4 FILLER_115_1210 ();
 FILLCELL_X2 FILLER_115_1238 ();
 FILLCELL_X2 FILLER_115_1244 ();
 FILLCELL_X4 FILLER_115_1254 ();
 FILLCELL_X1 FILLER_115_1258 ();
 FILLCELL_X2 FILLER_115_1270 ();
 FILLCELL_X1 FILLER_115_1275 ();
 FILLCELL_X2 FILLER_115_1283 ();
 FILLCELL_X1 FILLER_115_1285 ();
 FILLCELL_X2 FILLER_115_1295 ();
 FILLCELL_X1 FILLER_115_1297 ();
 FILLCELL_X2 FILLER_115_1304 ();
 FILLCELL_X1 FILLER_115_1306 ();
 FILLCELL_X1 FILLER_115_1313 ();
 FILLCELL_X8 FILLER_115_1359 ();
 FILLCELL_X1 FILLER_115_1379 ();
 FILLCELL_X1 FILLER_115_1396 ();
 FILLCELL_X1 FILLER_115_1403 ();
 FILLCELL_X1 FILLER_115_1410 ();
 FILLCELL_X4 FILLER_115_1417 ();
 FILLCELL_X2 FILLER_115_1421 ();
 FILLCELL_X1 FILLER_115_1423 ();
 FILLCELL_X2 FILLER_115_1434 ();
 FILLCELL_X1 FILLER_115_1436 ();
 FILLCELL_X2 FILLER_115_1447 ();
 FILLCELL_X2 FILLER_115_1459 ();
 FILLCELL_X1 FILLER_115_1461 ();
 FILLCELL_X2 FILLER_115_1468 ();
 FILLCELL_X1 FILLER_115_1470 ();
 FILLCELL_X2 FILLER_115_1481 ();
 FILLCELL_X32 FILLER_115_1492 ();
 FILLCELL_X32 FILLER_115_1524 ();
 FILLCELL_X32 FILLER_115_1556 ();
 FILLCELL_X32 FILLER_115_1588 ();
 FILLCELL_X16 FILLER_115_1620 ();
 FILLCELL_X8 FILLER_115_1636 ();
 FILLCELL_X4 FILLER_115_1644 ();
 FILLCELL_X2 FILLER_115_1648 ();
 FILLCELL_X1 FILLER_115_1650 ();
 FILLCELL_X8 FILLER_116_1 ();
 FILLCELL_X4 FILLER_116_9 ();
 FILLCELL_X1 FILLER_116_40 ();
 FILLCELL_X1 FILLER_116_81 ();
 FILLCELL_X1 FILLER_116_91 ();
 FILLCELL_X1 FILLER_116_99 ();
 FILLCELL_X1 FILLER_116_117 ();
 FILLCELL_X8 FILLER_116_141 ();
 FILLCELL_X2 FILLER_116_149 ();
 FILLCELL_X4 FILLER_116_158 ();
 FILLCELL_X2 FILLER_116_169 ();
 FILLCELL_X2 FILLER_116_176 ();
 FILLCELL_X1 FILLER_116_178 ();
 FILLCELL_X1 FILLER_116_199 ();
 FILLCELL_X2 FILLER_116_205 ();
 FILLCELL_X1 FILLER_116_207 ();
 FILLCELL_X4 FILLER_116_215 ();
 FILLCELL_X1 FILLER_116_219 ();
 FILLCELL_X4 FILLER_116_233 ();
 FILLCELL_X8 FILLER_116_265 ();
 FILLCELL_X2 FILLER_116_297 ();
 FILLCELL_X2 FILLER_116_307 ();
 FILLCELL_X1 FILLER_116_309 ();
 FILLCELL_X8 FILLER_116_313 ();
 FILLCELL_X4 FILLER_116_324 ();
 FILLCELL_X8 FILLER_116_333 ();
 FILLCELL_X2 FILLER_116_341 ();
 FILLCELL_X1 FILLER_116_343 ();
 FILLCELL_X2 FILLER_116_353 ();
 FILLCELL_X1 FILLER_116_355 ();
 FILLCELL_X8 FILLER_116_359 ();
 FILLCELL_X4 FILLER_116_367 ();
 FILLCELL_X1 FILLER_116_371 ();
 FILLCELL_X2 FILLER_116_397 ();
 FILLCELL_X1 FILLER_116_399 ();
 FILLCELL_X2 FILLER_116_409 ();
 FILLCELL_X1 FILLER_116_411 ();
 FILLCELL_X2 FILLER_116_432 ();
 FILLCELL_X1 FILLER_116_434 ();
 FILLCELL_X2 FILLER_116_467 ();
 FILLCELL_X1 FILLER_116_472 ();
 FILLCELL_X8 FILLER_116_480 ();
 FILLCELL_X2 FILLER_116_488 ();
 FILLCELL_X1 FILLER_116_490 ();
 FILLCELL_X1 FILLER_116_496 ();
 FILLCELL_X4 FILLER_116_520 ();
 FILLCELL_X1 FILLER_116_535 ();
 FILLCELL_X1 FILLER_116_539 ();
 FILLCELL_X8 FILLER_116_564 ();
 FILLCELL_X8 FILLER_116_576 ();
 FILLCELL_X4 FILLER_116_584 ();
 FILLCELL_X2 FILLER_116_592 ();
 FILLCELL_X1 FILLER_116_594 ();
 FILLCELL_X2 FILLER_116_632 ();
 FILLCELL_X2 FILLER_116_646 ();
 FILLCELL_X1 FILLER_116_648 ();
 FILLCELL_X2 FILLER_116_680 ();
 FILLCELL_X4 FILLER_116_688 ();
 FILLCELL_X4 FILLER_116_697 ();
 FILLCELL_X2 FILLER_116_701 ();
 FILLCELL_X1 FILLER_116_703 ();
 FILLCELL_X4 FILLER_116_707 ();
 FILLCELL_X1 FILLER_116_711 ();
 FILLCELL_X2 FILLER_116_715 ();
 FILLCELL_X8 FILLER_116_767 ();
 FILLCELL_X2 FILLER_116_802 ();
 FILLCELL_X8 FILLER_116_834 ();
 FILLCELL_X16 FILLER_116_892 ();
 FILLCELL_X2 FILLER_116_908 ();
 FILLCELL_X8 FILLER_116_923 ();
 FILLCELL_X1 FILLER_116_931 ();
 FILLCELL_X8 FILLER_116_939 ();
 FILLCELL_X4 FILLER_116_947 ();
 FILLCELL_X8 FILLER_116_960 ();
 FILLCELL_X2 FILLER_116_968 ();
 FILLCELL_X1 FILLER_116_970 ();
 FILLCELL_X8 FILLER_116_1031 ();
 FILLCELL_X4 FILLER_116_1039 ();
 FILLCELL_X1 FILLER_116_1050 ();
 FILLCELL_X2 FILLER_116_1071 ();
 FILLCELL_X4 FILLER_116_1080 ();
 FILLCELL_X2 FILLER_116_1084 ();
 FILLCELL_X4 FILLER_116_1114 ();
 FILLCELL_X2 FILLER_116_1118 ();
 FILLCELL_X1 FILLER_116_1141 ();
 FILLCELL_X4 FILLER_116_1152 ();
 FILLCELL_X2 FILLER_116_1156 ();
 FILLCELL_X1 FILLER_116_1158 ();
 FILLCELL_X2 FILLER_116_1180 ();
 FILLCELL_X2 FILLER_116_1204 ();
 FILLCELL_X1 FILLER_116_1206 ();
 FILLCELL_X8 FILLER_116_1229 ();
 FILLCELL_X1 FILLER_116_1237 ();
 FILLCELL_X1 FILLER_116_1301 ();
 FILLCELL_X1 FILLER_116_1313 ();
 FILLCELL_X1 FILLER_116_1319 ();
 FILLCELL_X8 FILLER_116_1325 ();
 FILLCELL_X4 FILLER_116_1336 ();
 FILLCELL_X1 FILLER_116_1340 ();
 FILLCELL_X4 FILLER_116_1385 ();
 FILLCELL_X1 FILLER_116_1389 ();
 FILLCELL_X4 FILLER_116_1400 ();
 FILLCELL_X1 FILLER_116_1404 ();
 FILLCELL_X4 FILLER_116_1415 ();
 FILLCELL_X4 FILLER_116_1425 ();
 FILLCELL_X4 FILLER_116_1435 ();
 FILLCELL_X2 FILLER_116_1461 ();
 FILLCELL_X1 FILLER_116_1469 ();
 FILLCELL_X32 FILLER_116_1480 ();
 FILLCELL_X32 FILLER_116_1512 ();
 FILLCELL_X32 FILLER_116_1544 ();
 FILLCELL_X32 FILLER_116_1576 ();
 FILLCELL_X32 FILLER_116_1608 ();
 FILLCELL_X8 FILLER_116_1640 ();
 FILLCELL_X2 FILLER_116_1648 ();
 FILLCELL_X1 FILLER_116_1650 ();
 FILLCELL_X1 FILLER_117_1 ();
 FILLCELL_X2 FILLER_117_29 ();
 FILLCELL_X1 FILLER_117_31 ();
 FILLCELL_X8 FILLER_117_51 ();
 FILLCELL_X2 FILLER_117_59 ();
 FILLCELL_X1 FILLER_117_61 ();
 FILLCELL_X1 FILLER_117_105 ();
 FILLCELL_X8 FILLER_117_114 ();
 FILLCELL_X2 FILLER_117_122 ();
 FILLCELL_X1 FILLER_117_124 ();
 FILLCELL_X1 FILLER_117_152 ();
 FILLCELL_X2 FILLER_117_160 ();
 FILLCELL_X8 FILLER_117_182 ();
 FILLCELL_X2 FILLER_117_190 ();
 FILLCELL_X4 FILLER_117_261 ();
 FILLCELL_X2 FILLER_117_265 ();
 FILLCELL_X1 FILLER_117_275 ();
 FILLCELL_X2 FILLER_117_333 ();
 FILLCELL_X8 FILLER_117_409 ();
 FILLCELL_X4 FILLER_117_417 ();
 FILLCELL_X2 FILLER_117_421 ();
 FILLCELL_X1 FILLER_117_423 ();
 FILLCELL_X8 FILLER_117_431 ();
 FILLCELL_X2 FILLER_117_439 ();
 FILLCELL_X1 FILLER_117_441 ();
 FILLCELL_X1 FILLER_117_454 ();
 FILLCELL_X1 FILLER_117_482 ();
 FILLCELL_X1 FILLER_117_503 ();
 FILLCELL_X2 FILLER_117_516 ();
 FILLCELL_X8 FILLER_117_534 ();
 FILLCELL_X2 FILLER_117_542 ();
 FILLCELL_X1 FILLER_117_544 ();
 FILLCELL_X1 FILLER_117_555 ();
 FILLCELL_X8 FILLER_117_576 ();
 FILLCELL_X2 FILLER_117_584 ();
 FILLCELL_X1 FILLER_117_642 ();
 FILLCELL_X4 FILLER_117_690 ();
 FILLCELL_X1 FILLER_117_694 ();
 FILLCELL_X4 FILLER_117_712 ();
 FILLCELL_X2 FILLER_117_716 ();
 FILLCELL_X1 FILLER_117_718 ();
 FILLCELL_X2 FILLER_117_726 ();
 FILLCELL_X1 FILLER_117_728 ();
 FILLCELL_X2 FILLER_117_738 ();
 FILLCELL_X8 FILLER_117_767 ();
 FILLCELL_X2 FILLER_117_779 ();
 FILLCELL_X4 FILLER_117_810 ();
 FILLCELL_X8 FILLER_117_821 ();
 FILLCELL_X4 FILLER_117_829 ();
 FILLCELL_X2 FILLER_117_833 ();
 FILLCELL_X8 FILLER_117_865 ();
 FILLCELL_X2 FILLER_117_873 ();
 FILLCELL_X1 FILLER_117_875 ();
 FILLCELL_X4 FILLER_117_879 ();
 FILLCELL_X1 FILLER_117_883 ();
 FILLCELL_X2 FILLER_117_916 ();
 FILLCELL_X8 FILLER_117_953 ();
 FILLCELL_X1 FILLER_117_985 ();
 FILLCELL_X8 FILLER_117_993 ();
 FILLCELL_X1 FILLER_117_1001 ();
 FILLCELL_X8 FILLER_117_1009 ();
 FILLCELL_X8 FILLER_117_1024 ();
 FILLCELL_X1 FILLER_117_1032 ();
 FILLCELL_X4 FILLER_117_1042 ();
 FILLCELL_X8 FILLER_117_1068 ();
 FILLCELL_X1 FILLER_117_1076 ();
 FILLCELL_X1 FILLER_117_1110 ();
 FILLCELL_X1 FILLER_117_1145 ();
 FILLCELL_X8 FILLER_117_1153 ();
 FILLCELL_X4 FILLER_117_1161 ();
 FILLCELL_X1 FILLER_117_1165 ();
 FILLCELL_X4 FILLER_117_1171 ();
 FILLCELL_X2 FILLER_117_1175 ();
 FILLCELL_X1 FILLER_117_1189 ();
 FILLCELL_X8 FILLER_117_1195 ();
 FILLCELL_X1 FILLER_117_1203 ();
 FILLCELL_X2 FILLER_117_1208 ();
 FILLCELL_X1 FILLER_117_1236 ();
 FILLCELL_X2 FILLER_117_1243 ();
 FILLCELL_X1 FILLER_117_1245 ();
 FILLCELL_X2 FILLER_117_1253 ();
 FILLCELL_X8 FILLER_117_1264 ();
 FILLCELL_X2 FILLER_117_1272 ();
 FILLCELL_X2 FILLER_117_1296 ();
 FILLCELL_X2 FILLER_117_1305 ();
 FILLCELL_X4 FILLER_117_1313 ();
 FILLCELL_X8 FILLER_117_1319 ();
 FILLCELL_X4 FILLER_117_1327 ();
 FILLCELL_X1 FILLER_117_1331 ();
 FILLCELL_X1 FILLER_117_1348 ();
 FILLCELL_X4 FILLER_117_1362 ();
 FILLCELL_X2 FILLER_117_1366 ();
 FILLCELL_X2 FILLER_117_1396 ();
 FILLCELL_X4 FILLER_117_1410 ();
 FILLCELL_X2 FILLER_117_1414 ();
 FILLCELL_X1 FILLER_117_1416 ();
 FILLCELL_X4 FILLER_117_1427 ();
 FILLCELL_X8 FILLER_117_1453 ();
 FILLCELL_X4 FILLER_117_1461 ();
 FILLCELL_X2 FILLER_117_1465 ();
 FILLCELL_X1 FILLER_117_1467 ();
 FILLCELL_X32 FILLER_117_1480 ();
 FILLCELL_X32 FILLER_117_1512 ();
 FILLCELL_X32 FILLER_117_1544 ();
 FILLCELL_X32 FILLER_117_1576 ();
 FILLCELL_X32 FILLER_117_1608 ();
 FILLCELL_X8 FILLER_117_1640 ();
 FILLCELL_X2 FILLER_117_1648 ();
 FILLCELL_X1 FILLER_117_1650 ();
 FILLCELL_X2 FILLER_118_1 ();
 FILLCELL_X1 FILLER_118_3 ();
 FILLCELL_X4 FILLER_118_31 ();
 FILLCELL_X2 FILLER_118_55 ();
 FILLCELL_X1 FILLER_118_71 ();
 FILLCELL_X4 FILLER_118_79 ();
 FILLCELL_X8 FILLER_118_114 ();
 FILLCELL_X1 FILLER_118_122 ();
 FILLCELL_X8 FILLER_118_167 ();
 FILLCELL_X2 FILLER_118_175 ();
 FILLCELL_X4 FILLER_118_184 ();
 FILLCELL_X16 FILLER_118_195 ();
 FILLCELL_X8 FILLER_118_211 ();
 FILLCELL_X4 FILLER_118_219 ();
 FILLCELL_X2 FILLER_118_223 ();
 FILLCELL_X1 FILLER_118_225 ();
 FILLCELL_X2 FILLER_118_230 ();
 FILLCELL_X8 FILLER_118_235 ();
 FILLCELL_X1 FILLER_118_243 ();
 FILLCELL_X8 FILLER_118_253 ();
 FILLCELL_X1 FILLER_118_295 ();
 FILLCELL_X8 FILLER_118_335 ();
 FILLCELL_X1 FILLER_118_343 ();
 FILLCELL_X2 FILLER_118_346 ();
 FILLCELL_X4 FILLER_118_368 ();
 FILLCELL_X1 FILLER_118_372 ();
 FILLCELL_X4 FILLER_118_377 ();
 FILLCELL_X2 FILLER_118_391 ();
 FILLCELL_X1 FILLER_118_397 ();
 FILLCELL_X1 FILLER_118_410 ();
 FILLCELL_X8 FILLER_118_415 ();
 FILLCELL_X2 FILLER_118_423 ();
 FILLCELL_X4 FILLER_118_476 ();
 FILLCELL_X2 FILLER_118_480 ();
 FILLCELL_X1 FILLER_118_485 ();
 FILLCELL_X2 FILLER_118_511 ();
 FILLCELL_X1 FILLER_118_513 ();
 FILLCELL_X16 FILLER_118_531 ();
 FILLCELL_X16 FILLER_118_582 ();
 FILLCELL_X8 FILLER_118_598 ();
 FILLCELL_X4 FILLER_118_606 ();
 FILLCELL_X2 FILLER_118_610 ();
 FILLCELL_X4 FILLER_118_620 ();
 FILLCELL_X2 FILLER_118_624 ();
 FILLCELL_X1 FILLER_118_626 ();
 FILLCELL_X2 FILLER_118_632 ();
 FILLCELL_X1 FILLER_118_634 ();
 FILLCELL_X4 FILLER_118_638 ();
 FILLCELL_X2 FILLER_118_642 ();
 FILLCELL_X1 FILLER_118_644 ();
 FILLCELL_X4 FILLER_118_670 ();
 FILLCELL_X1 FILLER_118_698 ();
 FILLCELL_X8 FILLER_118_703 ();
 FILLCELL_X1 FILLER_118_711 ();
 FILLCELL_X1 FILLER_118_732 ();
 FILLCELL_X1 FILLER_118_738 ();
 FILLCELL_X16 FILLER_118_744 ();
 FILLCELL_X8 FILLER_118_760 ();
 FILLCELL_X8 FILLER_118_792 ();
 FILLCELL_X1 FILLER_118_800 ();
 FILLCELL_X4 FILLER_118_819 ();
 FILLCELL_X1 FILLER_118_823 ();
 FILLCELL_X1 FILLER_118_851 ();
 FILLCELL_X8 FILLER_118_861 ();
 FILLCELL_X4 FILLER_118_869 ();
 FILLCELL_X1 FILLER_118_873 ();
 FILLCELL_X4 FILLER_118_896 ();
 FILLCELL_X1 FILLER_118_900 ();
 FILLCELL_X32 FILLER_118_921 ();
 FILLCELL_X8 FILLER_118_953 ();
 FILLCELL_X4 FILLER_118_961 ();
 FILLCELL_X4 FILLER_118_987 ();
 FILLCELL_X1 FILLER_118_991 ();
 FILLCELL_X2 FILLER_118_1014 ();
 FILLCELL_X4 FILLER_118_1050 ();
 FILLCELL_X2 FILLER_118_1054 ();
 FILLCELL_X1 FILLER_118_1056 ();
 FILLCELL_X8 FILLER_118_1109 ();
 FILLCELL_X1 FILLER_118_1117 ();
 FILLCELL_X4 FILLER_118_1127 ();
 FILLCELL_X8 FILLER_118_1177 ();
 FILLCELL_X4 FILLER_118_1185 ();
 FILLCELL_X2 FILLER_118_1189 ();
 FILLCELL_X2 FILLER_118_1219 ();
 FILLCELL_X1 FILLER_118_1221 ();
 FILLCELL_X2 FILLER_118_1253 ();
 FILLCELL_X1 FILLER_118_1255 ();
 FILLCELL_X2 FILLER_118_1264 ();
 FILLCELL_X1 FILLER_118_1266 ();
 FILLCELL_X8 FILLER_118_1271 ();
 FILLCELL_X1 FILLER_118_1279 ();
 FILLCELL_X4 FILLER_118_1285 ();
 FILLCELL_X1 FILLER_118_1289 ();
 FILLCELL_X2 FILLER_118_1293 ();
 FILLCELL_X1 FILLER_118_1295 ();
 FILLCELL_X2 FILLER_118_1303 ();
 FILLCELL_X8 FILLER_118_1360 ();
 FILLCELL_X4 FILLER_118_1368 ();
 FILLCELL_X2 FILLER_118_1372 ();
 FILLCELL_X1 FILLER_118_1392 ();
 FILLCELL_X8 FILLER_118_1399 ();
 FILLCELL_X1 FILLER_118_1413 ();
 FILLCELL_X2 FILLER_118_1454 ();
 FILLCELL_X1 FILLER_118_1456 ();
 FILLCELL_X32 FILLER_118_1487 ();
 FILLCELL_X32 FILLER_118_1519 ();
 FILLCELL_X32 FILLER_118_1551 ();
 FILLCELL_X32 FILLER_118_1583 ();
 FILLCELL_X32 FILLER_118_1615 ();
 FILLCELL_X4 FILLER_118_1647 ();
 FILLCELL_X8 FILLER_119_37 ();
 FILLCELL_X2 FILLER_119_45 ();
 FILLCELL_X16 FILLER_119_54 ();
 FILLCELL_X8 FILLER_119_70 ();
 FILLCELL_X2 FILLER_119_78 ();
 FILLCELL_X1 FILLER_119_80 ();
 FILLCELL_X4 FILLER_119_94 ();
 FILLCELL_X2 FILLER_119_98 ();
 FILLCELL_X4 FILLER_119_120 ();
 FILLCELL_X4 FILLER_119_142 ();
 FILLCELL_X2 FILLER_119_146 ();
 FILLCELL_X1 FILLER_119_155 ();
 FILLCELL_X2 FILLER_119_163 ();
 FILLCELL_X2 FILLER_119_185 ();
 FILLCELL_X1 FILLER_119_187 ();
 FILLCELL_X16 FILLER_119_208 ();
 FILLCELL_X2 FILLER_119_247 ();
 FILLCELL_X2 FILLER_119_260 ();
 FILLCELL_X1 FILLER_119_262 ();
 FILLCELL_X2 FILLER_119_266 ();
 FILLCELL_X1 FILLER_119_268 ();
 FILLCELL_X1 FILLER_119_276 ();
 FILLCELL_X2 FILLER_119_300 ();
 FILLCELL_X2 FILLER_119_322 ();
 FILLCELL_X1 FILLER_119_331 ();
 FILLCELL_X2 FILLER_119_352 ();
 FILLCELL_X4 FILLER_119_361 ();
 FILLCELL_X1 FILLER_119_365 ();
 FILLCELL_X16 FILLER_119_370 ();
 FILLCELL_X8 FILLER_119_386 ();
 FILLCELL_X4 FILLER_119_394 ();
 FILLCELL_X2 FILLER_119_398 ();
 FILLCELL_X8 FILLER_119_408 ();
 FILLCELL_X4 FILLER_119_416 ();
 FILLCELL_X1 FILLER_119_440 ();
 FILLCELL_X8 FILLER_119_448 ();
 FILLCELL_X1 FILLER_119_461 ();
 FILLCELL_X1 FILLER_119_537 ();
 FILLCELL_X2 FILLER_119_567 ();
 FILLCELL_X1 FILLER_119_609 ();
 FILLCELL_X16 FILLER_119_637 ();
 FILLCELL_X1 FILLER_119_653 ();
 FILLCELL_X8 FILLER_119_668 ();
 FILLCELL_X1 FILLER_119_683 ();
 FILLCELL_X2 FILLER_119_689 ();
 FILLCELL_X1 FILLER_119_711 ();
 FILLCELL_X2 FILLER_119_722 ();
 FILLCELL_X8 FILLER_119_763 ();
 FILLCELL_X2 FILLER_119_771 ();
 FILLCELL_X1 FILLER_119_783 ();
 FILLCELL_X2 FILLER_119_811 ();
 FILLCELL_X1 FILLER_119_813 ();
 FILLCELL_X4 FILLER_119_821 ();
 FILLCELL_X1 FILLER_119_825 ();
 FILLCELL_X8 FILLER_119_846 ();
 FILLCELL_X4 FILLER_119_854 ();
 FILLCELL_X1 FILLER_119_858 ();
 FILLCELL_X16 FILLER_119_862 ();
 FILLCELL_X8 FILLER_119_878 ();
 FILLCELL_X4 FILLER_119_886 ();
 FILLCELL_X2 FILLER_119_890 ();
 FILLCELL_X4 FILLER_119_905 ();
 FILLCELL_X1 FILLER_119_909 ();
 FILLCELL_X8 FILLER_119_930 ();
 FILLCELL_X2 FILLER_119_938 ();
 FILLCELL_X2 FILLER_119_969 ();
 FILLCELL_X16 FILLER_119_993 ();
 FILLCELL_X4 FILLER_119_1038 ();
 FILLCELL_X16 FILLER_119_1084 ();
 FILLCELL_X2 FILLER_119_1100 ();
 FILLCELL_X2 FILLER_119_1108 ();
 FILLCELL_X1 FILLER_119_1110 ();
 FILLCELL_X4 FILLER_119_1121 ();
 FILLCELL_X1 FILLER_119_1125 ();
 FILLCELL_X4 FILLER_119_1148 ();
 FILLCELL_X4 FILLER_119_1162 ();
 FILLCELL_X1 FILLER_119_1166 ();
 FILLCELL_X2 FILLER_119_1171 ();
 FILLCELL_X4 FILLER_119_1177 ();
 FILLCELL_X1 FILLER_119_1181 ();
 FILLCELL_X1 FILLER_119_1204 ();
 FILLCELL_X2 FILLER_119_1222 ();
 FILLCELL_X8 FILLER_119_1227 ();
 FILLCELL_X4 FILLER_119_1235 ();
 FILLCELL_X1 FILLER_119_1239 ();
 FILLCELL_X4 FILLER_119_1247 ();
 FILLCELL_X2 FILLER_119_1251 ();
 FILLCELL_X4 FILLER_119_1256 ();
 FILLCELL_X2 FILLER_119_1260 ();
 FILLCELL_X1 FILLER_119_1262 ();
 FILLCELL_X2 FILLER_119_1264 ();
 FILLCELL_X1 FILLER_119_1266 ();
 FILLCELL_X4 FILLER_119_1275 ();
 FILLCELL_X1 FILLER_119_1290 ();
 FILLCELL_X4 FILLER_119_1317 ();
 FILLCELL_X1 FILLER_119_1321 ();
 FILLCELL_X2 FILLER_119_1344 ();
 FILLCELL_X1 FILLER_119_1346 ();
 FILLCELL_X4 FILLER_119_1351 ();
 FILLCELL_X8 FILLER_119_1358 ();
 FILLCELL_X4 FILLER_119_1366 ();
 FILLCELL_X1 FILLER_119_1473 ();
 FILLCELL_X32 FILLER_119_1480 ();
 FILLCELL_X32 FILLER_119_1512 ();
 FILLCELL_X32 FILLER_119_1544 ();
 FILLCELL_X32 FILLER_119_1576 ();
 FILLCELL_X32 FILLER_119_1608 ();
 FILLCELL_X8 FILLER_119_1640 ();
 FILLCELL_X2 FILLER_119_1648 ();
 FILLCELL_X1 FILLER_119_1650 ();
 FILLCELL_X8 FILLER_120_1 ();
 FILLCELL_X2 FILLER_120_89 ();
 FILLCELL_X4 FILLER_120_96 ();
 FILLCELL_X16 FILLER_120_113 ();
 FILLCELL_X4 FILLER_120_149 ();
 FILLCELL_X1 FILLER_120_153 ();
 FILLCELL_X2 FILLER_120_179 ();
 FILLCELL_X1 FILLER_120_333 ();
 FILLCELL_X2 FILLER_120_354 ();
 FILLCELL_X1 FILLER_120_356 ();
 FILLCELL_X1 FILLER_120_377 ();
 FILLCELL_X2 FILLER_120_409 ();
 FILLCELL_X1 FILLER_120_411 ();
 FILLCELL_X4 FILLER_120_436 ();
 FILLCELL_X4 FILLER_120_484 ();
 FILLCELL_X2 FILLER_120_488 ();
 FILLCELL_X2 FILLER_120_492 ();
 FILLCELL_X4 FILLER_120_501 ();
 FILLCELL_X4 FILLER_120_510 ();
 FILLCELL_X1 FILLER_120_566 ();
 FILLCELL_X8 FILLER_120_639 ();
 FILLCELL_X2 FILLER_120_647 ();
 FILLCELL_X1 FILLER_120_649 ();
 FILLCELL_X8 FILLER_120_690 ();
 FILLCELL_X2 FILLER_120_698 ();
 FILLCELL_X1 FILLER_120_700 ();
 FILLCELL_X1 FILLER_120_704 ();
 FILLCELL_X4 FILLER_120_709 ();
 FILLCELL_X2 FILLER_120_713 ();
 FILLCELL_X1 FILLER_120_715 ();
 FILLCELL_X8 FILLER_120_743 ();
 FILLCELL_X1 FILLER_120_751 ();
 FILLCELL_X2 FILLER_120_783 ();
 FILLCELL_X2 FILLER_120_794 ();
 FILLCELL_X1 FILLER_120_796 ();
 FILLCELL_X2 FILLER_120_826 ();
 FILLCELL_X1 FILLER_120_828 ();
 FILLCELL_X4 FILLER_120_836 ();
 FILLCELL_X2 FILLER_120_840 ();
 FILLCELL_X2 FILLER_120_845 ();
 FILLCELL_X1 FILLER_120_847 ();
 FILLCELL_X2 FILLER_120_885 ();
 FILLCELL_X2 FILLER_120_927 ();
 FILLCELL_X16 FILLER_120_938 ();
 FILLCELL_X8 FILLER_120_954 ();
 FILLCELL_X2 FILLER_120_962 ();
 FILLCELL_X8 FILLER_120_978 ();
 FILLCELL_X1 FILLER_120_993 ();
 FILLCELL_X4 FILLER_120_1004 ();
 FILLCELL_X2 FILLER_120_1008 ();
 FILLCELL_X8 FILLER_120_1048 ();
 FILLCELL_X2 FILLER_120_1056 ();
 FILLCELL_X1 FILLER_120_1065 ();
 FILLCELL_X2 FILLER_120_1068 ();
 FILLCELL_X1 FILLER_120_1070 ();
 FILLCELL_X4 FILLER_120_1106 ();
 FILLCELL_X2 FILLER_120_1110 ();
 FILLCELL_X1 FILLER_120_1112 ();
 FILLCELL_X8 FILLER_120_1119 ();
 FILLCELL_X1 FILLER_120_1127 ();
 FILLCELL_X8 FILLER_120_1134 ();
 FILLCELL_X2 FILLER_120_1142 ();
 FILLCELL_X1 FILLER_120_1144 ();
 FILLCELL_X4 FILLER_120_1148 ();
 FILLCELL_X4 FILLER_120_1163 ();
 FILLCELL_X2 FILLER_120_1167 ();
 FILLCELL_X1 FILLER_120_1169 ();
 FILLCELL_X2 FILLER_120_1176 ();
 FILLCELL_X1 FILLER_120_1178 ();
 FILLCELL_X4 FILLER_120_1182 ();
 FILLCELL_X1 FILLER_120_1186 ();
 FILLCELL_X4 FILLER_120_1198 ();
 FILLCELL_X2 FILLER_120_1202 ();
 FILLCELL_X1 FILLER_120_1235 ();
 FILLCELL_X1 FILLER_120_1243 ();
 FILLCELL_X1 FILLER_120_1256 ();
 FILLCELL_X1 FILLER_120_1261 ();
 FILLCELL_X8 FILLER_120_1274 ();
 FILLCELL_X1 FILLER_120_1294 ();
 FILLCELL_X2 FILLER_120_1299 ();
 FILLCELL_X2 FILLER_120_1311 ();
 FILLCELL_X1 FILLER_120_1313 ();
 FILLCELL_X4 FILLER_120_1321 ();
 FILLCELL_X1 FILLER_120_1325 ();
 FILLCELL_X4 FILLER_120_1329 ();
 FILLCELL_X2 FILLER_120_1340 ();
 FILLCELL_X1 FILLER_120_1342 ();
 FILLCELL_X2 FILLER_120_1395 ();
 FILLCELL_X2 FILLER_120_1429 ();
 FILLCELL_X2 FILLER_120_1453 ();
 FILLCELL_X1 FILLER_120_1471 ();
 FILLCELL_X2 FILLER_120_1478 ();
 FILLCELL_X32 FILLER_120_1486 ();
 FILLCELL_X32 FILLER_120_1518 ();
 FILLCELL_X32 FILLER_120_1550 ();
 FILLCELL_X32 FILLER_120_1582 ();
 FILLCELL_X32 FILLER_120_1614 ();
 FILLCELL_X4 FILLER_120_1646 ();
 FILLCELL_X1 FILLER_120_1650 ();
 FILLCELL_X16 FILLER_121_1 ();
 FILLCELL_X8 FILLER_121_44 ();
 FILLCELL_X2 FILLER_121_52 ();
 FILLCELL_X1 FILLER_121_61 ();
 FILLCELL_X2 FILLER_121_66 ();
 FILLCELL_X1 FILLER_121_68 ();
 FILLCELL_X1 FILLER_121_82 ();
 FILLCELL_X1 FILLER_121_90 ();
 FILLCELL_X2 FILLER_121_111 ();
 FILLCELL_X4 FILLER_121_158 ();
 FILLCELL_X1 FILLER_121_162 ();
 FILLCELL_X2 FILLER_121_170 ();
 FILLCELL_X1 FILLER_121_189 ();
 FILLCELL_X2 FILLER_121_195 ();
 FILLCELL_X1 FILLER_121_197 ();
 FILLCELL_X1 FILLER_121_236 ();
 FILLCELL_X2 FILLER_121_241 ();
 FILLCELL_X4 FILLER_121_252 ();
 FILLCELL_X2 FILLER_121_256 ();
 FILLCELL_X1 FILLER_121_258 ();
 FILLCELL_X4 FILLER_121_263 ();
 FILLCELL_X1 FILLER_121_267 ();
 FILLCELL_X4 FILLER_121_271 ();
 FILLCELL_X1 FILLER_121_275 ();
 FILLCELL_X8 FILLER_121_299 ();
 FILLCELL_X1 FILLER_121_307 ();
 FILLCELL_X8 FILLER_121_317 ();
 FILLCELL_X1 FILLER_121_350 ();
 FILLCELL_X4 FILLER_121_355 ();
 FILLCELL_X2 FILLER_121_359 ();
 FILLCELL_X1 FILLER_121_361 ();
 FILLCELL_X2 FILLER_121_365 ();
 FILLCELL_X1 FILLER_121_367 ();
 FILLCELL_X2 FILLER_121_371 ();
 FILLCELL_X1 FILLER_121_397 ();
 FILLCELL_X16 FILLER_121_410 ();
 FILLCELL_X4 FILLER_121_426 ();
 FILLCELL_X2 FILLER_121_430 ();
 FILLCELL_X4 FILLER_121_450 ();
 FILLCELL_X2 FILLER_121_454 ();
 FILLCELL_X1 FILLER_121_456 ();
 FILLCELL_X16 FILLER_121_472 ();
 FILLCELL_X8 FILLER_121_488 ();
 FILLCELL_X2 FILLER_121_496 ();
 FILLCELL_X1 FILLER_121_498 ();
 FILLCELL_X2 FILLER_121_508 ();
 FILLCELL_X4 FILLER_121_517 ();
 FILLCELL_X2 FILLER_121_521 ();
 FILLCELL_X1 FILLER_121_544 ();
 FILLCELL_X2 FILLER_121_548 ();
 FILLCELL_X2 FILLER_121_555 ();
 FILLCELL_X1 FILLER_121_557 ();
 FILLCELL_X4 FILLER_121_583 ();
 FILLCELL_X2 FILLER_121_587 ();
 FILLCELL_X1 FILLER_121_593 ();
 FILLCELL_X16 FILLER_121_597 ();
 FILLCELL_X8 FILLER_121_613 ();
 FILLCELL_X2 FILLER_121_621 ();
 FILLCELL_X16 FILLER_121_633 ();
 FILLCELL_X4 FILLER_121_649 ();
 FILLCELL_X1 FILLER_121_653 ();
 FILLCELL_X2 FILLER_121_674 ();
 FILLCELL_X1 FILLER_121_676 ();
 FILLCELL_X1 FILLER_121_692 ();
 FILLCELL_X8 FILLER_121_698 ();
 FILLCELL_X2 FILLER_121_729 ();
 FILLCELL_X8 FILLER_121_756 ();
 FILLCELL_X4 FILLER_121_764 ();
 FILLCELL_X4 FILLER_121_795 ();
 FILLCELL_X2 FILLER_121_799 ();
 FILLCELL_X1 FILLER_121_808 ();
 FILLCELL_X2 FILLER_121_812 ();
 FILLCELL_X4 FILLER_121_817 ();
 FILLCELL_X1 FILLER_121_821 ();
 FILLCELL_X4 FILLER_121_842 ();
 FILLCELL_X1 FILLER_121_846 ();
 FILLCELL_X8 FILLER_121_871 ();
 FILLCELL_X4 FILLER_121_879 ();
 FILLCELL_X2 FILLER_121_883 ();
 FILLCELL_X1 FILLER_121_892 ();
 FILLCELL_X2 FILLER_121_900 ();
 FILLCELL_X4 FILLER_121_912 ();
 FILLCELL_X1 FILLER_121_916 ();
 FILLCELL_X4 FILLER_121_921 ();
 FILLCELL_X1 FILLER_121_925 ();
 FILLCELL_X2 FILLER_121_1011 ();
 FILLCELL_X4 FILLER_121_1023 ();
 FILLCELL_X2 FILLER_121_1027 ();
 FILLCELL_X4 FILLER_121_1036 ();
 FILLCELL_X2 FILLER_121_1040 ();
 FILLCELL_X8 FILLER_121_1064 ();
 FILLCELL_X4 FILLER_121_1072 ();
 FILLCELL_X1 FILLER_121_1076 ();
 FILLCELL_X8 FILLER_121_1083 ();
 FILLCELL_X1 FILLER_121_1091 ();
 FILLCELL_X4 FILLER_121_1098 ();
 FILLCELL_X1 FILLER_121_1102 ();
 FILLCELL_X2 FILLER_121_1112 ();
 FILLCELL_X1 FILLER_121_1114 ();
 FILLCELL_X1 FILLER_121_1138 ();
 FILLCELL_X8 FILLER_121_1150 ();
 FILLCELL_X2 FILLER_121_1158 ();
 FILLCELL_X1 FILLER_121_1170 ();
 FILLCELL_X4 FILLER_121_1197 ();
 FILLCELL_X2 FILLER_121_1201 ();
 FILLCELL_X1 FILLER_121_1203 ();
 FILLCELL_X2 FILLER_121_1208 ();
 FILLCELL_X1 FILLER_121_1214 ();
 FILLCELL_X8 FILLER_121_1219 ();
 FILLCELL_X2 FILLER_121_1227 ();
 FILLCELL_X1 FILLER_121_1229 ();
 FILLCELL_X4 FILLER_121_1244 ();
 FILLCELL_X1 FILLER_121_1248 ();
 FILLCELL_X2 FILLER_121_1298 ();
 FILLCELL_X2 FILLER_121_1302 ();
 FILLCELL_X4 FILLER_121_1314 ();
 FILLCELL_X1 FILLER_121_1318 ();
 FILLCELL_X4 FILLER_121_1326 ();
 FILLCELL_X2 FILLER_121_1330 ();
 FILLCELL_X1 FILLER_121_1332 ();
 FILLCELL_X8 FILLER_121_1338 ();
 FILLCELL_X2 FILLER_121_1349 ();
 FILLCELL_X1 FILLER_121_1351 ();
 FILLCELL_X16 FILLER_121_1356 ();
 FILLCELL_X8 FILLER_121_1372 ();
 FILLCELL_X1 FILLER_121_1380 ();
 FILLCELL_X4 FILLER_121_1387 ();
 FILLCELL_X2 FILLER_121_1415 ();
 FILLCELL_X4 FILLER_121_1423 ();
 FILLCELL_X2 FILLER_121_1437 ();
 FILLCELL_X2 FILLER_121_1445 ();
 FILLCELL_X2 FILLER_121_1457 ();
 FILLCELL_X1 FILLER_121_1459 ();
 FILLCELL_X32 FILLER_121_1472 ();
 FILLCELL_X32 FILLER_121_1504 ();
 FILLCELL_X32 FILLER_121_1536 ();
 FILLCELL_X32 FILLER_121_1568 ();
 FILLCELL_X32 FILLER_121_1600 ();
 FILLCELL_X16 FILLER_121_1632 ();
 FILLCELL_X2 FILLER_121_1648 ();
 FILLCELL_X1 FILLER_121_1650 ();
 FILLCELL_X1 FILLER_122_21 ();
 FILLCELL_X1 FILLER_122_29 ();
 FILLCELL_X2 FILLER_122_50 ();
 FILLCELL_X2 FILLER_122_72 ();
 FILLCELL_X1 FILLER_122_74 ();
 FILLCELL_X2 FILLER_122_82 ();
 FILLCELL_X1 FILLER_122_84 ();
 FILLCELL_X4 FILLER_122_105 ();
 FILLCELL_X2 FILLER_122_109 ();
 FILLCELL_X1 FILLER_122_111 ();
 FILLCELL_X1 FILLER_122_130 ();
 FILLCELL_X1 FILLER_122_151 ();
 FILLCELL_X1 FILLER_122_172 ();
 FILLCELL_X2 FILLER_122_177 ();
 FILLCELL_X8 FILLER_122_203 ();
 FILLCELL_X2 FILLER_122_211 ();
 FILLCELL_X1 FILLER_122_213 ();
 FILLCELL_X1 FILLER_122_237 ();
 FILLCELL_X1 FILLER_122_242 ();
 FILLCELL_X2 FILLER_122_250 ();
 FILLCELL_X2 FILLER_122_281 ();
 FILLCELL_X1 FILLER_122_283 ();
 FILLCELL_X4 FILLER_122_288 ();
 FILLCELL_X1 FILLER_122_292 ();
 FILLCELL_X16 FILLER_122_325 ();
 FILLCELL_X4 FILLER_122_341 ();
 FILLCELL_X2 FILLER_122_345 ();
 FILLCELL_X2 FILLER_122_379 ();
 FILLCELL_X1 FILLER_122_381 ();
 FILLCELL_X1 FILLER_122_386 ();
 FILLCELL_X4 FILLER_122_410 ();
 FILLCELL_X4 FILLER_122_421 ();
 FILLCELL_X2 FILLER_122_425 ();
 FILLCELL_X1 FILLER_122_454 ();
 FILLCELL_X1 FILLER_122_462 ();
 FILLCELL_X4 FILLER_122_470 ();
 FILLCELL_X2 FILLER_122_474 ();
 FILLCELL_X1 FILLER_122_476 ();
 FILLCELL_X2 FILLER_122_500 ();
 FILLCELL_X1 FILLER_122_502 ();
 FILLCELL_X1 FILLER_122_523 ();
 FILLCELL_X1 FILLER_122_547 ();
 FILLCELL_X8 FILLER_122_552 ();
 FILLCELL_X1 FILLER_122_560 ();
 FILLCELL_X2 FILLER_122_581 ();
 FILLCELL_X8 FILLER_122_603 ();
 FILLCELL_X4 FILLER_122_636 ();
 FILLCELL_X8 FILLER_122_643 ();
 FILLCELL_X4 FILLER_122_651 ();
 FILLCELL_X2 FILLER_122_655 ();
 FILLCELL_X1 FILLER_122_657 ();
 FILLCELL_X1 FILLER_122_702 ();
 FILLCELL_X4 FILLER_122_713 ();
 FILLCELL_X1 FILLER_122_717 ();
 FILLCELL_X8 FILLER_122_738 ();
 FILLCELL_X2 FILLER_122_746 ();
 FILLCELL_X1 FILLER_122_748 ();
 FILLCELL_X8 FILLER_122_756 ();
 FILLCELL_X2 FILLER_122_764 ();
 FILLCELL_X1 FILLER_122_766 ();
 FILLCELL_X8 FILLER_122_770 ();
 FILLCELL_X2 FILLER_122_778 ();
 FILLCELL_X8 FILLER_122_800 ();
 FILLCELL_X4 FILLER_122_808 ();
 FILLCELL_X1 FILLER_122_812 ();
 FILLCELL_X2 FILLER_122_817 ();
 FILLCELL_X1 FILLER_122_819 ();
 FILLCELL_X2 FILLER_122_823 ();
 FILLCELL_X2 FILLER_122_829 ();
 FILLCELL_X4 FILLER_122_854 ();
 FILLCELL_X2 FILLER_122_858 ();
 FILLCELL_X4 FILLER_122_863 ();
 FILLCELL_X8 FILLER_122_894 ();
 FILLCELL_X4 FILLER_122_902 ();
 FILLCELL_X2 FILLER_122_906 ();
 FILLCELL_X1 FILLER_122_908 ();
 FILLCELL_X2 FILLER_122_914 ();
 FILLCELL_X1 FILLER_122_916 ();
 FILLCELL_X4 FILLER_122_924 ();
 FILLCELL_X1 FILLER_122_928 ();
 FILLCELL_X4 FILLER_122_935 ();
 FILLCELL_X1 FILLER_122_939 ();
 FILLCELL_X4 FILLER_122_960 ();
 FILLCELL_X4 FILLER_122_977 ();
 FILLCELL_X1 FILLER_122_981 ();
 FILLCELL_X4 FILLER_122_1024 ();
 FILLCELL_X16 FILLER_122_1055 ();
 FILLCELL_X1 FILLER_122_1071 ();
 FILLCELL_X2 FILLER_122_1082 ();
 FILLCELL_X2 FILLER_122_1090 ();
 FILLCELL_X1 FILLER_122_1092 ();
 FILLCELL_X2 FILLER_122_1115 ();
 FILLCELL_X1 FILLER_122_1117 ();
 FILLCELL_X2 FILLER_122_1124 ();
 FILLCELL_X1 FILLER_122_1141 ();
 FILLCELL_X1 FILLER_122_1146 ();
 FILLCELL_X1 FILLER_122_1169 ();
 FILLCELL_X1 FILLER_122_1176 ();
 FILLCELL_X2 FILLER_122_1181 ();
 FILLCELL_X2 FILLER_122_1203 ();
 FILLCELL_X1 FILLER_122_1205 ();
 FILLCELL_X1 FILLER_122_1244 ();
 FILLCELL_X1 FILLER_122_1256 ();
 FILLCELL_X1 FILLER_122_1262 ();
 FILLCELL_X1 FILLER_122_1265 ();
 FILLCELL_X2 FILLER_122_1270 ();
 FILLCELL_X1 FILLER_122_1282 ();
 FILLCELL_X8 FILLER_122_1289 ();
 FILLCELL_X4 FILLER_122_1297 ();
 FILLCELL_X1 FILLER_122_1301 ();
 FILLCELL_X2 FILLER_122_1327 ();
 FILLCELL_X1 FILLER_122_1329 ();
 FILLCELL_X4 FILLER_122_1332 ();
 FILLCELL_X2 FILLER_122_1336 ();
 FILLCELL_X4 FILLER_122_1342 ();
 FILLCELL_X4 FILLER_122_1350 ();
 FILLCELL_X1 FILLER_122_1354 ();
 FILLCELL_X2 FILLER_122_1359 ();
 FILLCELL_X1 FILLER_122_1361 ();
 FILLCELL_X4 FILLER_122_1378 ();
 FILLCELL_X2 FILLER_122_1382 ();
 FILLCELL_X2 FILLER_122_1424 ();
 FILLCELL_X1 FILLER_122_1426 ();
 FILLCELL_X4 FILLER_122_1433 ();
 FILLCELL_X2 FILLER_122_1437 ();
 FILLCELL_X2 FILLER_122_1449 ();
 FILLCELL_X1 FILLER_122_1451 ();
 FILLCELL_X32 FILLER_122_1478 ();
 FILLCELL_X32 FILLER_122_1510 ();
 FILLCELL_X32 FILLER_122_1542 ();
 FILLCELL_X32 FILLER_122_1574 ();
 FILLCELL_X32 FILLER_122_1606 ();
 FILLCELL_X8 FILLER_122_1638 ();
 FILLCELL_X4 FILLER_122_1646 ();
 FILLCELL_X1 FILLER_122_1650 ();
 FILLCELL_X1 FILLER_123_1 ();
 FILLCELL_X4 FILLER_123_34 ();
 FILLCELL_X2 FILLER_123_38 ();
 FILLCELL_X1 FILLER_123_40 ();
 FILLCELL_X2 FILLER_123_58 ();
 FILLCELL_X1 FILLER_123_60 ();
 FILLCELL_X8 FILLER_123_93 ();
 FILLCELL_X4 FILLER_123_101 ();
 FILLCELL_X2 FILLER_123_105 ();
 FILLCELL_X8 FILLER_123_116 ();
 FILLCELL_X4 FILLER_123_124 ();
 FILLCELL_X1 FILLER_123_128 ();
 FILLCELL_X2 FILLER_123_156 ();
 FILLCELL_X1 FILLER_123_158 ();
 FILLCELL_X32 FILLER_123_184 ();
 FILLCELL_X1 FILLER_123_216 ();
 FILLCELL_X1 FILLER_123_238 ();
 FILLCELL_X4 FILLER_123_248 ();
 FILLCELL_X8 FILLER_123_298 ();
 FILLCELL_X2 FILLER_123_306 ();
 FILLCELL_X1 FILLER_123_308 ();
 FILLCELL_X2 FILLER_123_313 ();
 FILLCELL_X2 FILLER_123_326 ();
 FILLCELL_X1 FILLER_123_328 ();
 FILLCELL_X2 FILLER_123_369 ();
 FILLCELL_X2 FILLER_123_376 ();
 FILLCELL_X8 FILLER_123_398 ();
 FILLCELL_X2 FILLER_123_436 ();
 FILLCELL_X1 FILLER_123_438 ();
 FILLCELL_X1 FILLER_123_506 ();
 FILLCELL_X32 FILLER_123_535 ();
 FILLCELL_X8 FILLER_123_567 ();
 FILLCELL_X4 FILLER_123_575 ();
 FILLCELL_X2 FILLER_123_579 ();
 FILLCELL_X4 FILLER_123_615 ();
 FILLCELL_X1 FILLER_123_619 ();
 FILLCELL_X2 FILLER_123_627 ();
 FILLCELL_X1 FILLER_123_629 ();
 FILLCELL_X4 FILLER_123_633 ();
 FILLCELL_X16 FILLER_123_644 ();
 FILLCELL_X4 FILLER_123_660 ();
 FILLCELL_X2 FILLER_123_664 ();
 FILLCELL_X8 FILLER_123_706 ();
 FILLCELL_X4 FILLER_123_717 ();
 FILLCELL_X2 FILLER_123_773 ();
 FILLCELL_X4 FILLER_123_786 ();
 FILLCELL_X1 FILLER_123_790 ();
 FILLCELL_X1 FILLER_123_814 ();
 FILLCELL_X1 FILLER_123_822 ();
 FILLCELL_X8 FILLER_123_827 ();
 FILLCELL_X4 FILLER_123_835 ();
 FILLCELL_X1 FILLER_123_839 ();
 FILLCELL_X1 FILLER_123_865 ();
 FILLCELL_X2 FILLER_123_874 ();
 FILLCELL_X2 FILLER_123_940 ();
 FILLCELL_X1 FILLER_123_949 ();
 FILLCELL_X16 FILLER_123_977 ();
 FILLCELL_X8 FILLER_123_993 ();
 FILLCELL_X1 FILLER_123_1001 ();
 FILLCELL_X1 FILLER_123_1026 ();
 FILLCELL_X8 FILLER_123_1037 ();
 FILLCELL_X16 FILLER_123_1067 ();
 FILLCELL_X4 FILLER_123_1083 ();
 FILLCELL_X1 FILLER_123_1087 ();
 FILLCELL_X8 FILLER_123_1114 ();
 FILLCELL_X1 FILLER_123_1122 ();
 FILLCELL_X1 FILLER_123_1129 ();
 FILLCELL_X2 FILLER_123_1136 ();
 FILLCELL_X2 FILLER_123_1148 ();
 FILLCELL_X8 FILLER_123_1168 ();
 FILLCELL_X4 FILLER_123_1186 ();
 FILLCELL_X1 FILLER_123_1190 ();
 FILLCELL_X1 FILLER_123_1198 ();
 FILLCELL_X4 FILLER_123_1211 ();
 FILLCELL_X16 FILLER_123_1222 ();
 FILLCELL_X1 FILLER_123_1238 ();
 FILLCELL_X4 FILLER_123_1242 ();
 FILLCELL_X2 FILLER_123_1246 ();
 FILLCELL_X1 FILLER_123_1248 ();
 FILLCELL_X4 FILLER_123_1253 ();
 FILLCELL_X2 FILLER_123_1264 ();
 FILLCELL_X1 FILLER_123_1306 ();
 FILLCELL_X1 FILLER_123_1321 ();
 FILLCELL_X1 FILLER_123_1344 ();
 FILLCELL_X4 FILLER_123_1373 ();
 FILLCELL_X1 FILLER_123_1377 ();
 FILLCELL_X4 FILLER_123_1384 ();
 FILLCELL_X2 FILLER_123_1406 ();
 FILLCELL_X1 FILLER_123_1408 ();
 FILLCELL_X2 FILLER_123_1419 ();
 FILLCELL_X1 FILLER_123_1441 ();
 FILLCELL_X1 FILLER_123_1452 ();
 FILLCELL_X1 FILLER_123_1459 ();
 FILLCELL_X32 FILLER_123_1466 ();
 FILLCELL_X32 FILLER_123_1498 ();
 FILLCELL_X32 FILLER_123_1530 ();
 FILLCELL_X32 FILLER_123_1562 ();
 FILLCELL_X32 FILLER_123_1594 ();
 FILLCELL_X16 FILLER_123_1626 ();
 FILLCELL_X8 FILLER_123_1642 ();
 FILLCELL_X1 FILLER_123_1650 ();
 FILLCELL_X16 FILLER_124_1 ();
 FILLCELL_X8 FILLER_124_17 ();
 FILLCELL_X4 FILLER_124_25 ();
 FILLCELL_X16 FILLER_124_34 ();
 FILLCELL_X8 FILLER_124_50 ();
 FILLCELL_X2 FILLER_124_78 ();
 FILLCELL_X1 FILLER_124_80 ();
 FILLCELL_X4 FILLER_124_101 ();
 FILLCELL_X2 FILLER_124_105 ();
 FILLCELL_X1 FILLER_124_107 ();
 FILLCELL_X1 FILLER_124_127 ();
 FILLCELL_X1 FILLER_124_162 ();
 FILLCELL_X2 FILLER_124_170 ();
 FILLCELL_X1 FILLER_124_179 ();
 FILLCELL_X4 FILLER_124_189 ();
 FILLCELL_X2 FILLER_124_193 ();
 FILLCELL_X1 FILLER_124_195 ();
 FILLCELL_X2 FILLER_124_200 ();
 FILLCELL_X1 FILLER_124_202 ();
 FILLCELL_X2 FILLER_124_230 ();
 FILLCELL_X4 FILLER_124_261 ();
 FILLCELL_X1 FILLER_124_265 ();
 FILLCELL_X2 FILLER_124_274 ();
 FILLCELL_X1 FILLER_124_276 ();
 FILLCELL_X8 FILLER_124_297 ();
 FILLCELL_X2 FILLER_124_305 ();
 FILLCELL_X4 FILLER_124_327 ();
 FILLCELL_X1 FILLER_124_331 ();
 FILLCELL_X4 FILLER_124_361 ();
 FILLCELL_X2 FILLER_124_365 ();
 FILLCELL_X1 FILLER_124_367 ();
 FILLCELL_X4 FILLER_124_383 ();
 FILLCELL_X2 FILLER_124_387 ();
 FILLCELL_X1 FILLER_124_389 ();
 FILLCELL_X4 FILLER_124_393 ();
 FILLCELL_X2 FILLER_124_397 ();
 FILLCELL_X1 FILLER_124_399 ();
 FILLCELL_X32 FILLER_124_443 ();
 FILLCELL_X2 FILLER_124_475 ();
 FILLCELL_X1 FILLER_124_492 ();
 FILLCELL_X1 FILLER_124_497 ();
 FILLCELL_X2 FILLER_124_505 ();
 FILLCELL_X1 FILLER_124_507 ();
 FILLCELL_X2 FILLER_124_535 ();
 FILLCELL_X1 FILLER_124_546 ();
 FILLCELL_X4 FILLER_124_572 ();
 FILLCELL_X1 FILLER_124_576 ();
 FILLCELL_X2 FILLER_124_600 ();
 FILLCELL_X1 FILLER_124_626 ();
 FILLCELL_X1 FILLER_124_632 ();
 FILLCELL_X1 FILLER_124_636 ();
 FILLCELL_X4 FILLER_124_669 ();
 FILLCELL_X1 FILLER_124_673 ();
 FILLCELL_X8 FILLER_124_678 ();
 FILLCELL_X1 FILLER_124_686 ();
 FILLCELL_X8 FILLER_124_691 ();
 FILLCELL_X4 FILLER_124_702 ();
 FILLCELL_X2 FILLER_124_706 ();
 FILLCELL_X1 FILLER_124_712 ();
 FILLCELL_X1 FILLER_124_717 ();
 FILLCELL_X8 FILLER_124_721 ();
 FILLCELL_X2 FILLER_124_729 ();
 FILLCELL_X1 FILLER_124_731 ();
 FILLCELL_X4 FILLER_124_744 ();
 FILLCELL_X1 FILLER_124_753 ();
 FILLCELL_X4 FILLER_124_781 ();
 FILLCELL_X8 FILLER_124_792 ();
 FILLCELL_X8 FILLER_124_809 ();
 FILLCELL_X2 FILLER_124_817 ();
 FILLCELL_X2 FILLER_124_842 ();
 FILLCELL_X1 FILLER_124_869 ();
 FILLCELL_X1 FILLER_124_910 ();
 FILLCELL_X1 FILLER_124_936 ();
 FILLCELL_X1 FILLER_124_944 ();
 FILLCELL_X8 FILLER_124_953 ();
 FILLCELL_X2 FILLER_124_961 ();
 FILLCELL_X32 FILLER_124_972 ();
 FILLCELL_X4 FILLER_124_1004 ();
 FILLCELL_X2 FILLER_124_1037 ();
 FILLCELL_X4 FILLER_124_1047 ();
 FILLCELL_X2 FILLER_124_1051 ();
 FILLCELL_X1 FILLER_124_1053 ();
 FILLCELL_X32 FILLER_124_1061 ();
 FILLCELL_X2 FILLER_124_1093 ();
 FILLCELL_X1 FILLER_124_1105 ();
 FILLCELL_X1 FILLER_124_1116 ();
 FILLCELL_X1 FILLER_124_1133 ();
 FILLCELL_X1 FILLER_124_1140 ();
 FILLCELL_X2 FILLER_124_1209 ();
 FILLCELL_X4 FILLER_124_1283 ();
 FILLCELL_X1 FILLER_124_1287 ();
 FILLCELL_X4 FILLER_124_1298 ();
 FILLCELL_X2 FILLER_124_1302 ();
 FILLCELL_X1 FILLER_124_1304 ();
 FILLCELL_X4 FILLER_124_1317 ();
 FILLCELL_X2 FILLER_124_1321 ();
 FILLCELL_X1 FILLER_124_1323 ();
 FILLCELL_X4 FILLER_124_1335 ();
 FILLCELL_X1 FILLER_124_1346 ();
 FILLCELL_X2 FILLER_124_1350 ();
 FILLCELL_X8 FILLER_124_1355 ();
 FILLCELL_X2 FILLER_124_1363 ();
 FILLCELL_X1 FILLER_124_1399 ();
 FILLCELL_X1 FILLER_124_1410 ();
 FILLCELL_X8 FILLER_124_1417 ();
 FILLCELL_X4 FILLER_124_1425 ();
 FILLCELL_X2 FILLER_124_1429 ();
 FILLCELL_X1 FILLER_124_1431 ();
 FILLCELL_X1 FILLER_124_1450 ();
 FILLCELL_X32 FILLER_124_1463 ();
 FILLCELL_X32 FILLER_124_1495 ();
 FILLCELL_X32 FILLER_124_1527 ();
 FILLCELL_X32 FILLER_124_1559 ();
 FILLCELL_X32 FILLER_124_1591 ();
 FILLCELL_X16 FILLER_124_1623 ();
 FILLCELL_X8 FILLER_124_1639 ();
 FILLCELL_X4 FILLER_124_1647 ();
 FILLCELL_X16 FILLER_125_1 ();
 FILLCELL_X8 FILLER_125_17 ();
 FILLCELL_X4 FILLER_125_25 ();
 FILLCELL_X2 FILLER_125_29 ();
 FILLCELL_X2 FILLER_125_62 ();
 FILLCELL_X2 FILLER_125_104 ();
 FILLCELL_X16 FILLER_125_120 ();
 FILLCELL_X4 FILLER_125_136 ();
 FILLCELL_X1 FILLER_125_140 ();
 FILLCELL_X1 FILLER_125_160 ();
 FILLCELL_X16 FILLER_125_205 ();
 FILLCELL_X2 FILLER_125_221 ();
 FILLCELL_X4 FILLER_125_230 ();
 FILLCELL_X1 FILLER_125_234 ();
 FILLCELL_X4 FILLER_125_260 ();
 FILLCELL_X2 FILLER_125_288 ();
 FILLCELL_X1 FILLER_125_310 ();
 FILLCELL_X8 FILLER_125_324 ();
 FILLCELL_X1 FILLER_125_339 ();
 FILLCELL_X16 FILLER_125_352 ();
 FILLCELL_X1 FILLER_125_368 ();
 FILLCELL_X2 FILLER_125_374 ();
 FILLCELL_X1 FILLER_125_376 ();
 FILLCELL_X4 FILLER_125_431 ();
 FILLCELL_X1 FILLER_125_435 ();
 FILLCELL_X1 FILLER_125_445 ();
 FILLCELL_X1 FILLER_125_460 ();
 FILLCELL_X2 FILLER_125_470 ();
 FILLCELL_X2 FILLER_125_492 ();
 FILLCELL_X4 FILLER_125_514 ();
 FILLCELL_X2 FILLER_125_518 ();
 FILLCELL_X2 FILLER_125_524 ();
 FILLCELL_X2 FILLER_125_546 ();
 FILLCELL_X1 FILLER_125_548 ();
 FILLCELL_X16 FILLER_125_556 ();
 FILLCELL_X1 FILLER_125_592 ();
 FILLCELL_X4 FILLER_125_616 ();
 FILLCELL_X1 FILLER_125_620 ();
 FILLCELL_X4 FILLER_125_641 ();
 FILLCELL_X2 FILLER_125_645 ();
 FILLCELL_X1 FILLER_125_647 ();
 FILLCELL_X2 FILLER_125_679 ();
 FILLCELL_X1 FILLER_125_681 ();
 FILLCELL_X2 FILLER_125_719 ();
 FILLCELL_X4 FILLER_125_758 ();
 FILLCELL_X1 FILLER_125_762 ();
 FILLCELL_X1 FILLER_125_804 ();
 FILLCELL_X8 FILLER_125_841 ();
 FILLCELL_X1 FILLER_125_849 ();
 FILLCELL_X2 FILLER_125_857 ();
 FILLCELL_X1 FILLER_125_859 ();
 FILLCELL_X4 FILLER_125_879 ();
 FILLCELL_X1 FILLER_125_883 ();
 FILLCELL_X2 FILLER_125_889 ();
 FILLCELL_X1 FILLER_125_891 ();
 FILLCELL_X4 FILLER_125_902 ();
 FILLCELL_X2 FILLER_125_906 ();
 FILLCELL_X1 FILLER_125_908 ();
 FILLCELL_X32 FILLER_125_929 ();
 FILLCELL_X2 FILLER_125_961 ();
 FILLCELL_X1 FILLER_125_963 ();
 FILLCELL_X8 FILLER_125_973 ();
 FILLCELL_X4 FILLER_125_981 ();
 FILLCELL_X2 FILLER_125_985 ();
 FILLCELL_X8 FILLER_125_1000 ();
 FILLCELL_X4 FILLER_125_1008 ();
 FILLCELL_X1 FILLER_125_1012 ();
 FILLCELL_X8 FILLER_125_1023 ();
 FILLCELL_X4 FILLER_125_1031 ();
 FILLCELL_X2 FILLER_125_1035 ();
 FILLCELL_X1 FILLER_125_1037 ();
 FILLCELL_X4 FILLER_125_1044 ();
 FILLCELL_X8 FILLER_125_1085 ();
 FILLCELL_X4 FILLER_125_1093 ();
 FILLCELL_X2 FILLER_125_1107 ();
 FILLCELL_X2 FILLER_125_1119 ();
 FILLCELL_X1 FILLER_125_1121 ();
 FILLCELL_X2 FILLER_125_1185 ();
 FILLCELL_X1 FILLER_125_1187 ();
 FILLCELL_X1 FILLER_125_1192 ();
 FILLCELL_X8 FILLER_125_1205 ();
 FILLCELL_X2 FILLER_125_1213 ();
 FILLCELL_X8 FILLER_125_1226 ();
 FILLCELL_X4 FILLER_125_1234 ();
 FILLCELL_X1 FILLER_125_1238 ();
 FILLCELL_X4 FILLER_125_1246 ();
 FILLCELL_X2 FILLER_125_1250 ();
 FILLCELL_X1 FILLER_125_1252 ();
 FILLCELL_X1 FILLER_125_1258 ();
 FILLCELL_X1 FILLER_125_1262 ();
 FILLCELL_X2 FILLER_125_1270 ();
 FILLCELL_X2 FILLER_125_1302 ();
 FILLCELL_X1 FILLER_125_1304 ();
 FILLCELL_X4 FILLER_125_1319 ();
 FILLCELL_X1 FILLER_125_1323 ();
 FILLCELL_X4 FILLER_125_1339 ();
 FILLCELL_X2 FILLER_125_1343 ();
 FILLCELL_X1 FILLER_125_1345 ();
 FILLCELL_X2 FILLER_125_1349 ();
 FILLCELL_X8 FILLER_125_1355 ();
 FILLCELL_X4 FILLER_125_1363 ();
 FILLCELL_X4 FILLER_125_1373 ();
 FILLCELL_X1 FILLER_125_1377 ();
 FILLCELL_X1 FILLER_125_1384 ();
 FILLCELL_X1 FILLER_125_1391 ();
 FILLCELL_X1 FILLER_125_1398 ();
 FILLCELL_X2 FILLER_125_1405 ();
 FILLCELL_X1 FILLER_125_1439 ();
 FILLCELL_X32 FILLER_125_1456 ();
 FILLCELL_X32 FILLER_125_1488 ();
 FILLCELL_X32 FILLER_125_1520 ();
 FILLCELL_X32 FILLER_125_1552 ();
 FILLCELL_X32 FILLER_125_1584 ();
 FILLCELL_X32 FILLER_125_1616 ();
 FILLCELL_X2 FILLER_125_1648 ();
 FILLCELL_X1 FILLER_125_1650 ();
 FILLCELL_X8 FILLER_126_1 ();
 FILLCELL_X1 FILLER_126_9 ();
 FILLCELL_X8 FILLER_126_37 ();
 FILLCELL_X4 FILLER_126_45 ();
 FILLCELL_X16 FILLER_126_54 ();
 FILLCELL_X2 FILLER_126_70 ();
 FILLCELL_X1 FILLER_126_72 ();
 FILLCELL_X1 FILLER_126_81 ();
 FILLCELL_X16 FILLER_126_89 ();
 FILLCELL_X4 FILLER_126_105 ();
 FILLCELL_X8 FILLER_126_129 ();
 FILLCELL_X1 FILLER_126_137 ();
 FILLCELL_X4 FILLER_126_158 ();
 FILLCELL_X2 FILLER_126_162 ();
 FILLCELL_X4 FILLER_126_171 ();
 FILLCELL_X2 FILLER_126_175 ();
 FILLCELL_X4 FILLER_126_190 ();
 FILLCELL_X8 FILLER_126_203 ();
 FILLCELL_X4 FILLER_126_211 ();
 FILLCELL_X2 FILLER_126_258 ();
 FILLCELL_X1 FILLER_126_260 ();
 FILLCELL_X4 FILLER_126_265 ();
 FILLCELL_X4 FILLER_126_272 ();
 FILLCELL_X8 FILLER_126_279 ();
 FILLCELL_X4 FILLER_126_327 ();
 FILLCELL_X2 FILLER_126_354 ();
 FILLCELL_X2 FILLER_126_361 ();
 FILLCELL_X2 FILLER_126_391 ();
 FILLCELL_X1 FILLER_126_393 ();
 FILLCELL_X2 FILLER_126_431 ();
 FILLCELL_X8 FILLER_126_465 ();
 FILLCELL_X2 FILLER_126_473 ();
 FILLCELL_X1 FILLER_126_475 ();
 FILLCELL_X4 FILLER_126_480 ();
 FILLCELL_X1 FILLER_126_484 ();
 FILLCELL_X4 FILLER_126_508 ();
 FILLCELL_X1 FILLER_126_512 ();
 FILLCELL_X8 FILLER_126_515 ();
 FILLCELL_X4 FILLER_126_523 ();
 FILLCELL_X2 FILLER_126_527 ();
 FILLCELL_X8 FILLER_126_536 ();
 FILLCELL_X2 FILLER_126_544 ();
 FILLCELL_X4 FILLER_126_591 ();
 FILLCELL_X8 FILLER_126_620 ();
 FILLCELL_X2 FILLER_126_628 ();
 FILLCELL_X1 FILLER_126_630 ();
 FILLCELL_X2 FILLER_126_632 ();
 FILLCELL_X1 FILLER_126_634 ();
 FILLCELL_X2 FILLER_126_656 ();
 FILLCELL_X2 FILLER_126_661 ();
 FILLCELL_X1 FILLER_126_663 ();
 FILLCELL_X8 FILLER_126_684 ();
 FILLCELL_X2 FILLER_126_692 ();
 FILLCELL_X1 FILLER_126_694 ();
 FILLCELL_X2 FILLER_126_708 ();
 FILLCELL_X2 FILLER_126_721 ();
 FILLCELL_X1 FILLER_126_730 ();
 FILLCELL_X2 FILLER_126_734 ();
 FILLCELL_X1 FILLER_126_736 ();
 FILLCELL_X2 FILLER_126_755 ();
 FILLCELL_X1 FILLER_126_757 ();
 FILLCELL_X8 FILLER_126_765 ();
 FILLCELL_X2 FILLER_126_793 ();
 FILLCELL_X1 FILLER_126_795 ();
 FILLCELL_X16 FILLER_126_823 ();
 FILLCELL_X8 FILLER_126_839 ();
 FILLCELL_X2 FILLER_126_847 ();
 FILLCELL_X1 FILLER_126_849 ();
 FILLCELL_X2 FILLER_126_888 ();
 FILLCELL_X4 FILLER_126_915 ();
 FILLCELL_X2 FILLER_126_919 ();
 FILLCELL_X1 FILLER_126_928 ();
 FILLCELL_X4 FILLER_126_961 ();
 FILLCELL_X8 FILLER_126_981 ();
 FILLCELL_X1 FILLER_126_989 ();
 FILLCELL_X8 FILLER_126_999 ();
 FILLCELL_X2 FILLER_126_1007 ();
 FILLCELL_X1 FILLER_126_1009 ();
 FILLCELL_X16 FILLER_126_1024 ();
 FILLCELL_X8 FILLER_126_1043 ();
 FILLCELL_X2 FILLER_126_1051 ();
 FILLCELL_X1 FILLER_126_1053 ();
 FILLCELL_X16 FILLER_126_1061 ();
 FILLCELL_X4 FILLER_126_1077 ();
 FILLCELL_X2 FILLER_126_1081 ();
 FILLCELL_X4 FILLER_126_1105 ();
 FILLCELL_X2 FILLER_126_1109 ();
 FILLCELL_X1 FILLER_126_1117 ();
 FILLCELL_X2 FILLER_126_1148 ();
 FILLCELL_X4 FILLER_126_1153 ();
 FILLCELL_X2 FILLER_126_1160 ();
 FILLCELL_X4 FILLER_126_1167 ();
 FILLCELL_X4 FILLER_126_1187 ();
 FILLCELL_X16 FILLER_126_1196 ();
 FILLCELL_X2 FILLER_126_1212 ();
 FILLCELL_X1 FILLER_126_1214 ();
 FILLCELL_X4 FILLER_126_1222 ();
 FILLCELL_X2 FILLER_126_1226 ();
 FILLCELL_X1 FILLER_126_1228 ();
 FILLCELL_X4 FILLER_126_1254 ();
 FILLCELL_X8 FILLER_126_1270 ();
 FILLCELL_X2 FILLER_126_1278 ();
 FILLCELL_X16 FILLER_126_1287 ();
 FILLCELL_X2 FILLER_126_1303 ();
 FILLCELL_X8 FILLER_126_1319 ();
 FILLCELL_X4 FILLER_126_1327 ();
 FILLCELL_X1 FILLER_126_1331 ();
 FILLCELL_X8 FILLER_126_1337 ();
 FILLCELL_X4 FILLER_126_1345 ();
 FILLCELL_X2 FILLER_126_1349 ();
 FILLCELL_X8 FILLER_126_1373 ();
 FILLCELL_X4 FILLER_126_1381 ();
 FILLCELL_X1 FILLER_126_1385 ();
 FILLCELL_X2 FILLER_126_1408 ();
 FILLCELL_X4 FILLER_126_1416 ();
 FILLCELL_X2 FILLER_126_1420 ();
 FILLCELL_X2 FILLER_126_1428 ();
 FILLCELL_X1 FILLER_126_1436 ();
 FILLCELL_X32 FILLER_126_1443 ();
 FILLCELL_X32 FILLER_126_1475 ();
 FILLCELL_X32 FILLER_126_1507 ();
 FILLCELL_X32 FILLER_126_1539 ();
 FILLCELL_X32 FILLER_126_1571 ();
 FILLCELL_X32 FILLER_126_1603 ();
 FILLCELL_X16 FILLER_126_1635 ();
 FILLCELL_X16 FILLER_127_1 ();
 FILLCELL_X1 FILLER_127_17 ();
 FILLCELL_X4 FILLER_127_23 ();
 FILLCELL_X2 FILLER_127_27 ();
 FILLCELL_X1 FILLER_127_29 ();
 FILLCELL_X4 FILLER_127_57 ();
 FILLCELL_X2 FILLER_127_61 ();
 FILLCELL_X8 FILLER_127_110 ();
 FILLCELL_X4 FILLER_127_118 ();
 FILLCELL_X16 FILLER_127_127 ();
 FILLCELL_X2 FILLER_127_143 ();
 FILLCELL_X1 FILLER_127_145 ();
 FILLCELL_X8 FILLER_127_159 ();
 FILLCELL_X4 FILLER_127_167 ();
 FILLCELL_X2 FILLER_127_171 ();
 FILLCELL_X1 FILLER_127_173 ();
 FILLCELL_X8 FILLER_127_214 ();
 FILLCELL_X4 FILLER_127_222 ();
 FILLCELL_X2 FILLER_127_226 ();
 FILLCELL_X1 FILLER_127_228 ();
 FILLCELL_X8 FILLER_127_233 ();
 FILLCELL_X2 FILLER_127_241 ();
 FILLCELL_X1 FILLER_127_243 ();
 FILLCELL_X8 FILLER_127_280 ();
 FILLCELL_X4 FILLER_127_288 ();
 FILLCELL_X1 FILLER_127_315 ();
 FILLCELL_X8 FILLER_127_327 ();
 FILLCELL_X1 FILLER_127_335 ();
 FILLCELL_X1 FILLER_127_363 ();
 FILLCELL_X1 FILLER_127_369 ();
 FILLCELL_X4 FILLER_127_374 ();
 FILLCELL_X1 FILLER_127_378 ();
 FILLCELL_X1 FILLER_127_382 ();
 FILLCELL_X8 FILLER_127_392 ();
 FILLCELL_X4 FILLER_127_400 ();
 FILLCELL_X2 FILLER_127_411 ();
 FILLCELL_X16 FILLER_127_429 ();
 FILLCELL_X4 FILLER_127_445 ();
 FILLCELL_X1 FILLER_127_449 ();
 FILLCELL_X4 FILLER_127_462 ();
 FILLCELL_X2 FILLER_127_466 ();
 FILLCELL_X1 FILLER_127_492 ();
 FILLCELL_X1 FILLER_127_501 ();
 FILLCELL_X2 FILLER_127_539 ();
 FILLCELL_X8 FILLER_127_561 ();
 FILLCELL_X2 FILLER_127_577 ();
 FILLCELL_X1 FILLER_127_579 ();
 FILLCELL_X2 FILLER_127_583 ();
 FILLCELL_X1 FILLER_127_590 ();
 FILLCELL_X2 FILLER_127_597 ();
 FILLCELL_X2 FILLER_127_603 ();
 FILLCELL_X1 FILLER_127_605 ();
 FILLCELL_X8 FILLER_127_613 ();
 FILLCELL_X2 FILLER_127_621 ();
 FILLCELL_X1 FILLER_127_623 ();
 FILLCELL_X1 FILLER_127_664 ();
 FILLCELL_X1 FILLER_127_669 ();
 FILLCELL_X4 FILLER_127_677 ();
 FILLCELL_X2 FILLER_127_749 ();
 FILLCELL_X2 FILLER_127_771 ();
 FILLCELL_X1 FILLER_127_773 ();
 FILLCELL_X2 FILLER_127_781 ();
 FILLCELL_X1 FILLER_127_783 ();
 FILLCELL_X2 FILLER_127_791 ();
 FILLCELL_X1 FILLER_127_793 ();
 FILLCELL_X32 FILLER_127_806 ();
 FILLCELL_X16 FILLER_127_838 ();
 FILLCELL_X4 FILLER_127_900 ();
 FILLCELL_X2 FILLER_127_904 ();
 FILLCELL_X1 FILLER_127_906 ();
 FILLCELL_X1 FILLER_127_914 ();
 FILLCELL_X8 FILLER_127_996 ();
 FILLCELL_X4 FILLER_127_1004 ();
 FILLCELL_X2 FILLER_127_1008 ();
 FILLCELL_X2 FILLER_127_1032 ();
 FILLCELL_X4 FILLER_127_1049 ();
 FILLCELL_X1 FILLER_127_1053 ();
 FILLCELL_X1 FILLER_127_1086 ();
 FILLCELL_X4 FILLER_127_1097 ();
 FILLCELL_X2 FILLER_127_1101 ();
 FILLCELL_X1 FILLER_127_1103 ();
 FILLCELL_X1 FILLER_127_1110 ();
 FILLCELL_X2 FILLER_127_1123 ();
 FILLCELL_X1 FILLER_127_1125 ();
 FILLCELL_X16 FILLER_127_1144 ();
 FILLCELL_X4 FILLER_127_1160 ();
 FILLCELL_X1 FILLER_127_1164 ();
 FILLCELL_X1 FILLER_127_1170 ();
 FILLCELL_X4 FILLER_127_1222 ();
 FILLCELL_X1 FILLER_127_1226 ();
 FILLCELL_X4 FILLER_127_1234 ();
 FILLCELL_X1 FILLER_127_1238 ();
 FILLCELL_X1 FILLER_127_1264 ();
 FILLCELL_X1 FILLER_127_1292 ();
 FILLCELL_X1 FILLER_127_1350 ();
 FILLCELL_X32 FILLER_127_1383 ();
 FILLCELL_X2 FILLER_127_1415 ();
 FILLCELL_X1 FILLER_127_1417 ();
 FILLCELL_X1 FILLER_127_1424 ();
 FILLCELL_X32 FILLER_127_1441 ();
 FILLCELL_X32 FILLER_127_1473 ();
 FILLCELL_X32 FILLER_127_1505 ();
 FILLCELL_X32 FILLER_127_1537 ();
 FILLCELL_X32 FILLER_127_1569 ();
 FILLCELL_X32 FILLER_127_1601 ();
 FILLCELL_X16 FILLER_127_1633 ();
 FILLCELL_X2 FILLER_127_1649 ();
 FILLCELL_X8 FILLER_128_1 ();
 FILLCELL_X2 FILLER_128_9 ();
 FILLCELL_X1 FILLER_128_11 ();
 FILLCELL_X4 FILLER_128_42 ();
 FILLCELL_X2 FILLER_128_57 ();
 FILLCELL_X2 FILLER_128_88 ();
 FILLCELL_X1 FILLER_128_90 ();
 FILLCELL_X4 FILLER_128_98 ();
 FILLCELL_X1 FILLER_128_102 ();
 FILLCELL_X4 FILLER_128_110 ();
 FILLCELL_X1 FILLER_128_119 ();
 FILLCELL_X8 FILLER_128_139 ();
 FILLCELL_X1 FILLER_128_147 ();
 FILLCELL_X4 FILLER_128_168 ();
 FILLCELL_X1 FILLER_128_172 ();
 FILLCELL_X4 FILLER_128_184 ();
 FILLCELL_X4 FILLER_128_200 ();
 FILLCELL_X1 FILLER_128_204 ();
 FILLCELL_X8 FILLER_128_235 ();
 FILLCELL_X2 FILLER_128_243 ();
 FILLCELL_X4 FILLER_128_277 ();
 FILLCELL_X1 FILLER_128_281 ();
 FILLCELL_X2 FILLER_128_286 ();
 FILLCELL_X1 FILLER_128_288 ();
 FILLCELL_X4 FILLER_128_292 ();
 FILLCELL_X1 FILLER_128_296 ();
 FILLCELL_X4 FILLER_128_306 ();
 FILLCELL_X1 FILLER_128_310 ();
 FILLCELL_X4 FILLER_128_323 ();
 FILLCELL_X1 FILLER_128_327 ();
 FILLCELL_X1 FILLER_128_348 ();
 FILLCELL_X4 FILLER_128_369 ();
 FILLCELL_X2 FILLER_128_373 ();
 FILLCELL_X1 FILLER_128_375 ();
 FILLCELL_X16 FILLER_128_388 ();
 FILLCELL_X4 FILLER_128_404 ();
 FILLCELL_X2 FILLER_128_408 ();
 FILLCELL_X8 FILLER_128_430 ();
 FILLCELL_X2 FILLER_128_438 ();
 FILLCELL_X1 FILLER_128_440 ();
 FILLCELL_X1 FILLER_128_461 ();
 FILLCELL_X1 FILLER_128_467 ();
 FILLCELL_X2 FILLER_128_488 ();
 FILLCELL_X8 FILLER_128_493 ();
 FILLCELL_X8 FILLER_128_504 ();
 FILLCELL_X4 FILLER_128_512 ();
 FILLCELL_X2 FILLER_128_516 ();
 FILLCELL_X1 FILLER_128_518 ();
 FILLCELL_X4 FILLER_128_539 ();
 FILLCELL_X2 FILLER_128_543 ();
 FILLCELL_X1 FILLER_128_545 ();
 FILLCELL_X4 FILLER_128_560 ();
 FILLCELL_X1 FILLER_128_604 ();
 FILLCELL_X2 FILLER_128_625 ();
 FILLCELL_X8 FILLER_128_661 ();
 FILLCELL_X4 FILLER_128_669 ();
 FILLCELL_X8 FILLER_128_693 ();
 FILLCELL_X2 FILLER_128_701 ();
 FILLCELL_X1 FILLER_128_703 ();
 FILLCELL_X2 FILLER_128_724 ();
 FILLCELL_X8 FILLER_128_733 ();
 FILLCELL_X4 FILLER_128_741 ();
 FILLCELL_X1 FILLER_128_745 ();
 FILLCELL_X16 FILLER_128_768 ();
 FILLCELL_X2 FILLER_128_784 ();
 FILLCELL_X8 FILLER_128_833 ();
 FILLCELL_X2 FILLER_128_841 ();
 FILLCELL_X1 FILLER_128_843 ();
 FILLCELL_X8 FILLER_128_871 ();
 FILLCELL_X2 FILLER_128_906 ();
 FILLCELL_X2 FILLER_128_928 ();
 FILLCELL_X1 FILLER_128_930 ();
 FILLCELL_X2 FILLER_128_936 ();
 FILLCELL_X1 FILLER_128_938 ();
 FILLCELL_X8 FILLER_128_966 ();
 FILLCELL_X2 FILLER_128_974 ();
 FILLCELL_X8 FILLER_128_1003 ();
 FILLCELL_X4 FILLER_128_1011 ();
 FILLCELL_X1 FILLER_128_1015 ();
 FILLCELL_X1 FILLER_128_1036 ();
 FILLCELL_X1 FILLER_128_1046 ();
 FILLCELL_X2 FILLER_128_1054 ();
 FILLCELL_X1 FILLER_128_1056 ();
 FILLCELL_X4 FILLER_128_1063 ();
 FILLCELL_X2 FILLER_128_1067 ();
 FILLCELL_X1 FILLER_128_1069 ();
 FILLCELL_X4 FILLER_128_1088 ();
 FILLCELL_X1 FILLER_128_1092 ();
 FILLCELL_X4 FILLER_128_1111 ();
 FILLCELL_X1 FILLER_128_1115 ();
 FILLCELL_X1 FILLER_128_1126 ();
 FILLCELL_X4 FILLER_128_1139 ();
 FILLCELL_X1 FILLER_128_1143 ();
 FILLCELL_X8 FILLER_128_1159 ();
 FILLCELL_X2 FILLER_128_1167 ();
 FILLCELL_X4 FILLER_128_1181 ();
 FILLCELL_X1 FILLER_128_1202 ();
 FILLCELL_X4 FILLER_128_1208 ();
 FILLCELL_X2 FILLER_128_1212 ();
 FILLCELL_X4 FILLER_128_1218 ();
 FILLCELL_X4 FILLER_128_1229 ();
 FILLCELL_X1 FILLER_128_1233 ();
 FILLCELL_X8 FILLER_128_1248 ();
 FILLCELL_X4 FILLER_128_1256 ();
 FILLCELL_X2 FILLER_128_1260 ();
 FILLCELL_X4 FILLER_128_1265 ();
 FILLCELL_X8 FILLER_128_1276 ();
 FILLCELL_X4 FILLER_128_1284 ();
 FILLCELL_X1 FILLER_128_1288 ();
 FILLCELL_X4 FILLER_128_1296 ();
 FILLCELL_X1 FILLER_128_1339 ();
 FILLCELL_X2 FILLER_128_1343 ();
 FILLCELL_X2 FILLER_128_1349 ();
 FILLCELL_X1 FILLER_128_1351 ();
 FILLCELL_X2 FILLER_128_1359 ();
 FILLCELL_X16 FILLER_128_1368 ();
 FILLCELL_X8 FILLER_128_1384 ();
 FILLCELL_X4 FILLER_128_1392 ();
 FILLCELL_X2 FILLER_128_1396 ();
 FILLCELL_X1 FILLER_128_1398 ();
 FILLCELL_X4 FILLER_128_1403 ();
 FILLCELL_X1 FILLER_128_1407 ();
 FILLCELL_X32 FILLER_128_1415 ();
 FILLCELL_X32 FILLER_128_1447 ();
 FILLCELL_X32 FILLER_128_1479 ();
 FILLCELL_X32 FILLER_128_1511 ();
 FILLCELL_X32 FILLER_128_1543 ();
 FILLCELL_X32 FILLER_128_1575 ();
 FILLCELL_X32 FILLER_128_1607 ();
 FILLCELL_X8 FILLER_128_1639 ();
 FILLCELL_X4 FILLER_128_1647 ();
 FILLCELL_X2 FILLER_129_1 ();
 FILLCELL_X1 FILLER_129_3 ();
 FILLCELL_X1 FILLER_129_24 ();
 FILLCELL_X1 FILLER_129_32 ();
 FILLCELL_X1 FILLER_129_38 ();
 FILLCELL_X8 FILLER_129_68 ();
 FILLCELL_X1 FILLER_129_76 ();
 FILLCELL_X2 FILLER_129_120 ();
 FILLCELL_X8 FILLER_129_135 ();
 FILLCELL_X4 FILLER_129_143 ();
 FILLCELL_X2 FILLER_129_147 ();
 FILLCELL_X2 FILLER_129_210 ();
 FILLCELL_X1 FILLER_129_212 ();
 FILLCELL_X1 FILLER_129_236 ();
 FILLCELL_X4 FILLER_129_254 ();
 FILLCELL_X8 FILLER_129_268 ();
 FILLCELL_X4 FILLER_129_276 ();
 FILLCELL_X1 FILLER_129_280 ();
 FILLCELL_X4 FILLER_129_301 ();
 FILLCELL_X1 FILLER_129_305 ();
 FILLCELL_X8 FILLER_129_326 ();
 FILLCELL_X2 FILLER_129_334 ();
 FILLCELL_X4 FILLER_129_343 ();
 FILLCELL_X2 FILLER_129_355 ();
 FILLCELL_X2 FILLER_129_360 ();
 FILLCELL_X1 FILLER_129_362 ();
 FILLCELL_X4 FILLER_129_366 ();
 FILLCELL_X2 FILLER_129_370 ();
 FILLCELL_X16 FILLER_129_392 ();
 FILLCELL_X4 FILLER_129_408 ();
 FILLCELL_X1 FILLER_129_412 ();
 FILLCELL_X8 FILLER_129_433 ();
 FILLCELL_X2 FILLER_129_441 ();
 FILLCELL_X1 FILLER_129_443 ();
 FILLCELL_X4 FILLER_129_460 ();
 FILLCELL_X4 FILLER_129_491 ();
 FILLCELL_X8 FILLER_129_499 ();
 FILLCELL_X8 FILLER_129_510 ();
 FILLCELL_X1 FILLER_129_530 ();
 FILLCELL_X2 FILLER_129_536 ();
 FILLCELL_X2 FILLER_129_545 ();
 FILLCELL_X1 FILLER_129_551 ();
 FILLCELL_X2 FILLER_129_562 ();
 FILLCELL_X2 FILLER_129_587 ();
 FILLCELL_X2 FILLER_129_593 ();
 FILLCELL_X8 FILLER_129_598 ();
 FILLCELL_X2 FILLER_129_606 ();
 FILLCELL_X4 FILLER_129_615 ();
 FILLCELL_X2 FILLER_129_619 ();
 FILLCELL_X4 FILLER_129_641 ();
 FILLCELL_X2 FILLER_129_645 ();
 FILLCELL_X4 FILLER_129_667 ();
 FILLCELL_X1 FILLER_129_671 ();
 FILLCELL_X4 FILLER_129_692 ();
 FILLCELL_X8 FILLER_129_715 ();
 FILLCELL_X4 FILLER_129_723 ();
 FILLCELL_X1 FILLER_129_727 ();
 FILLCELL_X2 FILLER_129_748 ();
 FILLCELL_X1 FILLER_129_757 ();
 FILLCELL_X2 FILLER_129_778 ();
 FILLCELL_X1 FILLER_129_787 ();
 FILLCELL_X4 FILLER_129_795 ();
 FILLCELL_X1 FILLER_129_799 ();
 FILLCELL_X1 FILLER_129_825 ();
 FILLCELL_X4 FILLER_129_833 ();
 FILLCELL_X2 FILLER_129_837 ();
 FILLCELL_X2 FILLER_129_863 ();
 FILLCELL_X2 FILLER_129_872 ();
 FILLCELL_X4 FILLER_129_887 ();
 FILLCELL_X1 FILLER_129_911 ();
 FILLCELL_X2 FILLER_129_919 ();
 FILLCELL_X1 FILLER_129_928 ();
 FILLCELL_X2 FILLER_129_932 ();
 FILLCELL_X8 FILLER_129_941 ();
 FILLCELL_X2 FILLER_129_949 ();
 FILLCELL_X1 FILLER_129_951 ();
 FILLCELL_X16 FILLER_129_959 ();
 FILLCELL_X2 FILLER_129_975 ();
 FILLCELL_X4 FILLER_129_982 ();
 FILLCELL_X2 FILLER_129_986 ();
 FILLCELL_X16 FILLER_129_1008 ();
 FILLCELL_X4 FILLER_129_1024 ();
 FILLCELL_X2 FILLER_129_1028 ();
 FILLCELL_X1 FILLER_129_1030 ();
 FILLCELL_X32 FILLER_129_1033 ();
 FILLCELL_X16 FILLER_129_1065 ();
 FILLCELL_X2 FILLER_129_1090 ();
 FILLCELL_X4 FILLER_129_1104 ();
 FILLCELL_X1 FILLER_129_1124 ();
 FILLCELL_X1 FILLER_129_1137 ();
 FILLCELL_X16 FILLER_129_1144 ();
 FILLCELL_X4 FILLER_129_1160 ();
 FILLCELL_X2 FILLER_129_1164 ();
 FILLCELL_X4 FILLER_129_1176 ();
 FILLCELL_X8 FILLER_129_1189 ();
 FILLCELL_X2 FILLER_129_1197 ();
 FILLCELL_X4 FILLER_129_1221 ();
 FILLCELL_X2 FILLER_129_1225 ();
 FILLCELL_X4 FILLER_129_1233 ();
 FILLCELL_X4 FILLER_129_1257 ();
 FILLCELL_X2 FILLER_129_1261 ();
 FILLCELL_X1 FILLER_129_1264 ();
 FILLCELL_X4 FILLER_129_1275 ();
 FILLCELL_X8 FILLER_129_1284 ();
 FILLCELL_X2 FILLER_129_1300 ();
 FILLCELL_X1 FILLER_129_1309 ();
 FILLCELL_X2 FILLER_129_1341 ();
 FILLCELL_X8 FILLER_129_1365 ();
 FILLCELL_X4 FILLER_129_1373 ();
 FILLCELL_X4 FILLER_129_1387 ();
 FILLCELL_X2 FILLER_129_1416 ();
 FILLCELL_X8 FILLER_129_1427 ();
 FILLCELL_X1 FILLER_129_1435 ();
 FILLCELL_X32 FILLER_129_1443 ();
 FILLCELL_X32 FILLER_129_1475 ();
 FILLCELL_X32 FILLER_129_1507 ();
 FILLCELL_X32 FILLER_129_1539 ();
 FILLCELL_X32 FILLER_129_1571 ();
 FILLCELL_X32 FILLER_129_1603 ();
 FILLCELL_X16 FILLER_129_1635 ();
 FILLCELL_X1 FILLER_130_1 ();
 FILLCELL_X2 FILLER_130_29 ();
 FILLCELL_X4 FILLER_130_54 ();
 FILLCELL_X1 FILLER_130_58 ();
 FILLCELL_X8 FILLER_130_66 ();
 FILLCELL_X2 FILLER_130_74 ();
 FILLCELL_X8 FILLER_130_85 ();
 FILLCELL_X4 FILLER_130_93 ();
 FILLCELL_X2 FILLER_130_104 ();
 FILLCELL_X1 FILLER_130_106 ();
 FILLCELL_X8 FILLER_130_119 ();
 FILLCELL_X4 FILLER_130_127 ();
 FILLCELL_X16 FILLER_130_157 ();
 FILLCELL_X4 FILLER_130_173 ();
 FILLCELL_X8 FILLER_130_202 ();
 FILLCELL_X4 FILLER_130_210 ();
 FILLCELL_X4 FILLER_130_227 ();
 FILLCELL_X1 FILLER_130_231 ();
 FILLCELL_X2 FILLER_130_252 ();
 FILLCELL_X16 FILLER_130_301 ();
 FILLCELL_X4 FILLER_130_317 ();
 FILLCELL_X2 FILLER_130_321 ();
 FILLCELL_X8 FILLER_130_343 ();
 FILLCELL_X4 FILLER_130_351 ();
 FILLCELL_X1 FILLER_130_355 ();
 FILLCELL_X8 FILLER_130_407 ();
 FILLCELL_X2 FILLER_130_415 ();
 FILLCELL_X4 FILLER_130_424 ();
 FILLCELL_X1 FILLER_130_435 ();
 FILLCELL_X2 FILLER_130_465 ();
 FILLCELL_X1 FILLER_130_467 ();
 FILLCELL_X8 FILLER_130_475 ();
 FILLCELL_X4 FILLER_130_483 ();
 FILLCELL_X2 FILLER_130_487 ();
 FILLCELL_X1 FILLER_130_489 ();
 FILLCELL_X1 FILLER_130_522 ();
 FILLCELL_X2 FILLER_130_531 ();
 FILLCELL_X1 FILLER_130_533 ();
 FILLCELL_X8 FILLER_130_560 ();
 FILLCELL_X2 FILLER_130_568 ();
 FILLCELL_X4 FILLER_130_574 ();
 FILLCELL_X1 FILLER_130_578 ();
 FILLCELL_X4 FILLER_130_582 ();
 FILLCELL_X2 FILLER_130_586 ();
 FILLCELL_X1 FILLER_130_588 ();
 FILLCELL_X8 FILLER_130_623 ();
 FILLCELL_X8 FILLER_130_639 ();
 FILLCELL_X2 FILLER_130_647 ();
 FILLCELL_X1 FILLER_130_663 ();
 FILLCELL_X2 FILLER_130_677 ();
 FILLCELL_X2 FILLER_130_699 ();
 FILLCELL_X1 FILLER_130_701 ();
 FILLCELL_X16 FILLER_130_722 ();
 FILLCELL_X8 FILLER_130_738 ();
 FILLCELL_X2 FILLER_130_746 ();
 FILLCELL_X16 FILLER_130_768 ();
 FILLCELL_X4 FILLER_130_784 ();
 FILLCELL_X1 FILLER_130_788 ();
 FILLCELL_X2 FILLER_130_814 ();
 FILLCELL_X1 FILLER_130_827 ();
 FILLCELL_X4 FILLER_130_848 ();
 FILLCELL_X2 FILLER_130_852 ();
 FILLCELL_X8 FILLER_130_881 ();
 FILLCELL_X1 FILLER_130_909 ();
 FILLCELL_X1 FILLER_130_927 ();
 FILLCELL_X2 FILLER_130_932 ();
 FILLCELL_X1 FILLER_130_934 ();
 FILLCELL_X2 FILLER_130_955 ();
 FILLCELL_X4 FILLER_130_1003 ();
 FILLCELL_X1 FILLER_130_1007 ();
 FILLCELL_X8 FILLER_130_1021 ();
 FILLCELL_X4 FILLER_130_1036 ();
 FILLCELL_X8 FILLER_130_1060 ();
 FILLCELL_X4 FILLER_130_1068 ();
 FILLCELL_X2 FILLER_130_1072 ();
 FILLCELL_X1 FILLER_130_1100 ();
 FILLCELL_X4 FILLER_130_1107 ();
 FILLCELL_X2 FILLER_130_1137 ();
 FILLCELL_X1 FILLER_130_1149 ();
 FILLCELL_X4 FILLER_130_1156 ();
 FILLCELL_X4 FILLER_130_1176 ();
 FILLCELL_X16 FILLER_130_1196 ();
 FILLCELL_X16 FILLER_130_1260 ();
 FILLCELL_X2 FILLER_130_1276 ();
 FILLCELL_X1 FILLER_130_1278 ();
 FILLCELL_X8 FILLER_130_1299 ();
 FILLCELL_X2 FILLER_130_1311 ();
 FILLCELL_X1 FILLER_130_1313 ();
 FILLCELL_X8 FILLER_130_1317 ();
 FILLCELL_X1 FILLER_130_1325 ();
 FILLCELL_X1 FILLER_130_1351 ();
 FILLCELL_X4 FILLER_130_1374 ();
 FILLCELL_X1 FILLER_130_1391 ();
 FILLCELL_X1 FILLER_130_1406 ();
 FILLCELL_X1 FILLER_130_1416 ();
 FILLCELL_X8 FILLER_130_1424 ();
 FILLCELL_X4 FILLER_130_1432 ();
 FILLCELL_X2 FILLER_130_1436 ();
 FILLCELL_X16 FILLER_130_1454 ();
 FILLCELL_X8 FILLER_130_1470 ();
 FILLCELL_X32 FILLER_130_1494 ();
 FILLCELL_X32 FILLER_130_1526 ();
 FILLCELL_X32 FILLER_130_1558 ();
 FILLCELL_X32 FILLER_130_1590 ();
 FILLCELL_X16 FILLER_130_1622 ();
 FILLCELL_X8 FILLER_130_1638 ();
 FILLCELL_X4 FILLER_130_1646 ();
 FILLCELL_X1 FILLER_130_1650 ();
 FILLCELL_X2 FILLER_131_1 ();
 FILLCELL_X1 FILLER_131_3 ();
 FILLCELL_X8 FILLER_131_51 ();
 FILLCELL_X2 FILLER_131_59 ();
 FILLCELL_X4 FILLER_131_81 ();
 FILLCELL_X1 FILLER_131_85 ();
 FILLCELL_X4 FILLER_131_126 ();
 FILLCELL_X4 FILLER_131_176 ();
 FILLCELL_X1 FILLER_131_180 ();
 FILLCELL_X4 FILLER_131_188 ();
 FILLCELL_X1 FILLER_131_192 ();
 FILLCELL_X4 FILLER_131_206 ();
 FILLCELL_X1 FILLER_131_210 ();
 FILLCELL_X8 FILLER_131_228 ();
 FILLCELL_X1 FILLER_131_236 ();
 FILLCELL_X4 FILLER_131_261 ();
 FILLCELL_X2 FILLER_131_265 ();
 FILLCELL_X1 FILLER_131_267 ();
 FILLCELL_X2 FILLER_131_277 ();
 FILLCELL_X2 FILLER_131_282 ();
 FILLCELL_X2 FILLER_131_304 ();
 FILLCELL_X1 FILLER_131_306 ();
 FILLCELL_X8 FILLER_131_351 ();
 FILLCELL_X4 FILLER_131_359 ();
 FILLCELL_X2 FILLER_131_387 ();
 FILLCELL_X1 FILLER_131_421 ();
 FILLCELL_X4 FILLER_131_449 ();
 FILLCELL_X2 FILLER_131_453 ();
 FILLCELL_X1 FILLER_131_472 ();
 FILLCELL_X8 FILLER_131_480 ();
 FILLCELL_X4 FILLER_131_488 ();
 FILLCELL_X4 FILLER_131_519 ();
 FILLCELL_X2 FILLER_131_523 ();
 FILLCELL_X1 FILLER_131_525 ();
 FILLCELL_X4 FILLER_131_530 ();
 FILLCELL_X1 FILLER_131_534 ();
 FILLCELL_X8 FILLER_131_562 ();
 FILLCELL_X2 FILLER_131_570 ();
 FILLCELL_X1 FILLER_131_572 ();
 FILLCELL_X1 FILLER_131_674 ();
 FILLCELL_X1 FILLER_131_682 ();
 FILLCELL_X16 FILLER_131_695 ();
 FILLCELL_X8 FILLER_131_711 ();
 FILLCELL_X4 FILLER_131_719 ();
 FILLCELL_X1 FILLER_131_723 ();
 FILLCELL_X32 FILLER_131_731 ();
 FILLCELL_X2 FILLER_131_763 ();
 FILLCELL_X1 FILLER_131_765 ();
 FILLCELL_X2 FILLER_131_773 ();
 FILLCELL_X1 FILLER_131_775 ();
 FILLCELL_X4 FILLER_131_802 ();
 FILLCELL_X8 FILLER_131_813 ();
 FILLCELL_X2 FILLER_131_821 ();
 FILLCELL_X1 FILLER_131_823 ();
 FILLCELL_X1 FILLER_131_831 ();
 FILLCELL_X1 FILLER_131_859 ();
 FILLCELL_X8 FILLER_131_865 ();
 FILLCELL_X2 FILLER_131_873 ();
 FILLCELL_X1 FILLER_131_875 ();
 FILLCELL_X2 FILLER_131_913 ();
 FILLCELL_X2 FILLER_131_932 ();
 FILLCELL_X4 FILLER_131_946 ();
 FILLCELL_X2 FILLER_131_950 ();
 FILLCELL_X4 FILLER_131_1006 ();
 FILLCELL_X2 FILLER_131_1010 ();
 FILLCELL_X8 FILLER_131_1059 ();
 FILLCELL_X4 FILLER_131_1067 ();
 FILLCELL_X2 FILLER_131_1071 ();
 FILLCELL_X1 FILLER_131_1073 ();
 FILLCELL_X2 FILLER_131_1084 ();
 FILLCELL_X1 FILLER_131_1086 ();
 FILLCELL_X2 FILLER_131_1093 ();
 FILLCELL_X1 FILLER_131_1101 ();
 FILLCELL_X4 FILLER_131_1108 ();
 FILLCELL_X4 FILLER_131_1122 ();
 FILLCELL_X4 FILLER_131_1132 ();
 FILLCELL_X2 FILLER_131_1148 ();
 FILLCELL_X2 FILLER_131_1170 ();
 FILLCELL_X1 FILLER_131_1172 ();
 FILLCELL_X4 FILLER_131_1199 ();
 FILLCELL_X2 FILLER_131_1221 ();
 FILLCELL_X1 FILLER_131_1223 ();
 FILLCELL_X2 FILLER_131_1234 ();
 FILLCELL_X2 FILLER_131_1242 ();
 FILLCELL_X2 FILLER_131_1250 ();
 FILLCELL_X1 FILLER_131_1252 ();
 FILLCELL_X4 FILLER_131_1259 ();
 FILLCELL_X1 FILLER_131_1264 ();
 FILLCELL_X2 FILLER_131_1275 ();
 FILLCELL_X4 FILLER_131_1293 ();
 FILLCELL_X4 FILLER_131_1319 ();
 FILLCELL_X1 FILLER_131_1323 ();
 FILLCELL_X1 FILLER_131_1338 ();
 FILLCELL_X2 FILLER_131_1343 ();
 FILLCELL_X32 FILLER_131_1350 ();
 FILLCELL_X16 FILLER_131_1382 ();
 FILLCELL_X8 FILLER_131_1398 ();
 FILLCELL_X2 FILLER_131_1406 ();
 FILLCELL_X4 FILLER_131_1415 ();
 FILLCELL_X2 FILLER_131_1419 ();
 FILLCELL_X1 FILLER_131_1421 ();
 FILLCELL_X4 FILLER_131_1429 ();
 FILLCELL_X1 FILLER_131_1433 ();
 FILLCELL_X1 FILLER_131_1464 ();
 FILLCELL_X1 FILLER_131_1474 ();
 FILLCELL_X1 FILLER_131_1484 ();
 FILLCELL_X32 FILLER_131_1494 ();
 FILLCELL_X32 FILLER_131_1526 ();
 FILLCELL_X32 FILLER_131_1558 ();
 FILLCELL_X32 FILLER_131_1590 ();
 FILLCELL_X16 FILLER_131_1622 ();
 FILLCELL_X8 FILLER_131_1638 ();
 FILLCELL_X4 FILLER_131_1646 ();
 FILLCELL_X1 FILLER_131_1650 ();
 FILLCELL_X4 FILLER_132_1 ();
 FILLCELL_X2 FILLER_132_5 ();
 FILLCELL_X1 FILLER_132_27 ();
 FILLCELL_X4 FILLER_132_37 ();
 FILLCELL_X1 FILLER_132_75 ();
 FILLCELL_X2 FILLER_132_85 ();
 FILLCELL_X4 FILLER_132_94 ();
 FILLCELL_X2 FILLER_132_98 ();
 FILLCELL_X1 FILLER_132_100 ();
 FILLCELL_X8 FILLER_132_108 ();
 FILLCELL_X2 FILLER_132_116 ();
 FILLCELL_X4 FILLER_132_123 ();
 FILLCELL_X2 FILLER_132_127 ();
 FILLCELL_X1 FILLER_132_129 ();
 FILLCELL_X4 FILLER_132_150 ();
 FILLCELL_X2 FILLER_132_154 ();
 FILLCELL_X4 FILLER_132_208 ();
 FILLCELL_X2 FILLER_132_212 ();
 FILLCELL_X1 FILLER_132_237 ();
 FILLCELL_X2 FILLER_132_242 ();
 FILLCELL_X2 FILLER_132_247 ();
 FILLCELL_X16 FILLER_132_261 ();
 FILLCELL_X8 FILLER_132_277 ();
 FILLCELL_X4 FILLER_132_292 ();
 FILLCELL_X2 FILLER_132_296 ();
 FILLCELL_X2 FILLER_132_327 ();
 FILLCELL_X1 FILLER_132_394 ();
 FILLCELL_X1 FILLER_132_407 ();
 FILLCELL_X1 FILLER_132_422 ();
 FILLCELL_X8 FILLER_132_427 ();
 FILLCELL_X2 FILLER_132_435 ();
 FILLCELL_X1 FILLER_132_437 ();
 FILLCELL_X16 FILLER_132_445 ();
 FILLCELL_X4 FILLER_132_490 ();
 FILLCELL_X4 FILLER_132_514 ();
 FILLCELL_X8 FILLER_132_538 ();
 FILLCELL_X2 FILLER_132_546 ();
 FILLCELL_X8 FILLER_132_557 ();
 FILLCELL_X2 FILLER_132_565 ();
 FILLCELL_X1 FILLER_132_567 ();
 FILLCELL_X2 FILLER_132_598 ();
 FILLCELL_X1 FILLER_132_604 ();
 FILLCELL_X2 FILLER_132_614 ();
 FILLCELL_X1 FILLER_132_616 ();
 FILLCELL_X8 FILLER_132_620 ();
 FILLCELL_X2 FILLER_132_628 ();
 FILLCELL_X1 FILLER_132_630 ();
 FILLCELL_X4 FILLER_132_663 ();
 FILLCELL_X2 FILLER_132_667 ();
 FILLCELL_X1 FILLER_132_669 ();
 FILLCELL_X4 FILLER_132_694 ();
 FILLCELL_X2 FILLER_132_698 ();
 FILLCELL_X1 FILLER_132_705 ();
 FILLCELL_X4 FILLER_132_710 ();
 FILLCELL_X1 FILLER_132_744 ();
 FILLCELL_X4 FILLER_132_752 ();
 FILLCELL_X16 FILLER_132_780 ();
 FILLCELL_X2 FILLER_132_796 ();
 FILLCELL_X1 FILLER_132_798 ();
 FILLCELL_X4 FILLER_132_813 ();
 FILLCELL_X1 FILLER_132_817 ();
 FILLCELL_X4 FILLER_132_830 ();
 FILLCELL_X2 FILLER_132_834 ();
 FILLCELL_X1 FILLER_132_836 ();
 FILLCELL_X2 FILLER_132_844 ();
 FILLCELL_X1 FILLER_132_846 ();
 FILLCELL_X4 FILLER_132_854 ();
 FILLCELL_X2 FILLER_132_885 ();
 FILLCELL_X1 FILLER_132_887 ();
 FILLCELL_X4 FILLER_132_908 ();
 FILLCELL_X1 FILLER_132_912 ();
 FILLCELL_X16 FILLER_132_956 ();
 FILLCELL_X4 FILLER_132_972 ();
 FILLCELL_X2 FILLER_132_976 ();
 FILLCELL_X4 FILLER_132_985 ();
 FILLCELL_X2 FILLER_132_989 ();
 FILLCELL_X4 FILLER_132_996 ();
 FILLCELL_X1 FILLER_132_1000 ();
 FILLCELL_X8 FILLER_132_1019 ();
 FILLCELL_X4 FILLER_132_1027 ();
 FILLCELL_X2 FILLER_132_1031 ();
 FILLCELL_X1 FILLER_132_1033 ();
 FILLCELL_X16 FILLER_132_1041 ();
 FILLCELL_X8 FILLER_132_1057 ();
 FILLCELL_X4 FILLER_132_1065 ();
 FILLCELL_X1 FILLER_132_1069 ();
 FILLCELL_X4 FILLER_132_1080 ();
 FILLCELL_X4 FILLER_132_1122 ();
 FILLCELL_X1 FILLER_132_1126 ();
 FILLCELL_X8 FILLER_132_1167 ();
 FILLCELL_X1 FILLER_132_1175 ();
 FILLCELL_X2 FILLER_132_1185 ();
 FILLCELL_X1 FILLER_132_1187 ();
 FILLCELL_X2 FILLER_132_1194 ();
 FILLCELL_X1 FILLER_132_1196 ();
 FILLCELL_X8 FILLER_132_1203 ();
 FILLCELL_X2 FILLER_132_1211 ();
 FILLCELL_X2 FILLER_132_1253 ();
 FILLCELL_X4 FILLER_132_1267 ();
 FILLCELL_X1 FILLER_132_1271 ();
 FILLCELL_X2 FILLER_132_1282 ();
 FILLCELL_X8 FILLER_132_1298 ();
 FILLCELL_X4 FILLER_132_1306 ();
 FILLCELL_X2 FILLER_132_1310 ();
 FILLCELL_X1 FILLER_132_1312 ();
 FILLCELL_X8 FILLER_132_1320 ();
 FILLCELL_X2 FILLER_132_1331 ();
 FILLCELL_X1 FILLER_132_1333 ();
 FILLCELL_X2 FILLER_132_1337 ();
 FILLCELL_X16 FILLER_132_1346 ();
 FILLCELL_X4 FILLER_132_1362 ();
 FILLCELL_X1 FILLER_132_1366 ();
 FILLCELL_X16 FILLER_132_1376 ();
 FILLCELL_X2 FILLER_132_1392 ();
 FILLCELL_X1 FILLER_132_1394 ();
 FILLCELL_X2 FILLER_132_1401 ();
 FILLCELL_X1 FILLER_132_1403 ();
 FILLCELL_X4 FILLER_132_1411 ();
 FILLCELL_X2 FILLER_132_1415 ();
 FILLCELL_X2 FILLER_132_1420 ();
 FILLCELL_X2 FILLER_132_1454 ();
 FILLCELL_X4 FILLER_132_1470 ();
 FILLCELL_X2 FILLER_132_1474 ();
 FILLCELL_X1 FILLER_132_1476 ();
 FILLCELL_X1 FILLER_132_1495 ();
 FILLCELL_X8 FILLER_132_1505 ();
 FILLCELL_X4 FILLER_132_1513 ();
 FILLCELL_X2 FILLER_132_1517 ();
 FILLCELL_X4 FILLER_132_1526 ();
 FILLCELL_X1 FILLER_132_1535 ();
 FILLCELL_X2 FILLER_132_1543 ();
 FILLCELL_X32 FILLER_132_1552 ();
 FILLCELL_X32 FILLER_132_1584 ();
 FILLCELL_X32 FILLER_132_1616 ();
 FILLCELL_X2 FILLER_132_1648 ();
 FILLCELL_X1 FILLER_132_1650 ();
 FILLCELL_X16 FILLER_133_1 ();
 FILLCELL_X2 FILLER_133_17 ();
 FILLCELL_X8 FILLER_133_33 ();
 FILLCELL_X2 FILLER_133_41 ();
 FILLCELL_X1 FILLER_133_43 ();
 FILLCELL_X16 FILLER_133_64 ();
 FILLCELL_X2 FILLER_133_100 ();
 FILLCELL_X16 FILLER_133_129 ();
 FILLCELL_X1 FILLER_133_145 ();
 FILLCELL_X32 FILLER_133_153 ();
 FILLCELL_X8 FILLER_133_185 ();
 FILLCELL_X2 FILLER_133_193 ();
 FILLCELL_X1 FILLER_133_195 ();
 FILLCELL_X2 FILLER_133_216 ();
 FILLCELL_X1 FILLER_133_218 ();
 FILLCELL_X8 FILLER_133_247 ();
 FILLCELL_X2 FILLER_133_255 ();
 FILLCELL_X2 FILLER_133_262 ();
 FILLCELL_X1 FILLER_133_264 ();
 FILLCELL_X1 FILLER_133_289 ();
 FILLCELL_X2 FILLER_133_293 ();
 FILLCELL_X1 FILLER_133_300 ();
 FILLCELL_X2 FILLER_133_308 ();
 FILLCELL_X1 FILLER_133_313 ();
 FILLCELL_X1 FILLER_133_331 ();
 FILLCELL_X4 FILLER_133_336 ();
 FILLCELL_X4 FILLER_133_351 ();
 FILLCELL_X2 FILLER_133_355 ();
 FILLCELL_X4 FILLER_133_384 ();
 FILLCELL_X1 FILLER_133_388 ();
 FILLCELL_X1 FILLER_133_413 ();
 FILLCELL_X1 FILLER_133_419 ();
 FILLCELL_X8 FILLER_133_447 ();
 FILLCELL_X2 FILLER_133_455 ();
 FILLCELL_X1 FILLER_133_466 ();
 FILLCELL_X1 FILLER_133_478 ();
 FILLCELL_X2 FILLER_133_484 ();
 FILLCELL_X1 FILLER_133_486 ();
 FILLCELL_X8 FILLER_133_508 ();
 FILLCELL_X2 FILLER_133_516 ();
 FILLCELL_X4 FILLER_133_525 ();
 FILLCELL_X1 FILLER_133_529 ();
 FILLCELL_X4 FILLER_133_564 ();
 FILLCELL_X2 FILLER_133_568 ();
 FILLCELL_X1 FILLER_133_578 ();
 FILLCELL_X1 FILLER_133_582 ();
 FILLCELL_X1 FILLER_133_588 ();
 FILLCELL_X32 FILLER_133_617 ();
 FILLCELL_X2 FILLER_133_673 ();
 FILLCELL_X2 FILLER_133_682 ();
 FILLCELL_X1 FILLER_133_704 ();
 FILLCELL_X1 FILLER_133_725 ();
 FILLCELL_X1 FILLER_133_747 ();
 FILLCELL_X2 FILLER_133_762 ();
 FILLCELL_X1 FILLER_133_792 ();
 FILLCELL_X1 FILLER_133_873 ();
 FILLCELL_X8 FILLER_133_881 ();
 FILLCELL_X4 FILLER_133_889 ();
 FILLCELL_X2 FILLER_133_952 ();
 FILLCELL_X8 FILLER_133_961 ();
 FILLCELL_X1 FILLER_133_969 ();
 FILLCELL_X4 FILLER_133_977 ();
 FILLCELL_X2 FILLER_133_981 ();
 FILLCELL_X1 FILLER_133_983 ();
 FILLCELL_X4 FILLER_133_988 ();
 FILLCELL_X8 FILLER_133_999 ();
 FILLCELL_X8 FILLER_133_1016 ();
 FILLCELL_X16 FILLER_133_1044 ();
 FILLCELL_X8 FILLER_133_1060 ();
 FILLCELL_X2 FILLER_133_1068 ();
 FILLCELL_X1 FILLER_133_1070 ();
 FILLCELL_X1 FILLER_133_1097 ();
 FILLCELL_X2 FILLER_133_1108 ();
 FILLCELL_X1 FILLER_133_1110 ();
 FILLCELL_X4 FILLER_133_1121 ();
 FILLCELL_X1 FILLER_133_1141 ();
 FILLCELL_X2 FILLER_133_1152 ();
 FILLCELL_X2 FILLER_133_1157 ();
 FILLCELL_X2 FILLER_133_1181 ();
 FILLCELL_X8 FILLER_133_1213 ();
 FILLCELL_X1 FILLER_133_1221 ();
 FILLCELL_X4 FILLER_133_1232 ();
 FILLCELL_X4 FILLER_133_1258 ();
 FILLCELL_X1 FILLER_133_1262 ();
 FILLCELL_X4 FILLER_133_1286 ();
 FILLCELL_X2 FILLER_133_1290 ();
 FILLCELL_X1 FILLER_133_1292 ();
 FILLCELL_X1 FILLER_133_1328 ();
 FILLCELL_X4 FILLER_133_1336 ();
 FILLCELL_X2 FILLER_133_1340 ();
 FILLCELL_X1 FILLER_133_1359 ();
 FILLCELL_X1 FILLER_133_1369 ();
 FILLCELL_X2 FILLER_133_1386 ();
 FILLCELL_X4 FILLER_133_1406 ();
 FILLCELL_X1 FILLER_133_1410 ();
 FILLCELL_X2 FILLER_133_1415 ();
 FILLCELL_X4 FILLER_133_1426 ();
 FILLCELL_X2 FILLER_133_1430 ();
 FILLCELL_X8 FILLER_133_1439 ();
 FILLCELL_X2 FILLER_133_1447 ();
 FILLCELL_X2 FILLER_133_1453 ();
 FILLCELL_X8 FILLER_133_1483 ();
 FILLCELL_X1 FILLER_133_1503 ();
 FILLCELL_X1 FILLER_133_1533 ();
 FILLCELL_X32 FILLER_133_1543 ();
 FILLCELL_X32 FILLER_133_1575 ();
 FILLCELL_X32 FILLER_133_1607 ();
 FILLCELL_X8 FILLER_133_1639 ();
 FILLCELL_X4 FILLER_133_1647 ();
 FILLCELL_X16 FILLER_134_1 ();
 FILLCELL_X2 FILLER_134_17 ();
 FILLCELL_X1 FILLER_134_19 ();
 FILLCELL_X8 FILLER_134_27 ();
 FILLCELL_X4 FILLER_134_35 ();
 FILLCELL_X4 FILLER_134_47 ();
 FILLCELL_X8 FILLER_134_78 ();
 FILLCELL_X2 FILLER_134_86 ();
 FILLCELL_X8 FILLER_134_99 ();
 FILLCELL_X1 FILLER_134_107 ();
 FILLCELL_X2 FILLER_134_113 ();
 FILLCELL_X1 FILLER_134_115 ();
 FILLCELL_X4 FILLER_134_156 ();
 FILLCELL_X1 FILLER_134_187 ();
 FILLCELL_X1 FILLER_134_202 ();
 FILLCELL_X1 FILLER_134_207 ();
 FILLCELL_X1 FILLER_134_215 ();
 FILLCELL_X2 FILLER_134_224 ();
 FILLCELL_X2 FILLER_134_230 ();
 FILLCELL_X1 FILLER_134_255 ();
 FILLCELL_X1 FILLER_134_281 ();
 FILLCELL_X2 FILLER_134_306 ();
 FILLCELL_X4 FILLER_134_316 ();
 FILLCELL_X2 FILLER_134_320 ();
 FILLCELL_X1 FILLER_134_322 ();
 FILLCELL_X1 FILLER_134_326 ();
 FILLCELL_X16 FILLER_134_339 ();
 FILLCELL_X4 FILLER_134_355 ();
 FILLCELL_X2 FILLER_134_363 ();
 FILLCELL_X8 FILLER_134_368 ();
 FILLCELL_X1 FILLER_134_376 ();
 FILLCELL_X1 FILLER_134_442 ();
 FILLCELL_X1 FILLER_134_480 ();
 FILLCELL_X2 FILLER_134_491 ();
 FILLCELL_X1 FILLER_134_493 ();
 FILLCELL_X2 FILLER_134_508 ();
 FILLCELL_X1 FILLER_134_510 ();
 FILLCELL_X4 FILLER_134_524 ();
 FILLCELL_X2 FILLER_134_528 ();
 FILLCELL_X1 FILLER_134_530 ();
 FILLCELL_X2 FILLER_134_569 ();
 FILLCELL_X1 FILLER_134_571 ();
 FILLCELL_X8 FILLER_134_579 ();
 FILLCELL_X4 FILLER_134_587 ();
 FILLCELL_X2 FILLER_134_632 ();
 FILLCELL_X1 FILLER_134_634 ();
 FILLCELL_X4 FILLER_134_638 ();
 FILLCELL_X16 FILLER_134_673 ();
 FILLCELL_X2 FILLER_134_689 ();
 FILLCELL_X4 FILLER_134_695 ();
 FILLCELL_X8 FILLER_134_702 ();
 FILLCELL_X1 FILLER_134_710 ();
 FILLCELL_X4 FILLER_134_744 ();
 FILLCELL_X2 FILLER_134_748 ();
 FILLCELL_X1 FILLER_134_750 ();
 FILLCELL_X1 FILLER_134_758 ();
 FILLCELL_X8 FILLER_134_786 ();
 FILLCELL_X4 FILLER_134_794 ();
 FILLCELL_X4 FILLER_134_821 ();
 FILLCELL_X2 FILLER_134_825 ();
 FILLCELL_X1 FILLER_134_832 ();
 FILLCELL_X4 FILLER_134_838 ();
 FILLCELL_X8 FILLER_134_847 ();
 FILLCELL_X4 FILLER_134_855 ();
 FILLCELL_X16 FILLER_134_886 ();
 FILLCELL_X32 FILLER_134_909 ();
 FILLCELL_X8 FILLER_134_941 ();
 FILLCELL_X1 FILLER_134_949 ();
 FILLCELL_X4 FILLER_134_1010 ();
 FILLCELL_X2 FILLER_134_1014 ();
 FILLCELL_X2 FILLER_134_1036 ();
 FILLCELL_X8 FILLER_134_1058 ();
 FILLCELL_X4 FILLER_134_1066 ();
 FILLCELL_X1 FILLER_134_1080 ();
 FILLCELL_X1 FILLER_134_1087 ();
 FILLCELL_X1 FILLER_134_1094 ();
 FILLCELL_X1 FILLER_134_1123 ();
 FILLCELL_X1 FILLER_134_1130 ();
 FILLCELL_X2 FILLER_134_1141 ();
 FILLCELL_X4 FILLER_134_1163 ();
 FILLCELL_X8 FILLER_134_1174 ();
 FILLCELL_X1 FILLER_134_1182 ();
 FILLCELL_X1 FILLER_134_1201 ();
 FILLCELL_X2 FILLER_134_1208 ();
 FILLCELL_X1 FILLER_134_1267 ();
 FILLCELL_X2 FILLER_134_1278 ();
 FILLCELL_X16 FILLER_134_1300 ();
 FILLCELL_X2 FILLER_134_1316 ();
 FILLCELL_X8 FILLER_134_1325 ();
 FILLCELL_X8 FILLER_134_1336 ();
 FILLCELL_X2 FILLER_134_1344 ();
 FILLCELL_X1 FILLER_134_1359 ();
 FILLCELL_X1 FILLER_134_1367 ();
 FILLCELL_X8 FILLER_134_1381 ();
 FILLCELL_X4 FILLER_134_1389 ();
 FILLCELL_X2 FILLER_134_1393 ();
 FILLCELL_X16 FILLER_134_1413 ();
 FILLCELL_X4 FILLER_134_1450 ();
 FILLCELL_X2 FILLER_134_1454 ();
 FILLCELL_X1 FILLER_134_1456 ();
 FILLCELL_X2 FILLER_134_1471 ();
 FILLCELL_X1 FILLER_134_1493 ();
 FILLCELL_X2 FILLER_134_1513 ();
 FILLCELL_X1 FILLER_134_1536 ();
 FILLCELL_X32 FILLER_134_1546 ();
 FILLCELL_X32 FILLER_134_1578 ();
 FILLCELL_X32 FILLER_134_1610 ();
 FILLCELL_X8 FILLER_134_1642 ();
 FILLCELL_X1 FILLER_134_1650 ();
 FILLCELL_X8 FILLER_135_1 ();
 FILLCELL_X1 FILLER_135_9 ();
 FILLCELL_X1 FILLER_135_30 ();
 FILLCELL_X8 FILLER_135_58 ();
 FILLCELL_X2 FILLER_135_66 ();
 FILLCELL_X1 FILLER_135_68 ();
 FILLCELL_X8 FILLER_135_76 ();
 FILLCELL_X2 FILLER_135_84 ();
 FILLCELL_X1 FILLER_135_86 ();
 FILLCELL_X2 FILLER_135_114 ();
 FILLCELL_X1 FILLER_135_116 ();
 FILLCELL_X16 FILLER_135_135 ();
 FILLCELL_X1 FILLER_135_151 ();
 FILLCELL_X2 FILLER_135_156 ();
 FILLCELL_X4 FILLER_135_198 ();
 FILLCELL_X1 FILLER_135_202 ();
 FILLCELL_X16 FILLER_135_223 ();
 FILLCELL_X1 FILLER_135_267 ();
 FILLCELL_X2 FILLER_135_272 ();
 FILLCELL_X1 FILLER_135_274 ();
 FILLCELL_X4 FILLER_135_278 ();
 FILLCELL_X2 FILLER_135_282 ();
 FILLCELL_X1 FILLER_135_284 ();
 FILLCELL_X4 FILLER_135_289 ();
 FILLCELL_X2 FILLER_135_296 ();
 FILLCELL_X2 FILLER_135_301 ();
 FILLCELL_X2 FILLER_135_346 ();
 FILLCELL_X1 FILLER_135_348 ();
 FILLCELL_X16 FILLER_135_356 ();
 FILLCELL_X4 FILLER_135_372 ();
 FILLCELL_X2 FILLER_135_376 ();
 FILLCELL_X2 FILLER_135_385 ();
 FILLCELL_X4 FILLER_135_394 ();
 FILLCELL_X1 FILLER_135_398 ();
 FILLCELL_X1 FILLER_135_424 ();
 FILLCELL_X2 FILLER_135_429 ();
 FILLCELL_X8 FILLER_135_439 ();
 FILLCELL_X4 FILLER_135_447 ();
 FILLCELL_X2 FILLER_135_458 ();
 FILLCELL_X1 FILLER_135_460 ();
 FILLCELL_X2 FILLER_135_466 ();
 FILLCELL_X1 FILLER_135_468 ();
 FILLCELL_X16 FILLER_135_478 ();
 FILLCELL_X8 FILLER_135_494 ();
 FILLCELL_X1 FILLER_135_502 ();
 FILLCELL_X2 FILLER_135_510 ();
 FILLCELL_X1 FILLER_135_512 ();
 FILLCELL_X1 FILLER_135_516 ();
 FILLCELL_X16 FILLER_135_520 ();
 FILLCELL_X4 FILLER_135_536 ();
 FILLCELL_X1 FILLER_135_540 ();
 FILLCELL_X2 FILLER_135_548 ();
 FILLCELL_X1 FILLER_135_550 ();
 FILLCELL_X8 FILLER_135_588 ();
 FILLCELL_X2 FILLER_135_596 ();
 FILLCELL_X8 FILLER_135_601 ();
 FILLCELL_X2 FILLER_135_609 ();
 FILLCELL_X1 FILLER_135_611 ();
 FILLCELL_X4 FILLER_135_644 ();
 FILLCELL_X1 FILLER_135_648 ();
 FILLCELL_X2 FILLER_135_653 ();
 FILLCELL_X1 FILLER_135_655 ();
 FILLCELL_X1 FILLER_135_664 ();
 FILLCELL_X2 FILLER_135_707 ();
 FILLCELL_X16 FILLER_135_712 ();
 FILLCELL_X2 FILLER_135_728 ();
 FILLCELL_X2 FILLER_135_737 ();
 FILLCELL_X8 FILLER_135_759 ();
 FILLCELL_X4 FILLER_135_767 ();
 FILLCELL_X1 FILLER_135_771 ();
 FILLCELL_X2 FILLER_135_776 ();
 FILLCELL_X2 FILLER_135_780 ();
 FILLCELL_X8 FILLER_135_814 ();
 FILLCELL_X4 FILLER_135_822 ();
 FILLCELL_X1 FILLER_135_833 ();
 FILLCELL_X1 FILLER_135_861 ();
 FILLCELL_X16 FILLER_135_900 ();
 FILLCELL_X2 FILLER_135_916 ();
 FILLCELL_X1 FILLER_135_918 ();
 FILLCELL_X16 FILLER_135_939 ();
 FILLCELL_X4 FILLER_135_955 ();
 FILLCELL_X8 FILLER_135_964 ();
 FILLCELL_X1 FILLER_135_977 ();
 FILLCELL_X1 FILLER_135_983 ();
 FILLCELL_X2 FILLER_135_1022 ();
 FILLCELL_X2 FILLER_135_1031 ();
 FILLCELL_X2 FILLER_135_1040 ();
 FILLCELL_X1 FILLER_135_1042 ();
 FILLCELL_X2 FILLER_135_1050 ();
 FILLCELL_X1 FILLER_135_1052 ();
 FILLCELL_X2 FILLER_135_1073 ();
 FILLCELL_X1 FILLER_135_1081 ();
 FILLCELL_X4 FILLER_135_1101 ();
 FILLCELL_X4 FILLER_135_1115 ();
 FILLCELL_X1 FILLER_135_1119 ();
 FILLCELL_X8 FILLER_135_1130 ();
 FILLCELL_X4 FILLER_135_1138 ();
 FILLCELL_X1 FILLER_135_1142 ();
 FILLCELL_X4 FILLER_135_1158 ();
 FILLCELL_X1 FILLER_135_1162 ();
 FILLCELL_X4 FILLER_135_1169 ();
 FILLCELL_X2 FILLER_135_1173 ();
 FILLCELL_X4 FILLER_135_1179 ();
 FILLCELL_X2 FILLER_135_1190 ();
 FILLCELL_X1 FILLER_135_1192 ();
 FILLCELL_X8 FILLER_135_1199 ();
 FILLCELL_X2 FILLER_135_1207 ();
 FILLCELL_X1 FILLER_135_1215 ();
 FILLCELL_X4 FILLER_135_1226 ();
 FILLCELL_X4 FILLER_135_1246 ();
 FILLCELL_X1 FILLER_135_1256 ();
 FILLCELL_X4 FILLER_135_1292 ();
 FILLCELL_X1 FILLER_135_1296 ();
 FILLCELL_X2 FILLER_135_1300 ();
 FILLCELL_X1 FILLER_135_1306 ();
 FILLCELL_X2 FILLER_135_1327 ();
 FILLCELL_X16 FILLER_135_1333 ();
 FILLCELL_X1 FILLER_135_1349 ();
 FILLCELL_X2 FILLER_135_1354 ();
 FILLCELL_X4 FILLER_135_1363 ();
 FILLCELL_X2 FILLER_135_1367 ();
 FILLCELL_X1 FILLER_135_1369 ();
 FILLCELL_X8 FILLER_135_1379 ();
 FILLCELL_X4 FILLER_135_1387 ();
 FILLCELL_X1 FILLER_135_1391 ();
 FILLCELL_X4 FILLER_135_1406 ();
 FILLCELL_X2 FILLER_135_1410 ();
 FILLCELL_X4 FILLER_135_1426 ();
 FILLCELL_X2 FILLER_135_1433 ();
 FILLCELL_X1 FILLER_135_1435 ();
 FILLCELL_X4 FILLER_135_1439 ();
 FILLCELL_X1 FILLER_135_1443 ();
 FILLCELL_X2 FILLER_135_1449 ();
 FILLCELL_X1 FILLER_135_1451 ();
 FILLCELL_X4 FILLER_135_1478 ();
 FILLCELL_X1 FILLER_135_1491 ();
 FILLCELL_X1 FILLER_135_1503 ();
 FILLCELL_X4 FILLER_135_1508 ();
 FILLCELL_X1 FILLER_135_1512 ();
 FILLCELL_X4 FILLER_135_1522 ();
 FILLCELL_X2 FILLER_135_1526 ();
 FILLCELL_X1 FILLER_135_1528 ();
 FILLCELL_X4 FILLER_135_1536 ();
 FILLCELL_X2 FILLER_135_1540 ();
 FILLCELL_X1 FILLER_135_1542 ();
 FILLCELL_X32 FILLER_135_1546 ();
 FILLCELL_X32 FILLER_135_1578 ();
 FILLCELL_X32 FILLER_135_1610 ();
 FILLCELL_X8 FILLER_135_1642 ();
 FILLCELL_X1 FILLER_135_1650 ();
 FILLCELL_X4 FILLER_136_21 ();
 FILLCELL_X1 FILLER_136_25 ();
 FILLCELL_X4 FILLER_136_35 ();
 FILLCELL_X1 FILLER_136_39 ();
 FILLCELL_X2 FILLER_136_61 ();
 FILLCELL_X1 FILLER_136_63 ();
 FILLCELL_X2 FILLER_136_91 ();
 FILLCELL_X1 FILLER_136_93 ();
 FILLCELL_X2 FILLER_136_114 ();
 FILLCELL_X2 FILLER_136_134 ();
 FILLCELL_X1 FILLER_136_156 ();
 FILLCELL_X2 FILLER_136_178 ();
 FILLCELL_X1 FILLER_136_180 ();
 FILLCELL_X1 FILLER_136_188 ();
 FILLCELL_X2 FILLER_136_200 ();
 FILLCELL_X1 FILLER_136_202 ();
 FILLCELL_X16 FILLER_136_230 ();
 FILLCELL_X4 FILLER_136_246 ();
 FILLCELL_X2 FILLER_136_250 ();
 FILLCELL_X1 FILLER_136_256 ();
 FILLCELL_X2 FILLER_136_262 ();
 FILLCELL_X4 FILLER_136_267 ();
 FILLCELL_X2 FILLER_136_271 ();
 FILLCELL_X4 FILLER_136_293 ();
 FILLCELL_X2 FILLER_136_306 ();
 FILLCELL_X8 FILLER_136_316 ();
 FILLCELL_X4 FILLER_136_326 ();
 FILLCELL_X4 FILLER_136_335 ();
 FILLCELL_X1 FILLER_136_339 ();
 FILLCELL_X2 FILLER_136_371 ();
 FILLCELL_X8 FILLER_136_393 ();
 FILLCELL_X4 FILLER_136_401 ();
 FILLCELL_X2 FILLER_136_405 ();
 FILLCELL_X1 FILLER_136_407 ();
 FILLCELL_X4 FILLER_136_412 ();
 FILLCELL_X4 FILLER_136_419 ();
 FILLCELL_X2 FILLER_136_423 ();
 FILLCELL_X8 FILLER_136_432 ();
 FILLCELL_X4 FILLER_136_440 ();
 FILLCELL_X1 FILLER_136_444 ();
 FILLCELL_X4 FILLER_136_452 ();
 FILLCELL_X1 FILLER_136_456 ();
 FILLCELL_X1 FILLER_136_508 ();
 FILLCELL_X4 FILLER_136_533 ();
 FILLCELL_X2 FILLER_136_537 ();
 FILLCELL_X4 FILLER_136_544 ();
 FILLCELL_X2 FILLER_136_548 ();
 FILLCELL_X1 FILLER_136_550 ();
 FILLCELL_X1 FILLER_136_556 ();
 FILLCELL_X2 FILLER_136_568 ();
 FILLCELL_X4 FILLER_136_575 ();
 FILLCELL_X2 FILLER_136_579 ();
 FILLCELL_X4 FILLER_136_588 ();
 FILLCELL_X1 FILLER_136_592 ();
 FILLCELL_X4 FILLER_136_600 ();
 FILLCELL_X2 FILLER_136_604 ();
 FILLCELL_X1 FILLER_136_606 ();
 FILLCELL_X8 FILLER_136_611 ();
 FILLCELL_X2 FILLER_136_619 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X2 FILLER_136_632 ();
 FILLCELL_X1 FILLER_136_634 ();
 FILLCELL_X1 FILLER_136_662 ();
 FILLCELL_X4 FILLER_136_667 ();
 FILLCELL_X2 FILLER_136_671 ();
 FILLCELL_X1 FILLER_136_737 ();
 FILLCELL_X1 FILLER_136_763 ();
 FILLCELL_X2 FILLER_136_788 ();
 FILLCELL_X1 FILLER_136_790 ();
 FILLCELL_X4 FILLER_136_798 ();
 FILLCELL_X1 FILLER_136_802 ();
 FILLCELL_X2 FILLER_136_810 ();
 FILLCELL_X4 FILLER_136_857 ();
 FILLCELL_X4 FILLER_136_872 ();
 FILLCELL_X1 FILLER_136_876 ();
 FILLCELL_X1 FILLER_136_897 ();
 FILLCELL_X8 FILLER_136_905 ();
 FILLCELL_X4 FILLER_136_913 ();
 FILLCELL_X2 FILLER_136_917 ();
 FILLCELL_X1 FILLER_136_919 ();
 FILLCELL_X4 FILLER_136_933 ();
 FILLCELL_X1 FILLER_136_937 ();
 FILLCELL_X1 FILLER_136_978 ();
 FILLCELL_X2 FILLER_136_986 ();
 FILLCELL_X1 FILLER_136_988 ();
 FILLCELL_X1 FILLER_136_994 ();
 FILLCELL_X16 FILLER_136_1022 ();
 FILLCELL_X2 FILLER_136_1038 ();
 FILLCELL_X1 FILLER_136_1040 ();
 FILLCELL_X8 FILLER_136_1062 ();
 FILLCELL_X4 FILLER_136_1070 ();
 FILLCELL_X2 FILLER_136_1074 ();
 FILLCELL_X1 FILLER_136_1082 ();
 FILLCELL_X1 FILLER_136_1089 ();
 FILLCELL_X2 FILLER_136_1096 ();
 FILLCELL_X4 FILLER_136_1134 ();
 FILLCELL_X2 FILLER_136_1138 ();
 FILLCELL_X8 FILLER_136_1168 ();
 FILLCELL_X2 FILLER_136_1176 ();
 FILLCELL_X2 FILLER_136_1209 ();
 FILLCELL_X1 FILLER_136_1211 ();
 FILLCELL_X1 FILLER_136_1234 ();
 FILLCELL_X8 FILLER_136_1261 ();
 FILLCELL_X1 FILLER_136_1269 ();
 FILLCELL_X2 FILLER_136_1297 ();
 FILLCELL_X4 FILLER_136_1305 ();
 FILLCELL_X2 FILLER_136_1309 ();
 FILLCELL_X1 FILLER_136_1311 ();
 FILLCELL_X16 FILLER_136_1339 ();
 FILLCELL_X4 FILLER_136_1355 ();
 FILLCELL_X1 FILLER_136_1359 ();
 FILLCELL_X2 FILLER_136_1381 ();
 FILLCELL_X1 FILLER_136_1383 ();
 FILLCELL_X4 FILLER_136_1406 ();
 FILLCELL_X1 FILLER_136_1449 ();
 FILLCELL_X4 FILLER_136_1457 ();
 FILLCELL_X2 FILLER_136_1461 ();
 FILLCELL_X2 FILLER_136_1466 ();
 FILLCELL_X1 FILLER_136_1468 ();
 FILLCELL_X8 FILLER_136_1473 ();
 FILLCELL_X4 FILLER_136_1481 ();
 FILLCELL_X2 FILLER_136_1485 ();
 FILLCELL_X1 FILLER_136_1487 ();
 FILLCELL_X2 FILLER_136_1495 ();
 FILLCELL_X4 FILLER_136_1507 ();
 FILLCELL_X1 FILLER_136_1511 ();
 FILLCELL_X4 FILLER_136_1529 ();
 FILLCELL_X2 FILLER_136_1533 ();
 FILLCELL_X2 FILLER_136_1546 ();
 FILLCELL_X1 FILLER_136_1548 ();
 FILLCELL_X4 FILLER_136_1563 ();
 FILLCELL_X2 FILLER_136_1567 ();
 FILLCELL_X1 FILLER_136_1569 ();
 FILLCELL_X4 FILLER_136_1574 ();
 FILLCELL_X32 FILLER_136_1585 ();
 FILLCELL_X32 FILLER_136_1617 ();
 FILLCELL_X2 FILLER_136_1649 ();
 FILLCELL_X8 FILLER_137_1 ();
 FILLCELL_X2 FILLER_137_9 ();
 FILLCELL_X1 FILLER_137_11 ();
 FILLCELL_X1 FILLER_137_39 ();
 FILLCELL_X16 FILLER_137_67 ();
 FILLCELL_X4 FILLER_137_103 ();
 FILLCELL_X2 FILLER_137_107 ();
 FILLCELL_X2 FILLER_137_135 ();
 FILLCELL_X1 FILLER_137_137 ();
 FILLCELL_X4 FILLER_137_145 ();
 FILLCELL_X1 FILLER_137_154 ();
 FILLCELL_X4 FILLER_137_190 ();
 FILLCELL_X2 FILLER_137_194 ();
 FILLCELL_X8 FILLER_137_216 ();
 FILLCELL_X4 FILLER_137_224 ();
 FILLCELL_X1 FILLER_137_255 ();
 FILLCELL_X4 FILLER_137_269 ();
 FILLCELL_X2 FILLER_137_273 ();
 FILLCELL_X1 FILLER_137_275 ();
 FILLCELL_X2 FILLER_137_391 ();
 FILLCELL_X4 FILLER_137_397 ();
 FILLCELL_X1 FILLER_137_401 ();
 FILLCELL_X1 FILLER_137_442 ();
 FILLCELL_X1 FILLER_137_450 ();
 FILLCELL_X4 FILLER_137_460 ();
 FILLCELL_X1 FILLER_137_471 ();
 FILLCELL_X2 FILLER_137_509 ();
 FILLCELL_X2 FILLER_137_520 ();
 FILLCELL_X2 FILLER_137_527 ();
 FILLCELL_X4 FILLER_137_572 ();
 FILLCELL_X1 FILLER_137_576 ();
 FILLCELL_X4 FILLER_137_597 ();
 FILLCELL_X8 FILLER_137_635 ();
 FILLCELL_X2 FILLER_137_643 ();
 FILLCELL_X1 FILLER_137_652 ();
 FILLCELL_X1 FILLER_137_657 ();
 FILLCELL_X1 FILLER_137_661 ();
 FILLCELL_X1 FILLER_137_667 ();
 FILLCELL_X4 FILLER_137_696 ();
 FILLCELL_X4 FILLER_137_707 ();
 FILLCELL_X1 FILLER_137_711 ();
 FILLCELL_X8 FILLER_137_756 ();
 FILLCELL_X2 FILLER_137_764 ();
 FILLCELL_X1 FILLER_137_766 ();
 FILLCELL_X1 FILLER_137_778 ();
 FILLCELL_X2 FILLER_137_792 ();
 FILLCELL_X1 FILLER_137_794 ();
 FILLCELL_X8 FILLER_137_829 ();
 FILLCELL_X2 FILLER_137_837 ();
 FILLCELL_X2 FILLER_137_846 ();
 FILLCELL_X4 FILLER_137_868 ();
 FILLCELL_X2 FILLER_137_872 ();
 FILLCELL_X1 FILLER_137_874 ();
 FILLCELL_X16 FILLER_137_889 ();
 FILLCELL_X4 FILLER_137_959 ();
 FILLCELL_X1 FILLER_137_963 ();
 FILLCELL_X8 FILLER_137_968 ();
 FILLCELL_X2 FILLER_137_976 ();
 FILLCELL_X1 FILLER_137_978 ();
 FILLCELL_X1 FILLER_137_990 ();
 FILLCELL_X4 FILLER_137_1017 ();
 FILLCELL_X2 FILLER_137_1021 ();
 FILLCELL_X1 FILLER_137_1023 ();
 FILLCELL_X8 FILLER_137_1069 ();
 FILLCELL_X4 FILLER_137_1077 ();
 FILLCELL_X1 FILLER_137_1081 ();
 FILLCELL_X2 FILLER_137_1098 ();
 FILLCELL_X16 FILLER_137_1110 ();
 FILLCELL_X2 FILLER_137_1138 ();
 FILLCELL_X8 FILLER_137_1166 ();
 FILLCELL_X1 FILLER_137_1186 ();
 FILLCELL_X1 FILLER_137_1193 ();
 FILLCELL_X8 FILLER_137_1210 ();
 FILLCELL_X8 FILLER_137_1234 ();
 FILLCELL_X2 FILLER_137_1260 ();
 FILLCELL_X1 FILLER_137_1262 ();
 FILLCELL_X2 FILLER_137_1264 ();
 FILLCELL_X1 FILLER_137_1276 ();
 FILLCELL_X2 FILLER_137_1283 ();
 FILLCELL_X32 FILLER_137_1295 ();
 FILLCELL_X32 FILLER_137_1327 ();
 FILLCELL_X4 FILLER_137_1359 ();
 FILLCELL_X1 FILLER_137_1363 ();
 FILLCELL_X4 FILLER_137_1382 ();
 FILLCELL_X1 FILLER_137_1401 ();
 FILLCELL_X1 FILLER_137_1414 ();
 FILLCELL_X2 FILLER_137_1428 ();
 FILLCELL_X1 FILLER_137_1430 ();
 FILLCELL_X16 FILLER_137_1440 ();
 FILLCELL_X4 FILLER_137_1456 ();
 FILLCELL_X2 FILLER_137_1460 ();
 FILLCELL_X2 FILLER_137_1476 ();
 FILLCELL_X1 FILLER_137_1478 ();
 FILLCELL_X1 FILLER_137_1502 ();
 FILLCELL_X1 FILLER_137_1528 ();
 FILLCELL_X1 FILLER_137_1540 ();
 FILLCELL_X2 FILLER_137_1548 ();
 FILLCELL_X32 FILLER_137_1557 ();
 FILLCELL_X32 FILLER_137_1589 ();
 FILLCELL_X16 FILLER_137_1621 ();
 FILLCELL_X8 FILLER_137_1637 ();
 FILLCELL_X4 FILLER_137_1645 ();
 FILLCELL_X2 FILLER_137_1649 ();
 FILLCELL_X2 FILLER_138_21 ();
 FILLCELL_X2 FILLER_138_43 ();
 FILLCELL_X1 FILLER_138_45 ();
 FILLCELL_X16 FILLER_138_55 ();
 FILLCELL_X4 FILLER_138_71 ();
 FILLCELL_X16 FILLER_138_80 ();
 FILLCELL_X2 FILLER_138_96 ();
 FILLCELL_X1 FILLER_138_98 ();
 FILLCELL_X1 FILLER_138_138 ();
 FILLCELL_X2 FILLER_138_159 ();
 FILLCELL_X1 FILLER_138_161 ();
 FILLCELL_X4 FILLER_138_174 ();
 FILLCELL_X2 FILLER_138_178 ();
 FILLCELL_X1 FILLER_138_180 ();
 FILLCELL_X16 FILLER_138_188 ();
 FILLCELL_X2 FILLER_138_221 ();
 FILLCELL_X1 FILLER_138_223 ();
 FILLCELL_X2 FILLER_138_238 ();
 FILLCELL_X1 FILLER_138_240 ();
 FILLCELL_X4 FILLER_138_268 ();
 FILLCELL_X1 FILLER_138_272 ();
 FILLCELL_X1 FILLER_138_301 ();
 FILLCELL_X4 FILLER_138_308 ();
 FILLCELL_X1 FILLER_138_312 ();
 FILLCELL_X1 FILLER_138_369 ();
 FILLCELL_X4 FILLER_138_402 ();
 FILLCELL_X2 FILLER_138_406 ();
 FILLCELL_X4 FILLER_138_442 ();
 FILLCELL_X16 FILLER_138_468 ();
 FILLCELL_X8 FILLER_138_484 ();
 FILLCELL_X2 FILLER_138_492 ();
 FILLCELL_X1 FILLER_138_535 ();
 FILLCELL_X2 FILLER_138_556 ();
 FILLCELL_X1 FILLER_138_558 ();
 FILLCELL_X1 FILLER_138_632 ();
 FILLCELL_X8 FILLER_138_636 ();
 FILLCELL_X1 FILLER_138_644 ();
 FILLCELL_X16 FILLER_138_694 ();
 FILLCELL_X8 FILLER_138_710 ();
 FILLCELL_X4 FILLER_138_718 ();
 FILLCELL_X1 FILLER_138_768 ();
 FILLCELL_X2 FILLER_138_809 ();
 FILLCELL_X16 FILLER_138_816 ();
 FILLCELL_X4 FILLER_138_832 ();
 FILLCELL_X8 FILLER_138_840 ();
 FILLCELL_X4 FILLER_138_848 ();
 FILLCELL_X4 FILLER_138_859 ();
 FILLCELL_X2 FILLER_138_863 ();
 FILLCELL_X1 FILLER_138_865 ();
 FILLCELL_X8 FILLER_138_871 ();
 FILLCELL_X1 FILLER_138_879 ();
 FILLCELL_X4 FILLER_138_961 ();
 FILLCELL_X2 FILLER_138_965 ();
 FILLCELL_X1 FILLER_138_975 ();
 FILLCELL_X2 FILLER_138_996 ();
 FILLCELL_X1 FILLER_138_1005 ();
 FILLCELL_X2 FILLER_138_1018 ();
 FILLCELL_X1 FILLER_138_1020 ();
 FILLCELL_X8 FILLER_138_1028 ();
 FILLCELL_X2 FILLER_138_1036 ();
 FILLCELL_X1 FILLER_138_1038 ();
 FILLCELL_X4 FILLER_138_1042 ();
 FILLCELL_X16 FILLER_138_1073 ();
 FILLCELL_X4 FILLER_138_1089 ();
 FILLCELL_X1 FILLER_138_1093 ();
 FILLCELL_X1 FILLER_138_1110 ();
 FILLCELL_X4 FILLER_138_1117 ();
 FILLCELL_X1 FILLER_138_1121 ();
 FILLCELL_X16 FILLER_138_1131 ();
 FILLCELL_X8 FILLER_138_1147 ();
 FILLCELL_X8 FILLER_138_1171 ();
 FILLCELL_X1 FILLER_138_1203 ();
 FILLCELL_X4 FILLER_138_1210 ();
 FILLCELL_X1 FILLER_138_1214 ();
 FILLCELL_X2 FILLER_138_1231 ();
 FILLCELL_X1 FILLER_138_1239 ();
 FILLCELL_X1 FILLER_138_1246 ();
 FILLCELL_X2 FILLER_138_1263 ();
 FILLCELL_X1 FILLER_138_1265 ();
 FILLCELL_X2 FILLER_138_1286 ();
 FILLCELL_X32 FILLER_138_1306 ();
 FILLCELL_X32 FILLER_138_1338 ();
 FILLCELL_X2 FILLER_138_1370 ();
 FILLCELL_X1 FILLER_138_1372 ();
 FILLCELL_X4 FILLER_138_1430 ();
 FILLCELL_X2 FILLER_138_1434 ();
 FILLCELL_X2 FILLER_138_1467 ();
 FILLCELL_X2 FILLER_138_1474 ();
 FILLCELL_X1 FILLER_138_1476 ();
 FILLCELL_X4 FILLER_138_1495 ();
 FILLCELL_X8 FILLER_138_1502 ();
 FILLCELL_X1 FILLER_138_1510 ();
 FILLCELL_X4 FILLER_138_1520 ();
 FILLCELL_X2 FILLER_138_1524 ();
 FILLCELL_X1 FILLER_138_1526 ();
 FILLCELL_X4 FILLER_138_1530 ();
 FILLCELL_X2 FILLER_138_1534 ();
 FILLCELL_X1 FILLER_138_1536 ();
 FILLCELL_X32 FILLER_138_1564 ();
 FILLCELL_X32 FILLER_138_1596 ();
 FILLCELL_X16 FILLER_138_1628 ();
 FILLCELL_X4 FILLER_138_1644 ();
 FILLCELL_X2 FILLER_138_1648 ();
 FILLCELL_X1 FILLER_138_1650 ();
 FILLCELL_X8 FILLER_139_1 ();
 FILLCELL_X4 FILLER_139_9 ();
 FILLCELL_X1 FILLER_139_13 ();
 FILLCELL_X4 FILLER_139_33 ();
 FILLCELL_X16 FILLER_139_44 ();
 FILLCELL_X8 FILLER_139_88 ();
 FILLCELL_X2 FILLER_139_96 ();
 FILLCELL_X1 FILLER_139_98 ();
 FILLCELL_X4 FILLER_139_125 ();
 FILLCELL_X1 FILLER_139_129 ();
 FILLCELL_X4 FILLER_139_156 ();
 FILLCELL_X2 FILLER_139_160 ();
 FILLCELL_X1 FILLER_139_169 ();
 FILLCELL_X2 FILLER_139_177 ();
 FILLCELL_X1 FILLER_139_179 ();
 FILLCELL_X4 FILLER_139_207 ();
 FILLCELL_X8 FILLER_139_224 ();
 FILLCELL_X8 FILLER_139_256 ();
 FILLCELL_X4 FILLER_139_264 ();
 FILLCELL_X2 FILLER_139_268 ();
 FILLCELL_X4 FILLER_139_277 ();
 FILLCELL_X1 FILLER_139_281 ();
 FILLCELL_X2 FILLER_139_306 ();
 FILLCELL_X1 FILLER_139_326 ();
 FILLCELL_X1 FILLER_139_347 ();
 FILLCELL_X2 FILLER_139_353 ();
 FILLCELL_X1 FILLER_139_375 ();
 FILLCELL_X8 FILLER_139_399 ();
 FILLCELL_X2 FILLER_139_407 ();
 FILLCELL_X1 FILLER_139_409 ();
 FILLCELL_X1 FILLER_139_418 ();
 FILLCELL_X1 FILLER_139_422 ();
 FILLCELL_X4 FILLER_139_434 ();
 FILLCELL_X2 FILLER_139_445 ();
 FILLCELL_X2 FILLER_139_454 ();
 FILLCELL_X1 FILLER_139_456 ();
 FILLCELL_X1 FILLER_139_462 ();
 FILLCELL_X2 FILLER_139_472 ();
 FILLCELL_X1 FILLER_139_474 ();
 FILLCELL_X8 FILLER_139_484 ();
 FILLCELL_X1 FILLER_139_492 ();
 FILLCELL_X4 FILLER_139_503 ();
 FILLCELL_X2 FILLER_139_507 ();
 FILLCELL_X1 FILLER_139_509 ();
 FILLCELL_X2 FILLER_139_517 ();
 FILLCELL_X2 FILLER_139_522 ();
 FILLCELL_X1 FILLER_139_524 ();
 FILLCELL_X2 FILLER_139_529 ();
 FILLCELL_X1 FILLER_139_531 ();
 FILLCELL_X8 FILLER_139_535 ();
 FILLCELL_X2 FILLER_139_543 ();
 FILLCELL_X16 FILLER_139_568 ();
 FILLCELL_X1 FILLER_139_605 ();
 FILLCELL_X1 FILLER_139_615 ();
 FILLCELL_X1 FILLER_139_620 ();
 FILLCELL_X1 FILLER_139_624 ();
 FILLCELL_X4 FILLER_139_664 ();
 FILLCELL_X1 FILLER_139_668 ();
 FILLCELL_X1 FILLER_139_673 ();
 FILLCELL_X1 FILLER_139_677 ();
 FILLCELL_X2 FILLER_139_681 ();
 FILLCELL_X1 FILLER_139_686 ();
 FILLCELL_X1 FILLER_139_694 ();
 FILLCELL_X2 FILLER_139_722 ();
 FILLCELL_X2 FILLER_139_733 ();
 FILLCELL_X16 FILLER_139_742 ();
 FILLCELL_X2 FILLER_139_758 ();
 FILLCELL_X1 FILLER_139_760 ();
 FILLCELL_X8 FILLER_139_781 ();
 FILLCELL_X4 FILLER_139_789 ();
 FILLCELL_X1 FILLER_139_793 ();
 FILLCELL_X2 FILLER_139_801 ();
 FILLCELL_X4 FILLER_139_810 ();
 FILLCELL_X1 FILLER_139_814 ();
 FILLCELL_X8 FILLER_139_818 ();
 FILLCELL_X4 FILLER_139_862 ();
 FILLCELL_X1 FILLER_139_866 ();
 FILLCELL_X8 FILLER_139_874 ();
 FILLCELL_X8 FILLER_139_895 ();
 FILLCELL_X8 FILLER_139_908 ();
 FILLCELL_X2 FILLER_139_916 ();
 FILLCELL_X1 FILLER_139_918 ();
 FILLCELL_X1 FILLER_139_994 ();
 FILLCELL_X16 FILLER_139_1056 ();
 FILLCELL_X2 FILLER_139_1072 ();
 FILLCELL_X4 FILLER_139_1082 ();
 FILLCELL_X1 FILLER_139_1086 ();
 FILLCELL_X8 FILLER_139_1097 ();
 FILLCELL_X2 FILLER_139_1144 ();
 FILLCELL_X2 FILLER_139_1152 ();
 FILLCELL_X1 FILLER_139_1160 ();
 FILLCELL_X8 FILLER_139_1167 ();
 FILLCELL_X2 FILLER_139_1175 ();
 FILLCELL_X1 FILLER_139_1177 ();
 FILLCELL_X4 FILLER_139_1194 ();
 FILLCELL_X2 FILLER_139_1198 ();
 FILLCELL_X1 FILLER_139_1200 ();
 FILLCELL_X2 FILLER_139_1211 ();
 FILLCELL_X1 FILLER_139_1213 ();
 FILLCELL_X1 FILLER_139_1224 ();
 FILLCELL_X2 FILLER_139_1251 ();
 FILLCELL_X1 FILLER_139_1264 ();
 FILLCELL_X1 FILLER_139_1275 ();
 FILLCELL_X32 FILLER_139_1309 ();
 FILLCELL_X16 FILLER_139_1341 ();
 FILLCELL_X8 FILLER_139_1357 ();
 FILLCELL_X1 FILLER_139_1365 ();
 FILLCELL_X4 FILLER_139_1384 ();
 FILLCELL_X1 FILLER_139_1388 ();
 FILLCELL_X2 FILLER_139_1406 ();
 FILLCELL_X4 FILLER_139_1412 ();
 FILLCELL_X2 FILLER_139_1416 ();
 FILLCELL_X1 FILLER_139_1418 ();
 FILLCELL_X8 FILLER_139_1458 ();
 FILLCELL_X2 FILLER_139_1466 ();
 FILLCELL_X1 FILLER_139_1468 ();
 FILLCELL_X4 FILLER_139_1473 ();
 FILLCELL_X1 FILLER_139_1477 ();
 FILLCELL_X4 FILLER_139_1514 ();
 FILLCELL_X2 FILLER_139_1518 ();
 FILLCELL_X1 FILLER_139_1520 ();
 FILLCELL_X2 FILLER_139_1524 ();
 FILLCELL_X2 FILLER_139_1535 ();
 FILLCELL_X4 FILLER_139_1558 ();
 FILLCELL_X1 FILLER_139_1562 ();
 FILLCELL_X32 FILLER_139_1572 ();
 FILLCELL_X32 FILLER_139_1604 ();
 FILLCELL_X8 FILLER_139_1636 ();
 FILLCELL_X4 FILLER_139_1644 ();
 FILLCELL_X2 FILLER_139_1648 ();
 FILLCELL_X1 FILLER_139_1650 ();
 FILLCELL_X16 FILLER_140_1 ();
 FILLCELL_X2 FILLER_140_17 ();
 FILLCELL_X1 FILLER_140_39 ();
 FILLCELL_X2 FILLER_140_47 ();
 FILLCELL_X4 FILLER_140_56 ();
 FILLCELL_X2 FILLER_140_60 ();
 FILLCELL_X1 FILLER_140_66 ();
 FILLCELL_X1 FILLER_140_95 ();
 FILLCELL_X1 FILLER_140_123 ();
 FILLCELL_X2 FILLER_140_144 ();
 FILLCELL_X1 FILLER_140_146 ();
 FILLCELL_X2 FILLER_140_160 ();
 FILLCELL_X1 FILLER_140_162 ();
 FILLCELL_X2 FILLER_140_170 ();
 FILLCELL_X1 FILLER_140_172 ();
 FILLCELL_X2 FILLER_140_222 ();
 FILLCELL_X1 FILLER_140_224 ();
 FILLCELL_X4 FILLER_140_245 ();
 FILLCELL_X2 FILLER_140_249 ();
 FILLCELL_X1 FILLER_140_251 ();
 FILLCELL_X4 FILLER_140_255 ();
 FILLCELL_X1 FILLER_140_259 ();
 FILLCELL_X2 FILLER_140_287 ();
 FILLCELL_X1 FILLER_140_289 ();
 FILLCELL_X2 FILLER_140_310 ();
 FILLCELL_X1 FILLER_140_332 ();
 FILLCELL_X2 FILLER_140_359 ();
 FILLCELL_X1 FILLER_140_361 ();
 FILLCELL_X4 FILLER_140_366 ();
 FILLCELL_X2 FILLER_140_370 ();
 FILLCELL_X2 FILLER_140_375 ();
 FILLCELL_X1 FILLER_140_377 ();
 FILLCELL_X4 FILLER_140_382 ();
 FILLCELL_X2 FILLER_140_386 ();
 FILLCELL_X4 FILLER_140_402 ();
 FILLCELL_X1 FILLER_140_406 ();
 FILLCELL_X8 FILLER_140_441 ();
 FILLCELL_X1 FILLER_140_481 ();
 FILLCELL_X1 FILLER_140_522 ();
 FILLCELL_X2 FILLER_140_553 ();
 FILLCELL_X2 FILLER_140_575 ();
 FILLCELL_X1 FILLER_140_577 ();
 FILLCELL_X1 FILLER_140_598 ();
 FILLCELL_X2 FILLER_140_603 ();
 FILLCELL_X1 FILLER_140_605 ();
 FILLCELL_X1 FILLER_140_609 ();
 FILLCELL_X8 FILLER_140_613 ();
 FILLCELL_X4 FILLER_140_621 ();
 FILLCELL_X1 FILLER_140_625 ();
 FILLCELL_X16 FILLER_140_632 ();
 FILLCELL_X2 FILLER_140_648 ();
 FILLCELL_X1 FILLER_140_650 ();
 FILLCELL_X16 FILLER_140_658 ();
 FILLCELL_X8 FILLER_140_674 ();
 FILLCELL_X1 FILLER_140_682 ();
 FILLCELL_X1 FILLER_140_776 ();
 FILLCELL_X1 FILLER_140_797 ();
 FILLCELL_X2 FILLER_140_807 ();
 FILLCELL_X1 FILLER_140_809 ();
 FILLCELL_X8 FILLER_140_838 ();
 FILLCELL_X4 FILLER_140_846 ();
 FILLCELL_X2 FILLER_140_850 ();
 FILLCELL_X1 FILLER_140_852 ();
 FILLCELL_X8 FILLER_140_860 ();
 FILLCELL_X1 FILLER_140_868 ();
 FILLCELL_X4 FILLER_140_885 ();
 FILLCELL_X2 FILLER_140_889 ();
 FILLCELL_X1 FILLER_140_891 ();
 FILLCELL_X2 FILLER_140_899 ();
 FILLCELL_X4 FILLER_140_921 ();
 FILLCELL_X8 FILLER_140_942 ();
 FILLCELL_X4 FILLER_140_950 ();
 FILLCELL_X2 FILLER_140_954 ();
 FILLCELL_X8 FILLER_140_959 ();
 FILLCELL_X4 FILLER_140_967 ();
 FILLCELL_X2 FILLER_140_971 ();
 FILLCELL_X1 FILLER_140_973 ();
 FILLCELL_X4 FILLER_140_981 ();
 FILLCELL_X16 FILLER_140_1012 ();
 FILLCELL_X4 FILLER_140_1028 ();
 FILLCELL_X2 FILLER_140_1032 ();
 FILLCELL_X1 FILLER_140_1034 ();
 FILLCELL_X4 FILLER_140_1042 ();
 FILLCELL_X2 FILLER_140_1046 ();
 FILLCELL_X1 FILLER_140_1048 ();
 FILLCELL_X16 FILLER_140_1054 ();
 FILLCELL_X8 FILLER_140_1070 ();
 FILLCELL_X2 FILLER_140_1078 ();
 FILLCELL_X1 FILLER_140_1080 ();
 FILLCELL_X2 FILLER_140_1091 ();
 FILLCELL_X1 FILLER_140_1093 ();
 FILLCELL_X1 FILLER_140_1104 ();
 FILLCELL_X4 FILLER_140_1121 ();
 FILLCELL_X16 FILLER_140_1159 ();
 FILLCELL_X1 FILLER_140_1175 ();
 FILLCELL_X1 FILLER_140_1182 ();
 FILLCELL_X1 FILLER_140_1193 ();
 FILLCELL_X1 FILLER_140_1204 ();
 FILLCELL_X4 FILLER_140_1221 ();
 FILLCELL_X2 FILLER_140_1234 ();
 FILLCELL_X1 FILLER_140_1236 ();
 FILLCELL_X2 FILLER_140_1255 ();
 FILLCELL_X1 FILLER_140_1272 ();
 FILLCELL_X1 FILLER_140_1298 ();
 FILLCELL_X32 FILLER_140_1305 ();
 FILLCELL_X32 FILLER_140_1337 ();
 FILLCELL_X8 FILLER_140_1369 ();
 FILLCELL_X4 FILLER_140_1377 ();
 FILLCELL_X1 FILLER_140_1381 ();
 FILLCELL_X2 FILLER_140_1394 ();
 FILLCELL_X2 FILLER_140_1405 ();
 FILLCELL_X2 FILLER_140_1427 ();
 FILLCELL_X4 FILLER_140_1436 ();
 FILLCELL_X2 FILLER_140_1440 ();
 FILLCELL_X2 FILLER_140_1449 ();
 FILLCELL_X2 FILLER_140_1455 ();
 FILLCELL_X1 FILLER_140_1484 ();
 FILLCELL_X2 FILLER_140_1488 ();
 FILLCELL_X4 FILLER_140_1500 ();
 FILLCELL_X2 FILLER_140_1504 ();
 FILLCELL_X2 FILLER_140_1520 ();
 FILLCELL_X8 FILLER_140_1531 ();
 FILLCELL_X2 FILLER_140_1539 ();
 FILLCELL_X1 FILLER_140_1541 ();
 FILLCELL_X2 FILLER_140_1549 ();
 FILLCELL_X2 FILLER_140_1558 ();
 FILLCELL_X32 FILLER_140_1567 ();
 FILLCELL_X32 FILLER_140_1599 ();
 FILLCELL_X16 FILLER_140_1631 ();
 FILLCELL_X4 FILLER_140_1647 ();
 FILLCELL_X16 FILLER_141_1 ();
 FILLCELL_X2 FILLER_141_17 ();
 FILLCELL_X1 FILLER_141_39 ();
 FILLCELL_X2 FILLER_141_47 ();
 FILLCELL_X2 FILLER_141_73 ();
 FILLCELL_X1 FILLER_141_75 ();
 FILLCELL_X2 FILLER_141_94 ();
 FILLCELL_X1 FILLER_141_96 ();
 FILLCELL_X8 FILLER_141_110 ();
 FILLCELL_X2 FILLER_141_118 ();
 FILLCELL_X16 FILLER_141_148 ();
 FILLCELL_X2 FILLER_141_164 ();
 FILLCELL_X1 FILLER_141_186 ();
 FILLCELL_X1 FILLER_141_207 ();
 FILLCELL_X4 FILLER_141_213 ();
 FILLCELL_X2 FILLER_141_217 ();
 FILLCELL_X1 FILLER_141_226 ();
 FILLCELL_X1 FILLER_141_254 ();
 FILLCELL_X8 FILLER_141_284 ();
 FILLCELL_X8 FILLER_141_296 ();
 FILLCELL_X2 FILLER_141_304 ();
 FILLCELL_X2 FILLER_141_318 ();
 FILLCELL_X1 FILLER_141_340 ();
 FILLCELL_X2 FILLER_141_346 ();
 FILLCELL_X1 FILLER_141_348 ();
 FILLCELL_X4 FILLER_141_358 ();
 FILLCELL_X2 FILLER_141_362 ();
 FILLCELL_X1 FILLER_141_364 ();
 FILLCELL_X2 FILLER_141_401 ();
 FILLCELL_X1 FILLER_141_403 ();
 FILLCELL_X1 FILLER_141_413 ();
 FILLCELL_X8 FILLER_141_421 ();
 FILLCELL_X4 FILLER_141_429 ();
 FILLCELL_X1 FILLER_141_433 ();
 FILLCELL_X8 FILLER_141_441 ();
 FILLCELL_X1 FILLER_141_472 ();
 FILLCELL_X1 FILLER_141_477 ();
 FILLCELL_X8 FILLER_141_483 ();
 FILLCELL_X1 FILLER_141_491 ();
 FILLCELL_X2 FILLER_141_507 ();
 FILLCELL_X1 FILLER_141_509 ();
 FILLCELL_X1 FILLER_141_556 ();
 FILLCELL_X4 FILLER_141_628 ();
 FILLCELL_X2 FILLER_141_632 ();
 FILLCELL_X4 FILLER_141_654 ();
 FILLCELL_X2 FILLER_141_658 ();
 FILLCELL_X1 FILLER_141_660 ();
 FILLCELL_X1 FILLER_141_665 ();
 FILLCELL_X1 FILLER_141_670 ();
 FILLCELL_X4 FILLER_141_674 ();
 FILLCELL_X2 FILLER_141_678 ();
 FILLCELL_X1 FILLER_141_680 ();
 FILLCELL_X2 FILLER_141_685 ();
 FILLCELL_X1 FILLER_141_687 ();
 FILLCELL_X8 FILLER_141_692 ();
 FILLCELL_X4 FILLER_141_700 ();
 FILLCELL_X2 FILLER_141_704 ();
 FILLCELL_X2 FILLER_141_726 ();
 FILLCELL_X2 FILLER_141_760 ();
 FILLCELL_X1 FILLER_141_762 ();
 FILLCELL_X1 FILLER_141_770 ();
 FILLCELL_X2 FILLER_141_805 ();
 FILLCELL_X2 FILLER_141_827 ();
 FILLCELL_X1 FILLER_141_829 ();
 FILLCELL_X4 FILLER_141_839 ();
 FILLCELL_X1 FILLER_141_843 ();
 FILLCELL_X2 FILLER_141_864 ();
 FILLCELL_X4 FILLER_141_886 ();
 FILLCELL_X1 FILLER_141_890 ();
 FILLCELL_X8 FILLER_141_911 ();
 FILLCELL_X4 FILLER_141_919 ();
 FILLCELL_X1 FILLER_141_923 ();
 FILLCELL_X16 FILLER_141_937 ();
 FILLCELL_X4 FILLER_141_953 ();
 FILLCELL_X2 FILLER_141_957 ();
 FILLCELL_X1 FILLER_141_959 ();
 FILLCELL_X8 FILLER_141_964 ();
 FILLCELL_X1 FILLER_141_972 ();
 FILLCELL_X2 FILLER_141_993 ();
 FILLCELL_X1 FILLER_141_995 ();
 FILLCELL_X16 FILLER_141_1023 ();
 FILLCELL_X8 FILLER_141_1076 ();
 FILLCELL_X4 FILLER_141_1084 ();
 FILLCELL_X2 FILLER_141_1088 ();
 FILLCELL_X2 FILLER_141_1112 ();
 FILLCELL_X1 FILLER_141_1114 ();
 FILLCELL_X1 FILLER_141_1131 ();
 FILLCELL_X1 FILLER_141_1142 ();
 FILLCELL_X8 FILLER_141_1161 ();
 FILLCELL_X4 FILLER_141_1169 ();
 FILLCELL_X2 FILLER_141_1183 ();
 FILLCELL_X2 FILLER_141_1195 ();
 FILLCELL_X8 FILLER_141_1203 ();
 FILLCELL_X1 FILLER_141_1211 ();
 FILLCELL_X8 FILLER_141_1222 ();
 FILLCELL_X2 FILLER_141_1230 ();
 FILLCELL_X1 FILLER_141_1232 ();
 FILLCELL_X2 FILLER_141_1245 ();
 FILLCELL_X8 FILLER_141_1264 ();
 FILLCELL_X1 FILLER_141_1272 ();
 FILLCELL_X4 FILLER_141_1283 ();
 FILLCELL_X4 FILLER_141_1315 ();
 FILLCELL_X2 FILLER_141_1319 ();
 FILLCELL_X32 FILLER_141_1328 ();
 FILLCELL_X16 FILLER_141_1360 ();
 FILLCELL_X2 FILLER_141_1376 ();
 FILLCELL_X4 FILLER_141_1387 ();
 FILLCELL_X2 FILLER_141_1391 ();
 FILLCELL_X4 FILLER_141_1398 ();
 FILLCELL_X2 FILLER_141_1402 ();
 FILLCELL_X1 FILLER_141_1404 ();
 FILLCELL_X4 FILLER_141_1416 ();
 FILLCELL_X2 FILLER_141_1420 ();
 FILLCELL_X2 FILLER_141_1429 ();
 FILLCELL_X1 FILLER_141_1431 ();
 FILLCELL_X1 FILLER_141_1440 ();
 FILLCELL_X2 FILLER_141_1453 ();
 FILLCELL_X4 FILLER_141_1466 ();
 FILLCELL_X2 FILLER_141_1470 ();
 FILLCELL_X1 FILLER_141_1483 ();
 FILLCELL_X4 FILLER_141_1495 ();
 FILLCELL_X2 FILLER_141_1499 ();
 FILLCELL_X1 FILLER_141_1501 ();
 FILLCELL_X4 FILLER_141_1509 ();
 FILLCELL_X4 FILLER_141_1537 ();
 FILLCELL_X4 FILLER_141_1556 ();
 FILLCELL_X4 FILLER_141_1564 ();
 FILLCELL_X2 FILLER_141_1568 ();
 FILLCELL_X32 FILLER_141_1577 ();
 FILLCELL_X32 FILLER_141_1609 ();
 FILLCELL_X8 FILLER_141_1641 ();
 FILLCELL_X2 FILLER_141_1649 ();
 FILLCELL_X2 FILLER_142_1 ();
 FILLCELL_X1 FILLER_142_3 ();
 FILLCELL_X4 FILLER_142_24 ();
 FILLCELL_X2 FILLER_142_28 ();
 FILLCELL_X2 FILLER_142_37 ();
 FILLCELL_X1 FILLER_142_39 ();
 FILLCELL_X8 FILLER_142_45 ();
 FILLCELL_X4 FILLER_142_53 ();
 FILLCELL_X1 FILLER_142_57 ();
 FILLCELL_X2 FILLER_142_83 ();
 FILLCELL_X8 FILLER_142_106 ();
 FILLCELL_X2 FILLER_142_114 ();
 FILLCELL_X1 FILLER_142_123 ();
 FILLCELL_X2 FILLER_142_138 ();
 FILLCELL_X4 FILLER_142_160 ();
 FILLCELL_X2 FILLER_142_164 ();
 FILLCELL_X1 FILLER_142_166 ();
 FILLCELL_X2 FILLER_142_174 ();
 FILLCELL_X1 FILLER_142_176 ();
 FILLCELL_X4 FILLER_142_184 ();
 FILLCELL_X4 FILLER_142_213 ();
 FILLCELL_X2 FILLER_142_217 ();
 FILLCELL_X2 FILLER_142_226 ();
 FILLCELL_X4 FILLER_142_230 ();
 FILLCELL_X1 FILLER_142_234 ();
 FILLCELL_X4 FILLER_142_263 ();
 FILLCELL_X8 FILLER_142_281 ();
 FILLCELL_X4 FILLER_142_289 ();
 FILLCELL_X4 FILLER_142_300 ();
 FILLCELL_X2 FILLER_142_304 ();
 FILLCELL_X1 FILLER_142_306 ();
 FILLCELL_X4 FILLER_142_314 ();
 FILLCELL_X1 FILLER_142_318 ();
 FILLCELL_X4 FILLER_142_322 ();
 FILLCELL_X2 FILLER_142_326 ();
 FILLCELL_X4 FILLER_142_335 ();
 FILLCELL_X1 FILLER_142_339 ();
 FILLCELL_X4 FILLER_142_349 ();
 FILLCELL_X2 FILLER_142_353 ();
 FILLCELL_X1 FILLER_142_359 ();
 FILLCELL_X4 FILLER_142_363 ();
 FILLCELL_X2 FILLER_142_367 ();
 FILLCELL_X8 FILLER_142_373 ();
 FILLCELL_X1 FILLER_142_381 ();
 FILLCELL_X8 FILLER_142_392 ();
 FILLCELL_X2 FILLER_142_404 ();
 FILLCELL_X1 FILLER_142_406 ();
 FILLCELL_X2 FILLER_142_433 ();
 FILLCELL_X2 FILLER_142_456 ();
 FILLCELL_X4 FILLER_142_465 ();
 FILLCELL_X2 FILLER_142_469 ();
 FILLCELL_X1 FILLER_142_471 ();
 FILLCELL_X2 FILLER_142_479 ();
 FILLCELL_X1 FILLER_142_488 ();
 FILLCELL_X2 FILLER_142_496 ();
 FILLCELL_X1 FILLER_142_498 ();
 FILLCELL_X4 FILLER_142_513 ();
 FILLCELL_X2 FILLER_142_521 ();
 FILLCELL_X1 FILLER_142_523 ();
 FILLCELL_X2 FILLER_142_527 ();
 FILLCELL_X1 FILLER_142_529 ();
 FILLCELL_X4 FILLER_142_534 ();
 FILLCELL_X1 FILLER_142_538 ();
 FILLCELL_X1 FILLER_142_543 ();
 FILLCELL_X8 FILLER_142_550 ();
 FILLCELL_X4 FILLER_142_558 ();
 FILLCELL_X1 FILLER_142_562 ();
 FILLCELL_X2 FILLER_142_567 ();
 FILLCELL_X4 FILLER_142_572 ();
 FILLCELL_X2 FILLER_142_581 ();
 FILLCELL_X2 FILLER_142_587 ();
 FILLCELL_X2 FILLER_142_593 ();
 FILLCELL_X8 FILLER_142_598 ();
 FILLCELL_X2 FILLER_142_606 ();
 FILLCELL_X4 FILLER_142_632 ();
 FILLCELL_X4 FILLER_142_643 ();
 FILLCELL_X1 FILLER_142_650 ();
 FILLCELL_X4 FILLER_142_656 ();
 FILLCELL_X2 FILLER_142_660 ();
 FILLCELL_X1 FILLER_142_693 ();
 FILLCELL_X4 FILLER_142_696 ();
 FILLCELL_X2 FILLER_142_700 ();
 FILLCELL_X1 FILLER_142_702 ();
 FILLCELL_X4 FILLER_142_710 ();
 FILLCELL_X1 FILLER_142_714 ();
 FILLCELL_X4 FILLER_142_720 ();
 FILLCELL_X1 FILLER_142_731 ();
 FILLCELL_X2 FILLER_142_766 ();
 FILLCELL_X1 FILLER_142_768 ();
 FILLCELL_X4 FILLER_142_776 ();
 FILLCELL_X1 FILLER_142_780 ();
 FILLCELL_X2 FILLER_142_790 ();
 FILLCELL_X4 FILLER_142_799 ();
 FILLCELL_X4 FILLER_142_806 ();
 FILLCELL_X4 FILLER_142_830 ();
 FILLCELL_X4 FILLER_142_908 ();
 FILLCELL_X1 FILLER_142_912 ();
 FILLCELL_X2 FILLER_142_926 ();
 FILLCELL_X4 FILLER_142_931 ();
 FILLCELL_X8 FILLER_142_966 ();
 FILLCELL_X2 FILLER_142_981 ();
 FILLCELL_X1 FILLER_142_996 ();
 FILLCELL_X1 FILLER_142_1044 ();
 FILLCELL_X2 FILLER_142_1051 ();
 FILLCELL_X1 FILLER_142_1053 ();
 FILLCELL_X1 FILLER_142_1061 ();
 FILLCELL_X4 FILLER_142_1082 ();
 FILLCELL_X1 FILLER_142_1086 ();
 FILLCELL_X4 FILLER_142_1097 ();
 FILLCELL_X2 FILLER_142_1101 ();
 FILLCELL_X2 FILLER_142_1119 ();
 FILLCELL_X2 FILLER_142_1131 ();
 FILLCELL_X4 FILLER_142_1139 ();
 FILLCELL_X2 FILLER_142_1149 ();
 FILLCELL_X2 FILLER_142_1157 ();
 FILLCELL_X1 FILLER_142_1159 ();
 FILLCELL_X2 FILLER_142_1170 ();
 FILLCELL_X1 FILLER_142_1172 ();
 FILLCELL_X2 FILLER_142_1179 ();
 FILLCELL_X2 FILLER_142_1197 ();
 FILLCELL_X1 FILLER_142_1199 ();
 FILLCELL_X1 FILLER_142_1206 ();
 FILLCELL_X2 FILLER_142_1235 ();
 FILLCELL_X4 FILLER_142_1243 ();
 FILLCELL_X1 FILLER_142_1247 ();
 FILLCELL_X1 FILLER_142_1264 ();
 FILLCELL_X1 FILLER_142_1275 ();
 FILLCELL_X1 FILLER_142_1282 ();
 FILLCELL_X16 FILLER_142_1295 ();
 FILLCELL_X32 FILLER_142_1335 ();
 FILLCELL_X8 FILLER_142_1367 ();
 FILLCELL_X1 FILLER_142_1397 ();
 FILLCELL_X4 FILLER_142_1407 ();
 FILLCELL_X1 FILLER_142_1416 ();
 FILLCELL_X2 FILLER_142_1420 ();
 FILLCELL_X1 FILLER_142_1422 ();
 FILLCELL_X16 FILLER_142_1433 ();
 FILLCELL_X1 FILLER_142_1449 ();
 FILLCELL_X2 FILLER_142_1480 ();
 FILLCELL_X16 FILLER_142_1485 ();
 FILLCELL_X2 FILLER_142_1501 ();
 FILLCELL_X2 FILLER_142_1507 ();
 FILLCELL_X1 FILLER_142_1509 ();
 FILLCELL_X8 FILLER_142_1522 ();
 FILLCELL_X1 FILLER_142_1530 ();
 FILLCELL_X4 FILLER_142_1535 ();
 FILLCELL_X2 FILLER_142_1539 ();
 FILLCELL_X1 FILLER_142_1541 ();
 FILLCELL_X8 FILLER_142_1561 ();
 FILLCELL_X4 FILLER_142_1569 ();
 FILLCELL_X1 FILLER_142_1573 ();
 FILLCELL_X2 FILLER_142_1578 ();
 FILLCELL_X1 FILLER_142_1580 ();
 FILLCELL_X32 FILLER_142_1592 ();
 FILLCELL_X16 FILLER_142_1624 ();
 FILLCELL_X8 FILLER_142_1640 ();
 FILLCELL_X2 FILLER_142_1648 ();
 FILLCELL_X1 FILLER_142_1650 ();
 FILLCELL_X8 FILLER_143_1 ();
 FILLCELL_X4 FILLER_143_9 ();
 FILLCELL_X8 FILLER_143_67 ();
 FILLCELL_X4 FILLER_143_82 ();
 FILLCELL_X2 FILLER_143_86 ();
 FILLCELL_X2 FILLER_143_135 ();
 FILLCELL_X8 FILLER_143_157 ();
 FILLCELL_X4 FILLER_143_165 ();
 FILLCELL_X2 FILLER_143_169 ();
 FILLCELL_X8 FILLER_143_178 ();
 FILLCELL_X1 FILLER_143_199 ();
 FILLCELL_X8 FILLER_143_256 ();
 FILLCELL_X4 FILLER_143_264 ();
 FILLCELL_X1 FILLER_143_268 ();
 FILLCELL_X2 FILLER_143_278 ();
 FILLCELL_X2 FILLER_143_300 ();
 FILLCELL_X4 FILLER_143_322 ();
 FILLCELL_X1 FILLER_143_350 ();
 FILLCELL_X2 FILLER_143_371 ();
 FILLCELL_X2 FILLER_143_393 ();
 FILLCELL_X2 FILLER_143_415 ();
 FILLCELL_X8 FILLER_143_446 ();
 FILLCELL_X2 FILLER_143_454 ();
 FILLCELL_X8 FILLER_143_463 ();
 FILLCELL_X4 FILLER_143_471 ();
 FILLCELL_X2 FILLER_143_475 ();
 FILLCELL_X4 FILLER_143_484 ();
 FILLCELL_X2 FILLER_143_488 ();
 FILLCELL_X1 FILLER_143_490 ();
 FILLCELL_X2 FILLER_143_512 ();
 FILLCELL_X1 FILLER_143_521 ();
 FILLCELL_X2 FILLER_143_526 ();
 FILLCELL_X1 FILLER_143_528 ();
 FILLCELL_X1 FILLER_143_549 ();
 FILLCELL_X8 FILLER_143_557 ();
 FILLCELL_X4 FILLER_143_565 ();
 FILLCELL_X2 FILLER_143_569 ();
 FILLCELL_X1 FILLER_143_571 ();
 FILLCELL_X4 FILLER_143_586 ();
 FILLCELL_X2 FILLER_143_590 ();
 FILLCELL_X1 FILLER_143_612 ();
 FILLCELL_X1 FILLER_143_617 ();
 FILLCELL_X4 FILLER_143_621 ();
 FILLCELL_X1 FILLER_143_625 ();
 FILLCELL_X4 FILLER_143_650 ();
 FILLCELL_X4 FILLER_143_661 ();
 FILLCELL_X1 FILLER_143_665 ();
 FILLCELL_X2 FILLER_143_670 ();
 FILLCELL_X1 FILLER_143_677 ();
 FILLCELL_X8 FILLER_143_752 ();
 FILLCELL_X2 FILLER_143_760 ();
 FILLCELL_X1 FILLER_143_762 ();
 FILLCELL_X8 FILLER_143_823 ();
 FILLCELL_X4 FILLER_143_831 ();
 FILLCELL_X2 FILLER_143_885 ();
 FILLCELL_X2 FILLER_143_923 ();
 FILLCELL_X1 FILLER_143_929 ();
 FILLCELL_X4 FILLER_143_937 ();
 FILLCELL_X2 FILLER_143_961 ();
 FILLCELL_X2 FILLER_143_972 ();
 FILLCELL_X1 FILLER_143_974 ();
 FILLCELL_X16 FILLER_143_982 ();
 FILLCELL_X2 FILLER_143_998 ();
 FILLCELL_X8 FILLER_143_1016 ();
 FILLCELL_X1 FILLER_143_1032 ();
 FILLCELL_X2 FILLER_143_1037 ();
 FILLCELL_X1 FILLER_143_1039 ();
 FILLCELL_X1 FILLER_143_1045 ();
 FILLCELL_X2 FILLER_143_1057 ();
 FILLCELL_X1 FILLER_143_1059 ();
 FILLCELL_X4 FILLER_143_1074 ();
 FILLCELL_X2 FILLER_143_1078 ();
 FILLCELL_X4 FILLER_143_1092 ();
 FILLCELL_X2 FILLER_143_1106 ();
 FILLCELL_X1 FILLER_143_1108 ();
 FILLCELL_X1 FILLER_143_1125 ();
 FILLCELL_X4 FILLER_143_1142 ();
 FILLCELL_X1 FILLER_143_1146 ();
 FILLCELL_X8 FILLER_143_1165 ();
 FILLCELL_X4 FILLER_143_1179 ();
 FILLCELL_X2 FILLER_143_1183 ();
 FILLCELL_X4 FILLER_143_1191 ();
 FILLCELL_X2 FILLER_143_1195 ();
 FILLCELL_X16 FILLER_143_1207 ();
 FILLCELL_X2 FILLER_143_1229 ();
 FILLCELL_X1 FILLER_143_1255 ();
 FILLCELL_X1 FILLER_143_1262 ();
 FILLCELL_X16 FILLER_143_1286 ();
 FILLCELL_X8 FILLER_143_1302 ();
 FILLCELL_X32 FILLER_143_1330 ();
 FILLCELL_X4 FILLER_143_1362 ();
 FILLCELL_X1 FILLER_143_1366 ();
 FILLCELL_X8 FILLER_143_1380 ();
 FILLCELL_X2 FILLER_143_1388 ();
 FILLCELL_X1 FILLER_143_1396 ();
 FILLCELL_X1 FILLER_143_1409 ();
 FILLCELL_X2 FILLER_143_1449 ();
 FILLCELL_X1 FILLER_143_1455 ();
 FILLCELL_X2 FILLER_143_1461 ();
 FILLCELL_X1 FILLER_143_1477 ();
 FILLCELL_X16 FILLER_143_1489 ();
 FILLCELL_X2 FILLER_143_1505 ();
 FILLCELL_X1 FILLER_143_1507 ();
 FILLCELL_X2 FILLER_143_1512 ();
 FILLCELL_X1 FILLER_143_1527 ();
 FILLCELL_X1 FILLER_143_1533 ();
 FILLCELL_X1 FILLER_143_1541 ();
 FILLCELL_X1 FILLER_143_1551 ();
 FILLCELL_X2 FILLER_143_1559 ();
 FILLCELL_X4 FILLER_143_1576 ();
 FILLCELL_X2 FILLER_143_1580 ();
 FILLCELL_X1 FILLER_143_1582 ();
 FILLCELL_X32 FILLER_143_1585 ();
 FILLCELL_X32 FILLER_143_1617 ();
 FILLCELL_X2 FILLER_143_1649 ();
 FILLCELL_X16 FILLER_144_1 ();
 FILLCELL_X8 FILLER_144_17 ();
 FILLCELL_X1 FILLER_144_25 ();
 FILLCELL_X4 FILLER_144_33 ();
 FILLCELL_X1 FILLER_144_37 ();
 FILLCELL_X16 FILLER_144_114 ();
 FILLCELL_X8 FILLER_144_130 ();
 FILLCELL_X1 FILLER_144_138 ();
 FILLCELL_X4 FILLER_144_155 ();
 FILLCELL_X2 FILLER_144_159 ();
 FILLCELL_X8 FILLER_144_201 ();
 FILLCELL_X2 FILLER_144_209 ();
 FILLCELL_X1 FILLER_144_236 ();
 FILLCELL_X8 FILLER_144_239 ();
 FILLCELL_X4 FILLER_144_247 ();
 FILLCELL_X2 FILLER_144_251 ();
 FILLCELL_X4 FILLER_144_293 ();
 FILLCELL_X1 FILLER_144_329 ();
 FILLCELL_X8 FILLER_144_359 ();
 FILLCELL_X8 FILLER_144_392 ();
 FILLCELL_X1 FILLER_144_400 ();
 FILLCELL_X2 FILLER_144_407 ();
 FILLCELL_X1 FILLER_144_409 ();
 FILLCELL_X4 FILLER_144_415 ();
 FILLCELL_X2 FILLER_144_419 ();
 FILLCELL_X8 FILLER_144_425 ();
 FILLCELL_X16 FILLER_144_436 ();
 FILLCELL_X2 FILLER_144_452 ();
 FILLCELL_X1 FILLER_144_461 ();
 FILLCELL_X1 FILLER_144_476 ();
 FILLCELL_X2 FILLER_144_498 ();
 FILLCELL_X2 FILLER_144_507 ();
 FILLCELL_X1 FILLER_144_509 ();
 FILLCELL_X2 FILLER_144_568 ();
 FILLCELL_X4 FILLER_144_590 ();
 FILLCELL_X1 FILLER_144_632 ();
 FILLCELL_X2 FILLER_144_636 ();
 FILLCELL_X1 FILLER_144_638 ();
 FILLCELL_X1 FILLER_144_660 ();
 FILLCELL_X2 FILLER_144_681 ();
 FILLCELL_X8 FILLER_144_710 ();
 FILLCELL_X1 FILLER_144_725 ();
 FILLCELL_X16 FILLER_144_766 ();
 FILLCELL_X2 FILLER_144_782 ();
 FILLCELL_X8 FILLER_144_791 ();
 FILLCELL_X1 FILLER_144_799 ();
 FILLCELL_X2 FILLER_144_814 ();
 FILLCELL_X1 FILLER_144_816 ();
 FILLCELL_X8 FILLER_144_826 ();
 FILLCELL_X1 FILLER_144_834 ();
 FILLCELL_X8 FILLER_144_848 ();
 FILLCELL_X4 FILLER_144_856 ();
 FILLCELL_X2 FILLER_144_860 ();
 FILLCELL_X4 FILLER_144_875 ();
 FILLCELL_X4 FILLER_144_933 ();
 FILLCELL_X1 FILLER_144_937 ();
 FILLCELL_X8 FILLER_144_945 ();
 FILLCELL_X4 FILLER_144_953 ();
 FILLCELL_X2 FILLER_144_957 ();
 FILLCELL_X4 FILLER_144_999 ();
 FILLCELL_X2 FILLER_144_1003 ();
 FILLCELL_X1 FILLER_144_1025 ();
 FILLCELL_X8 FILLER_144_1030 ();
 FILLCELL_X1 FILLER_144_1038 ();
 FILLCELL_X2 FILLER_144_1051 ();
 FILLCELL_X1 FILLER_144_1093 ();
 FILLCELL_X2 FILLER_144_1125 ();
 FILLCELL_X1 FILLER_144_1153 ();
 FILLCELL_X1 FILLER_144_1183 ();
 FILLCELL_X1 FILLER_144_1194 ();
 FILLCELL_X1 FILLER_144_1205 ();
 FILLCELL_X4 FILLER_144_1212 ();
 FILLCELL_X1 FILLER_144_1216 ();
 FILLCELL_X4 FILLER_144_1277 ();
 FILLCELL_X2 FILLER_144_1281 ();
 FILLCELL_X2 FILLER_144_1293 ();
 FILLCELL_X32 FILLER_144_1325 ();
 FILLCELL_X16 FILLER_144_1357 ();
 FILLCELL_X8 FILLER_144_1373 ();
 FILLCELL_X4 FILLER_144_1381 ();
 FILLCELL_X2 FILLER_144_1385 ();
 FILLCELL_X8 FILLER_144_1401 ();
 FILLCELL_X2 FILLER_144_1414 ();
 FILLCELL_X8 FILLER_144_1436 ();
 FILLCELL_X1 FILLER_144_1444 ();
 FILLCELL_X2 FILLER_144_1454 ();
 FILLCELL_X1 FILLER_144_1456 ();
 FILLCELL_X1 FILLER_144_1477 ();
 FILLCELL_X2 FILLER_144_1504 ();
 FILLCELL_X4 FILLER_144_1531 ();
 FILLCELL_X2 FILLER_144_1535 ();
 FILLCELL_X32 FILLER_144_1586 ();
 FILLCELL_X32 FILLER_144_1618 ();
 FILLCELL_X1 FILLER_144_1650 ();
 FILLCELL_X4 FILLER_145_1 ();
 FILLCELL_X2 FILLER_145_5 ();
 FILLCELL_X1 FILLER_145_27 ();
 FILLCELL_X2 FILLER_145_35 ();
 FILLCELL_X1 FILLER_145_37 ();
 FILLCELL_X1 FILLER_145_64 ();
 FILLCELL_X4 FILLER_145_72 ();
 FILLCELL_X2 FILLER_145_76 ();
 FILLCELL_X16 FILLER_145_85 ();
 FILLCELL_X2 FILLER_145_101 ();
 FILLCELL_X2 FILLER_145_112 ();
 FILLCELL_X2 FILLER_145_141 ();
 FILLCELL_X4 FILLER_145_152 ();
 FILLCELL_X4 FILLER_145_176 ();
 FILLCELL_X1 FILLER_145_180 ();
 FILLCELL_X2 FILLER_145_188 ();
 FILLCELL_X2 FILLER_145_203 ();
 FILLCELL_X1 FILLER_145_205 ();
 FILLCELL_X4 FILLER_145_228 ();
 FILLCELL_X2 FILLER_145_232 ();
 FILLCELL_X1 FILLER_145_234 ();
 FILLCELL_X4 FILLER_145_238 ();
 FILLCELL_X2 FILLER_145_242 ();
 FILLCELL_X4 FILLER_145_258 ();
 FILLCELL_X2 FILLER_145_262 ();
 FILLCELL_X1 FILLER_145_272 ();
 FILLCELL_X4 FILLER_145_276 ();
 FILLCELL_X4 FILLER_145_284 ();
 FILLCELL_X2 FILLER_145_291 ();
 FILLCELL_X1 FILLER_145_293 ();
 FILLCELL_X2 FILLER_145_303 ();
 FILLCELL_X1 FILLER_145_309 ();
 FILLCELL_X8 FILLER_145_327 ();
 FILLCELL_X2 FILLER_145_339 ();
 FILLCELL_X2 FILLER_145_344 ();
 FILLCELL_X1 FILLER_145_346 ();
 FILLCELL_X1 FILLER_145_352 ();
 FILLCELL_X2 FILLER_145_357 ();
 FILLCELL_X8 FILLER_145_363 ();
 FILLCELL_X2 FILLER_145_371 ();
 FILLCELL_X1 FILLER_145_373 ();
 FILLCELL_X2 FILLER_145_381 ();
 FILLCELL_X4 FILLER_145_386 ();
 FILLCELL_X1 FILLER_145_410 ();
 FILLCELL_X8 FILLER_145_414 ();
 FILLCELL_X4 FILLER_145_422 ();
 FILLCELL_X1 FILLER_145_426 ();
 FILLCELL_X2 FILLER_145_459 ();
 FILLCELL_X1 FILLER_145_461 ();
 FILLCELL_X1 FILLER_145_483 ();
 FILLCELL_X2 FILLER_145_498 ();
 FILLCELL_X4 FILLER_145_522 ();
 FILLCELL_X2 FILLER_145_526 ();
 FILLCELL_X1 FILLER_145_528 ();
 FILLCELL_X2 FILLER_145_532 ();
 FILLCELL_X8 FILLER_145_538 ();
 FILLCELL_X2 FILLER_145_546 ();
 FILLCELL_X1 FILLER_145_548 ();
 FILLCELL_X4 FILLER_145_582 ();
 FILLCELL_X2 FILLER_145_595 ();
 FILLCELL_X1 FILLER_145_597 ();
 FILLCELL_X4 FILLER_145_609 ();
 FILLCELL_X2 FILLER_145_613 ();
 FILLCELL_X1 FILLER_145_643 ();
 FILLCELL_X4 FILLER_145_664 ();
 FILLCELL_X1 FILLER_145_668 ();
 FILLCELL_X2 FILLER_145_672 ();
 FILLCELL_X8 FILLER_145_723 ();
 FILLCELL_X16 FILLER_145_749 ();
 FILLCELL_X8 FILLER_145_765 ();
 FILLCELL_X4 FILLER_145_773 ();
 FILLCELL_X16 FILLER_145_794 ();
 FILLCELL_X8 FILLER_145_810 ();
 FILLCELL_X4 FILLER_145_818 ();
 FILLCELL_X1 FILLER_145_822 ();
 FILLCELL_X16 FILLER_145_830 ();
 FILLCELL_X1 FILLER_145_846 ();
 FILLCELL_X16 FILLER_145_869 ();
 FILLCELL_X32 FILLER_145_890 ();
 FILLCELL_X2 FILLER_145_922 ();
 FILLCELL_X4 FILLER_145_929 ();
 FILLCELL_X4 FILLER_145_953 ();
 FILLCELL_X4 FILLER_145_973 ();
 FILLCELL_X2 FILLER_145_977 ();
 FILLCELL_X8 FILLER_145_1015 ();
 FILLCELL_X1 FILLER_145_1023 ();
 FILLCELL_X1 FILLER_145_1046 ();
 FILLCELL_X16 FILLER_145_1067 ();
 FILLCELL_X8 FILLER_145_1083 ();
 FILLCELL_X2 FILLER_145_1091 ();
 FILLCELL_X1 FILLER_145_1138 ();
 FILLCELL_X2 FILLER_145_1151 ();
 FILLCELL_X8 FILLER_145_1159 ();
 FILLCELL_X1 FILLER_145_1167 ();
 FILLCELL_X16 FILLER_145_1174 ();
 FILLCELL_X8 FILLER_145_1190 ();
 FILLCELL_X1 FILLER_145_1198 ();
 FILLCELL_X4 FILLER_145_1219 ();
 FILLCELL_X1 FILLER_145_1223 ();
 FILLCELL_X2 FILLER_145_1230 ();
 FILLCELL_X8 FILLER_145_1242 ();
 FILLCELL_X1 FILLER_145_1250 ();
 FILLCELL_X4 FILLER_145_1257 ();
 FILLCELL_X2 FILLER_145_1261 ();
 FILLCELL_X8 FILLER_145_1264 ();
 FILLCELL_X4 FILLER_145_1272 ();
 FILLCELL_X2 FILLER_145_1276 ();
 FILLCELL_X1 FILLER_145_1278 ();
 FILLCELL_X8 FILLER_145_1288 ();
 FILLCELL_X1 FILLER_145_1308 ();
 FILLCELL_X32 FILLER_145_1313 ();
 FILLCELL_X32 FILLER_145_1345 ();
 FILLCELL_X16 FILLER_145_1377 ();
 FILLCELL_X8 FILLER_145_1393 ();
 FILLCELL_X4 FILLER_145_1423 ();
 FILLCELL_X2 FILLER_145_1427 ();
 FILLCELL_X1 FILLER_145_1429 ();
 FILLCELL_X1 FILLER_145_1433 ();
 FILLCELL_X8 FILLER_145_1439 ();
 FILLCELL_X1 FILLER_145_1447 ();
 FILLCELL_X16 FILLER_145_1457 ();
 FILLCELL_X1 FILLER_145_1473 ();
 FILLCELL_X2 FILLER_145_1493 ();
 FILLCELL_X1 FILLER_145_1495 ();
 FILLCELL_X8 FILLER_145_1509 ();
 FILLCELL_X4 FILLER_145_1517 ();
 FILLCELL_X2 FILLER_145_1521 ();
 FILLCELL_X4 FILLER_145_1527 ();
 FILLCELL_X2 FILLER_145_1531 ();
 FILLCELL_X4 FILLER_145_1536 ();
 FILLCELL_X2 FILLER_145_1540 ();
 FILLCELL_X2 FILLER_145_1551 ();
 FILLCELL_X1 FILLER_145_1562 ();
 FILLCELL_X32 FILLER_145_1568 ();
 FILLCELL_X32 FILLER_145_1600 ();
 FILLCELL_X16 FILLER_145_1632 ();
 FILLCELL_X2 FILLER_145_1648 ();
 FILLCELL_X1 FILLER_145_1650 ();
 FILLCELL_X8 FILLER_146_1 ();
 FILLCELL_X4 FILLER_146_9 ();
 FILLCELL_X4 FILLER_146_40 ();
 FILLCELL_X2 FILLER_146_44 ();
 FILLCELL_X1 FILLER_146_46 ();
 FILLCELL_X1 FILLER_146_67 ();
 FILLCELL_X1 FILLER_146_88 ();
 FILLCELL_X4 FILLER_146_98 ();
 FILLCELL_X1 FILLER_146_115 ();
 FILLCELL_X1 FILLER_146_123 ();
 FILLCELL_X8 FILLER_146_144 ();
 FILLCELL_X2 FILLER_146_152 ();
 FILLCELL_X1 FILLER_146_154 ();
 FILLCELL_X4 FILLER_146_162 ();
 FILLCELL_X1 FILLER_146_186 ();
 FILLCELL_X4 FILLER_146_239 ();
 FILLCELL_X2 FILLER_146_243 ();
 FILLCELL_X2 FILLER_146_268 ();
 FILLCELL_X1 FILLER_146_270 ();
 FILLCELL_X4 FILLER_146_303 ();
 FILLCELL_X2 FILLER_146_312 ();
 FILLCELL_X4 FILLER_146_325 ();
 FILLCELL_X8 FILLER_146_333 ();
 FILLCELL_X2 FILLER_146_341 ();
 FILLCELL_X1 FILLER_146_343 ();
 FILLCELL_X1 FILLER_146_356 ();
 FILLCELL_X8 FILLER_146_377 ();
 FILLCELL_X2 FILLER_146_385 ();
 FILLCELL_X1 FILLER_146_387 ();
 FILLCELL_X2 FILLER_146_392 ();
 FILLCELL_X1 FILLER_146_401 ();
 FILLCELL_X8 FILLER_146_436 ();
 FILLCELL_X2 FILLER_146_444 ();
 FILLCELL_X1 FILLER_146_446 ();
 FILLCELL_X2 FILLER_146_468 ();
 FILLCELL_X1 FILLER_146_470 ();
 FILLCELL_X8 FILLER_146_478 ();
 FILLCELL_X1 FILLER_146_486 ();
 FILLCELL_X2 FILLER_146_494 ();
 FILLCELL_X16 FILLER_146_516 ();
 FILLCELL_X2 FILLER_146_532 ();
 FILLCELL_X16 FILLER_146_537 ();
 FILLCELL_X2 FILLER_146_553 ();
 FILLCELL_X1 FILLER_146_555 ();
 FILLCELL_X1 FILLER_146_569 ();
 FILLCELL_X8 FILLER_146_621 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X2 FILLER_146_632 ();
 FILLCELL_X4 FILLER_146_639 ();
 FILLCELL_X1 FILLER_146_643 ();
 FILLCELL_X4 FILLER_146_648 ();
 FILLCELL_X2 FILLER_146_652 ();
 FILLCELL_X1 FILLER_146_654 ();
 FILLCELL_X1 FILLER_146_658 ();
 FILLCELL_X2 FILLER_146_724 ();
 FILLCELL_X1 FILLER_146_730 ();
 FILLCELL_X1 FILLER_146_734 ();
 FILLCELL_X1 FILLER_146_755 ();
 FILLCELL_X1 FILLER_146_776 ();
 FILLCELL_X1 FILLER_146_784 ();
 FILLCELL_X4 FILLER_146_805 ();
 FILLCELL_X2 FILLER_146_809 ();
 FILLCELL_X1 FILLER_146_833 ();
 FILLCELL_X2 FILLER_146_886 ();
 FILLCELL_X1 FILLER_146_888 ();
 FILLCELL_X1 FILLER_146_934 ();
 FILLCELL_X4 FILLER_146_942 ();
 FILLCELL_X2 FILLER_146_1009 ();
 FILLCELL_X1 FILLER_146_1031 ();
 FILLCELL_X2 FILLER_146_1044 ();
 FILLCELL_X1 FILLER_146_1046 ();
 FILLCELL_X8 FILLER_146_1052 ();
 FILLCELL_X2 FILLER_146_1060 ();
 FILLCELL_X1 FILLER_146_1062 ();
 FILLCELL_X4 FILLER_146_1090 ();
 FILLCELL_X2 FILLER_146_1094 ();
 FILLCELL_X1 FILLER_146_1118 ();
 FILLCELL_X4 FILLER_146_1128 ();
 FILLCELL_X2 FILLER_146_1144 ();
 FILLCELL_X1 FILLER_146_1146 ();
 FILLCELL_X16 FILLER_146_1163 ();
 FILLCELL_X4 FILLER_146_1179 ();
 FILLCELL_X2 FILLER_146_1183 ();
 FILLCELL_X1 FILLER_146_1185 ();
 FILLCELL_X8 FILLER_146_1207 ();
 FILLCELL_X1 FILLER_146_1215 ();
 FILLCELL_X2 FILLER_146_1225 ();
 FILLCELL_X2 FILLER_146_1232 ();
 FILLCELL_X1 FILLER_146_1234 ();
 FILLCELL_X2 FILLER_146_1248 ();
 FILLCELL_X1 FILLER_146_1250 ();
 FILLCELL_X1 FILLER_146_1255 ();
 FILLCELL_X8 FILLER_146_1260 ();
 FILLCELL_X2 FILLER_146_1268 ();
 FILLCELL_X4 FILLER_146_1289 ();
 FILLCELL_X32 FILLER_146_1319 ();
 FILLCELL_X32 FILLER_146_1351 ();
 FILLCELL_X4 FILLER_146_1383 ();
 FILLCELL_X2 FILLER_146_1387 ();
 FILLCELL_X1 FILLER_146_1389 ();
 FILLCELL_X1 FILLER_146_1400 ();
 FILLCELL_X4 FILLER_146_1410 ();
 FILLCELL_X2 FILLER_146_1423 ();
 FILLCELL_X2 FILLER_146_1436 ();
 FILLCELL_X1 FILLER_146_1438 ();
 FILLCELL_X4 FILLER_146_1443 ();
 FILLCELL_X1 FILLER_146_1447 ();
 FILLCELL_X2 FILLER_146_1452 ();
 FILLCELL_X16 FILLER_146_1457 ();
 FILLCELL_X8 FILLER_146_1500 ();
 FILLCELL_X1 FILLER_146_1508 ();
 FILLCELL_X8 FILLER_146_1530 ();
 FILLCELL_X4 FILLER_146_1538 ();
 FILLCELL_X2 FILLER_146_1542 ();
 FILLCELL_X1 FILLER_146_1544 ();
 FILLCELL_X4 FILLER_146_1548 ();
 FILLCELL_X1 FILLER_146_1552 ();
 FILLCELL_X32 FILLER_146_1557 ();
 FILLCELL_X32 FILLER_146_1589 ();
 FILLCELL_X16 FILLER_146_1621 ();
 FILLCELL_X8 FILLER_146_1637 ();
 FILLCELL_X4 FILLER_146_1645 ();
 FILLCELL_X2 FILLER_146_1649 ();
 FILLCELL_X16 FILLER_147_1 ();
 FILLCELL_X2 FILLER_147_17 ();
 FILLCELL_X1 FILLER_147_19 ();
 FILLCELL_X8 FILLER_147_49 ();
 FILLCELL_X4 FILLER_147_57 ();
 FILLCELL_X2 FILLER_147_61 ();
 FILLCELL_X1 FILLER_147_63 ();
 FILLCELL_X1 FILLER_147_73 ();
 FILLCELL_X1 FILLER_147_81 ();
 FILLCELL_X2 FILLER_147_89 ();
 FILLCELL_X1 FILLER_147_111 ();
 FILLCELL_X8 FILLER_147_119 ();
 FILLCELL_X2 FILLER_147_127 ();
 FILLCELL_X1 FILLER_147_129 ();
 FILLCELL_X4 FILLER_147_172 ();
 FILLCELL_X2 FILLER_147_176 ();
 FILLCELL_X1 FILLER_147_178 ();
 FILLCELL_X4 FILLER_147_202 ();
 FILLCELL_X1 FILLER_147_206 ();
 FILLCELL_X4 FILLER_147_211 ();
 FILLCELL_X1 FILLER_147_215 ();
 FILLCELL_X1 FILLER_147_248 ();
 FILLCELL_X4 FILLER_147_276 ();
 FILLCELL_X2 FILLER_147_280 ();
 FILLCELL_X16 FILLER_147_286 ();
 FILLCELL_X1 FILLER_147_302 ();
 FILLCELL_X2 FILLER_147_353 ();
 FILLCELL_X8 FILLER_147_363 ();
 FILLCELL_X1 FILLER_147_371 ();
 FILLCELL_X2 FILLER_147_404 ();
 FILLCELL_X2 FILLER_147_413 ();
 FILLCELL_X1 FILLER_147_418 ();
 FILLCELL_X8 FILLER_147_446 ();
 FILLCELL_X2 FILLER_147_454 ();
 FILLCELL_X1 FILLER_147_456 ();
 FILLCELL_X1 FILLER_147_471 ();
 FILLCELL_X8 FILLER_147_479 ();
 FILLCELL_X1 FILLER_147_487 ();
 FILLCELL_X1 FILLER_147_493 ();
 FILLCELL_X16 FILLER_147_501 ();
 FILLCELL_X2 FILLER_147_554 ();
 FILLCELL_X8 FILLER_147_574 ();
 FILLCELL_X4 FILLER_147_582 ();
 FILLCELL_X8 FILLER_147_610 ();
 FILLCELL_X2 FILLER_147_618 ();
 FILLCELL_X2 FILLER_147_623 ();
 FILLCELL_X1 FILLER_147_625 ();
 FILLCELL_X8 FILLER_147_630 ();
 FILLCELL_X2 FILLER_147_638 ();
 FILLCELL_X1 FILLER_147_665 ();
 FILLCELL_X4 FILLER_147_745 ();
 FILLCELL_X2 FILLER_147_802 ();
 FILLCELL_X4 FILLER_147_854 ();
 FILLCELL_X2 FILLER_147_858 ();
 FILLCELL_X2 FILLER_147_919 ();
 FILLCELL_X1 FILLER_147_927 ();
 FILLCELL_X8 FILLER_147_935 ();
 FILLCELL_X1 FILLER_147_943 ();
 FILLCELL_X2 FILLER_147_951 ();
 FILLCELL_X8 FILLER_147_976 ();
 FILLCELL_X4 FILLER_147_984 ();
 FILLCELL_X2 FILLER_147_988 ();
 FILLCELL_X1 FILLER_147_990 ();
 FILLCELL_X4 FILLER_147_1000 ();
 FILLCELL_X4 FILLER_147_1036 ();
 FILLCELL_X16 FILLER_147_1060 ();
 FILLCELL_X8 FILLER_147_1076 ();
 FILLCELL_X1 FILLER_147_1084 ();
 FILLCELL_X16 FILLER_147_1092 ();
 FILLCELL_X2 FILLER_147_1108 ();
 FILLCELL_X1 FILLER_147_1110 ();
 FILLCELL_X16 FILLER_147_1116 ();
 FILLCELL_X8 FILLER_147_1132 ();
 FILLCELL_X4 FILLER_147_1140 ();
 FILLCELL_X1 FILLER_147_1144 ();
 FILLCELL_X16 FILLER_147_1167 ();
 FILLCELL_X8 FILLER_147_1183 ();
 FILLCELL_X4 FILLER_147_1191 ();
 FILLCELL_X2 FILLER_147_1195 ();
 FILLCELL_X2 FILLER_147_1200 ();
 FILLCELL_X4 FILLER_147_1221 ();
 FILLCELL_X1 FILLER_147_1225 ();
 FILLCELL_X2 FILLER_147_1255 ();
 FILLCELL_X1 FILLER_147_1257 ();
 FILLCELL_X32 FILLER_147_1308 ();
 FILLCELL_X32 FILLER_147_1340 ();
 FILLCELL_X16 FILLER_147_1372 ();
 FILLCELL_X2 FILLER_147_1388 ();
 FILLCELL_X1 FILLER_147_1398 ();
 FILLCELL_X1 FILLER_147_1402 ();
 FILLCELL_X8 FILLER_147_1410 ();
 FILLCELL_X1 FILLER_147_1418 ();
 FILLCELL_X2 FILLER_147_1434 ();
 FILLCELL_X2 FILLER_147_1443 ();
 FILLCELL_X16 FILLER_147_1455 ();
 FILLCELL_X4 FILLER_147_1484 ();
 FILLCELL_X2 FILLER_147_1492 ();
 FILLCELL_X2 FILLER_147_1499 ();
 FILLCELL_X1 FILLER_147_1501 ();
 FILLCELL_X8 FILLER_147_1506 ();
 FILLCELL_X1 FILLER_147_1514 ();
 FILLCELL_X2 FILLER_147_1524 ();
 FILLCELL_X2 FILLER_147_1535 ();
 FILLCELL_X4 FILLER_147_1541 ();
 FILLCELL_X4 FILLER_147_1562 ();
 FILLCELL_X2 FILLER_147_1566 ();
 FILLCELL_X1 FILLER_147_1568 ();
 FILLCELL_X32 FILLER_147_1576 ();
 FILLCELL_X32 FILLER_147_1608 ();
 FILLCELL_X8 FILLER_147_1640 ();
 FILLCELL_X2 FILLER_147_1648 ();
 FILLCELL_X1 FILLER_147_1650 ();
 FILLCELL_X16 FILLER_148_1 ();
 FILLCELL_X4 FILLER_148_17 ();
 FILLCELL_X2 FILLER_148_21 ();
 FILLCELL_X2 FILLER_148_43 ();
 FILLCELL_X4 FILLER_148_72 ();
 FILLCELL_X1 FILLER_148_76 ();
 FILLCELL_X32 FILLER_148_102 ();
 FILLCELL_X8 FILLER_148_134 ();
 FILLCELL_X4 FILLER_148_142 ();
 FILLCELL_X2 FILLER_148_146 ();
 FILLCELL_X1 FILLER_148_148 ();
 FILLCELL_X2 FILLER_148_154 ();
 FILLCELL_X2 FILLER_148_163 ();
 FILLCELL_X1 FILLER_148_165 ();
 FILLCELL_X1 FILLER_148_193 ();
 FILLCELL_X1 FILLER_148_199 ();
 FILLCELL_X2 FILLER_148_207 ();
 FILLCELL_X2 FILLER_148_229 ();
 FILLCELL_X2 FILLER_148_244 ();
 FILLCELL_X2 FILLER_148_253 ();
 FILLCELL_X1 FILLER_148_275 ();
 FILLCELL_X1 FILLER_148_279 ();
 FILLCELL_X4 FILLER_148_300 ();
 FILLCELL_X1 FILLER_148_308 ();
 FILLCELL_X1 FILLER_148_313 ();
 FILLCELL_X1 FILLER_148_317 ();
 FILLCELL_X1 FILLER_148_327 ();
 FILLCELL_X2 FILLER_148_348 ();
 FILLCELL_X8 FILLER_148_409 ();
 FILLCELL_X2 FILLER_148_417 ();
 FILLCELL_X1 FILLER_148_419 ();
 FILLCELL_X8 FILLER_148_434 ();
 FILLCELL_X4 FILLER_148_442 ();
 FILLCELL_X1 FILLER_148_446 ();
 FILLCELL_X4 FILLER_148_454 ();
 FILLCELL_X2 FILLER_148_472 ();
 FILLCELL_X2 FILLER_148_488 ();
 FILLCELL_X2 FILLER_148_497 ();
 FILLCELL_X1 FILLER_148_499 ();
 FILLCELL_X1 FILLER_148_504 ();
 FILLCELL_X2 FILLER_148_510 ();
 FILLCELL_X1 FILLER_148_512 ();
 FILLCELL_X4 FILLER_148_517 ();
 FILLCELL_X1 FILLER_148_528 ();
 FILLCELL_X8 FILLER_148_566 ();
 FILLCELL_X1 FILLER_148_578 ();
 FILLCELL_X1 FILLER_148_586 ();
 FILLCELL_X1 FILLER_148_590 ();
 FILLCELL_X2 FILLER_148_596 ();
 FILLCELL_X1 FILLER_148_618 ();
 FILLCELL_X2 FILLER_148_675 ();
 FILLCELL_X1 FILLER_148_680 ();
 FILLCELL_X1 FILLER_148_710 ();
 FILLCELL_X4 FILLER_148_721 ();
 FILLCELL_X1 FILLER_148_725 ();
 FILLCELL_X4 FILLER_148_737 ();
 FILLCELL_X2 FILLER_148_768 ();
 FILLCELL_X1 FILLER_148_770 ();
 FILLCELL_X4 FILLER_148_792 ();
 FILLCELL_X1 FILLER_148_796 ();
 FILLCELL_X2 FILLER_148_825 ();
 FILLCELL_X8 FILLER_148_859 ();
 FILLCELL_X2 FILLER_148_867 ();
 FILLCELL_X4 FILLER_148_876 ();
 FILLCELL_X2 FILLER_148_880 ();
 FILLCELL_X2 FILLER_148_905 ();
 FILLCELL_X1 FILLER_148_907 ();
 FILLCELL_X4 FILLER_148_915 ();
 FILLCELL_X1 FILLER_148_924 ();
 FILLCELL_X1 FILLER_148_950 ();
 FILLCELL_X8 FILLER_148_983 ();
 FILLCELL_X4 FILLER_148_991 ();
 FILLCELL_X1 FILLER_148_1031 ();
 FILLCELL_X2 FILLER_148_1081 ();
 FILLCELL_X1 FILLER_148_1083 ();
 FILLCELL_X32 FILLER_148_1111 ();
 FILLCELL_X32 FILLER_148_1143 ();
 FILLCELL_X16 FILLER_148_1175 ();
 FILLCELL_X2 FILLER_148_1191 ();
 FILLCELL_X1 FILLER_148_1193 ();
 FILLCELL_X16 FILLER_148_1210 ();
 FILLCELL_X2 FILLER_148_1226 ();
 FILLCELL_X1 FILLER_148_1228 ();
 FILLCELL_X4 FILLER_148_1234 ();
 FILLCELL_X1 FILLER_148_1238 ();
 FILLCELL_X1 FILLER_148_1247 ();
 FILLCELL_X32 FILLER_148_1293 ();
 FILLCELL_X32 FILLER_148_1325 ();
 FILLCELL_X16 FILLER_148_1357 ();
 FILLCELL_X8 FILLER_148_1373 ();
 FILLCELL_X4 FILLER_148_1381 ();
 FILLCELL_X2 FILLER_148_1385 ();
 FILLCELL_X1 FILLER_148_1387 ();
 FILLCELL_X1 FILLER_148_1402 ();
 FILLCELL_X1 FILLER_148_1419 ();
 FILLCELL_X2 FILLER_148_1440 ();
 FILLCELL_X1 FILLER_148_1442 ();
 FILLCELL_X8 FILLER_148_1461 ();
 FILLCELL_X2 FILLER_148_1469 ();
 FILLCELL_X8 FILLER_148_1483 ();
 FILLCELL_X4 FILLER_148_1493 ();
 FILLCELL_X2 FILLER_148_1497 ();
 FILLCELL_X8 FILLER_148_1509 ();
 FILLCELL_X2 FILLER_148_1517 ();
 FILLCELL_X1 FILLER_148_1526 ();
 FILLCELL_X1 FILLER_148_1533 ();
 FILLCELL_X4 FILLER_148_1543 ();
 FILLCELL_X8 FILLER_148_1550 ();
 FILLCELL_X32 FILLER_148_1572 ();
 FILLCELL_X32 FILLER_148_1604 ();
 FILLCELL_X8 FILLER_148_1636 ();
 FILLCELL_X4 FILLER_148_1644 ();
 FILLCELL_X2 FILLER_148_1648 ();
 FILLCELL_X1 FILLER_148_1650 ();
 FILLCELL_X16 FILLER_149_1 ();
 FILLCELL_X2 FILLER_149_17 ();
 FILLCELL_X1 FILLER_149_19 ();
 FILLCELL_X8 FILLER_149_28 ();
 FILLCELL_X2 FILLER_149_36 ();
 FILLCELL_X4 FILLER_149_45 ();
 FILLCELL_X32 FILLER_149_56 ();
 FILLCELL_X8 FILLER_149_88 ();
 FILLCELL_X4 FILLER_149_96 ();
 FILLCELL_X2 FILLER_149_100 ();
 FILLCELL_X2 FILLER_149_122 ();
 FILLCELL_X1 FILLER_149_124 ();
 FILLCELL_X1 FILLER_149_154 ();
 FILLCELL_X16 FILLER_149_168 ();
 FILLCELL_X1 FILLER_149_184 ();
 FILLCELL_X2 FILLER_149_205 ();
 FILLCELL_X4 FILLER_149_221 ();
 FILLCELL_X2 FILLER_149_225 ();
 FILLCELL_X1 FILLER_149_227 ();
 FILLCELL_X4 FILLER_149_260 ();
 FILLCELL_X4 FILLER_149_268 ();
 FILLCELL_X2 FILLER_149_272 ();
 FILLCELL_X4 FILLER_149_277 ();
 FILLCELL_X8 FILLER_149_323 ();
 FILLCELL_X2 FILLER_149_331 ();
 FILLCELL_X1 FILLER_149_333 ();
 FILLCELL_X1 FILLER_149_338 ();
 FILLCELL_X16 FILLER_149_342 ();
 FILLCELL_X1 FILLER_149_358 ();
 FILLCELL_X4 FILLER_149_363 ();
 FILLCELL_X2 FILLER_149_367 ();
 FILLCELL_X8 FILLER_149_372 ();
 FILLCELL_X4 FILLER_149_380 ();
 FILLCELL_X2 FILLER_149_384 ();
 FILLCELL_X1 FILLER_149_386 ();
 FILLCELL_X4 FILLER_149_391 ();
 FILLCELL_X1 FILLER_149_395 ();
 FILLCELL_X4 FILLER_149_404 ();
 FILLCELL_X1 FILLER_149_408 ();
 FILLCELL_X8 FILLER_149_413 ();
 FILLCELL_X2 FILLER_149_421 ();
 FILLCELL_X2 FILLER_149_444 ();
 FILLCELL_X2 FILLER_149_449 ();
 FILLCELL_X1 FILLER_149_451 ();
 FILLCELL_X4 FILLER_149_459 ();
 FILLCELL_X1 FILLER_149_463 ();
 FILLCELL_X1 FILLER_149_471 ();
 FILLCELL_X4 FILLER_149_489 ();
 FILLCELL_X1 FILLER_149_513 ();
 FILLCELL_X2 FILLER_149_536 ();
 FILLCELL_X2 FILLER_149_541 ();
 FILLCELL_X1 FILLER_149_543 ();
 FILLCELL_X8 FILLER_149_548 ();
 FILLCELL_X4 FILLER_149_556 ();
 FILLCELL_X2 FILLER_149_589 ();
 FILLCELL_X1 FILLER_149_591 ();
 FILLCELL_X2 FILLER_149_595 ();
 FILLCELL_X1 FILLER_149_648 ();
 FILLCELL_X2 FILLER_149_652 ();
 FILLCELL_X1 FILLER_149_654 ();
 FILLCELL_X4 FILLER_149_659 ();
 FILLCELL_X1 FILLER_149_753 ();
 FILLCELL_X2 FILLER_149_794 ();
 FILLCELL_X1 FILLER_149_796 ();
 FILLCELL_X2 FILLER_149_827 ();
 FILLCELL_X4 FILLER_149_836 ();
 FILLCELL_X4 FILLER_149_847 ();
 FILLCELL_X1 FILLER_149_851 ();
 FILLCELL_X4 FILLER_149_879 ();
 FILLCELL_X1 FILLER_149_890 ();
 FILLCELL_X4 FILLER_149_945 ();
 FILLCELL_X2 FILLER_149_949 ();
 FILLCELL_X1 FILLER_149_991 ();
 FILLCELL_X8 FILLER_149_1027 ();
 FILLCELL_X2 FILLER_149_1035 ();
 FILLCELL_X2 FILLER_149_1057 ();
 FILLCELL_X1 FILLER_149_1059 ();
 FILLCELL_X32 FILLER_149_1093 ();
 FILLCELL_X32 FILLER_149_1125 ();
 FILLCELL_X32 FILLER_149_1157 ();
 FILLCELL_X32 FILLER_149_1189 ();
 FILLCELL_X8 FILLER_149_1221 ();
 FILLCELL_X2 FILLER_149_1241 ();
 FILLCELL_X1 FILLER_149_1243 ();
 FILLCELL_X8 FILLER_149_1254 ();
 FILLCELL_X1 FILLER_149_1262 ();
 FILLCELL_X1 FILLER_149_1275 ();
 FILLCELL_X32 FILLER_149_1279 ();
 FILLCELL_X32 FILLER_149_1311 ();
 FILLCELL_X32 FILLER_149_1343 ();
 FILLCELL_X16 FILLER_149_1375 ();
 FILLCELL_X4 FILLER_149_1391 ();
 FILLCELL_X2 FILLER_149_1438 ();
 FILLCELL_X1 FILLER_149_1440 ();
 FILLCELL_X2 FILLER_149_1445 ();
 FILLCELL_X1 FILLER_149_1447 ();
 FILLCELL_X16 FILLER_149_1455 ();
 FILLCELL_X8 FILLER_149_1482 ();
 FILLCELL_X1 FILLER_149_1490 ();
 FILLCELL_X8 FILLER_149_1496 ();
 FILLCELL_X4 FILLER_149_1513 ();
 FILLCELL_X1 FILLER_149_1517 ();
 FILLCELL_X4 FILLER_149_1522 ();
 FILLCELL_X1 FILLER_149_1529 ();
 FILLCELL_X1 FILLER_149_1534 ();
 FILLCELL_X4 FILLER_149_1554 ();
 FILLCELL_X1 FILLER_149_1558 ();
 FILLCELL_X32 FILLER_149_1569 ();
 FILLCELL_X32 FILLER_149_1601 ();
 FILLCELL_X16 FILLER_149_1633 ();
 FILLCELL_X2 FILLER_149_1649 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X16 FILLER_150_33 ();
 FILLCELL_X1 FILLER_150_49 ();
 FILLCELL_X8 FILLER_150_106 ();
 FILLCELL_X2 FILLER_150_114 ();
 FILLCELL_X1 FILLER_150_123 ();
 FILLCELL_X4 FILLER_150_135 ();
 FILLCELL_X1 FILLER_150_139 ();
 FILLCELL_X4 FILLER_150_149 ();
 FILLCELL_X8 FILLER_150_180 ();
 FILLCELL_X2 FILLER_150_192 ();
 FILLCELL_X1 FILLER_150_194 ();
 FILLCELL_X4 FILLER_150_199 ();
 FILLCELL_X2 FILLER_150_203 ();
 FILLCELL_X1 FILLER_150_205 ();
 FILLCELL_X8 FILLER_150_231 ();
 FILLCELL_X4 FILLER_150_239 ();
 FILLCELL_X1 FILLER_150_243 ();
 FILLCELL_X4 FILLER_150_271 ();
 FILLCELL_X2 FILLER_150_275 ();
 FILLCELL_X4 FILLER_150_301 ();
 FILLCELL_X2 FILLER_150_305 ();
 FILLCELL_X2 FILLER_150_311 ();
 FILLCELL_X1 FILLER_150_313 ();
 FILLCELL_X2 FILLER_150_338 ();
 FILLCELL_X1 FILLER_150_340 ();
 FILLCELL_X8 FILLER_150_344 ();
 FILLCELL_X2 FILLER_150_376 ();
 FILLCELL_X1 FILLER_150_378 ();
 FILLCELL_X1 FILLER_150_402 ();
 FILLCELL_X4 FILLER_150_457 ();
 FILLCELL_X2 FILLER_150_461 ();
 FILLCELL_X4 FILLER_150_487 ();
 FILLCELL_X2 FILLER_150_491 ();
 FILLCELL_X1 FILLER_150_493 ();
 FILLCELL_X8 FILLER_150_501 ();
 FILLCELL_X1 FILLER_150_509 ();
 FILLCELL_X4 FILLER_150_513 ();
 FILLCELL_X2 FILLER_150_564 ();
 FILLCELL_X1 FILLER_150_566 ();
 FILLCELL_X8 FILLER_150_597 ();
 FILLCELL_X4 FILLER_150_605 ();
 FILLCELL_X8 FILLER_150_616 ();
 FILLCELL_X4 FILLER_150_624 ();
 FILLCELL_X2 FILLER_150_628 ();
 FILLCELL_X1 FILLER_150_630 ();
 FILLCELL_X8 FILLER_150_641 ();
 FILLCELL_X2 FILLER_150_649 ();
 FILLCELL_X8 FILLER_150_658 ();
 FILLCELL_X2 FILLER_150_670 ();
 FILLCELL_X1 FILLER_150_672 ();
 FILLCELL_X1 FILLER_150_680 ();
 FILLCELL_X2 FILLER_150_684 ();
 FILLCELL_X2 FILLER_150_689 ();
 FILLCELL_X1 FILLER_150_691 ();
 FILLCELL_X4 FILLER_150_697 ();
 FILLCELL_X2 FILLER_150_701 ();
 FILLCELL_X8 FILLER_150_710 ();
 FILLCELL_X4 FILLER_150_718 ();
 FILLCELL_X2 FILLER_150_722 ();
 FILLCELL_X1 FILLER_150_724 ();
 FILLCELL_X8 FILLER_150_737 ();
 FILLCELL_X4 FILLER_150_745 ();
 FILLCELL_X2 FILLER_150_749 ();
 FILLCELL_X1 FILLER_150_751 ();
 FILLCELL_X4 FILLER_150_789 ();
 FILLCELL_X1 FILLER_150_793 ();
 FILLCELL_X1 FILLER_150_801 ();
 FILLCELL_X4 FILLER_150_826 ();
 FILLCELL_X2 FILLER_150_850 ();
 FILLCELL_X1 FILLER_150_852 ();
 FILLCELL_X1 FILLER_150_858 ();
 FILLCELL_X2 FILLER_150_864 ();
 FILLCELL_X2 FILLER_150_893 ();
 FILLCELL_X1 FILLER_150_895 ();
 FILLCELL_X8 FILLER_150_903 ();
 FILLCELL_X4 FILLER_150_911 ();
 FILLCELL_X2 FILLER_150_915 ();
 FILLCELL_X2 FILLER_150_922 ();
 FILLCELL_X1 FILLER_150_944 ();
 FILLCELL_X1 FILLER_150_952 ();
 FILLCELL_X1 FILLER_150_960 ();
 FILLCELL_X1 FILLER_150_970 ();
 FILLCELL_X1 FILLER_150_978 ();
 FILLCELL_X1 FILLER_150_1006 ();
 FILLCELL_X2 FILLER_150_1014 ();
 FILLCELL_X8 FILLER_150_1036 ();
 FILLCELL_X32 FILLER_150_1085 ();
 FILLCELL_X32 FILLER_150_1117 ();
 FILLCELL_X32 FILLER_150_1149 ();
 FILLCELL_X32 FILLER_150_1181 ();
 FILLCELL_X4 FILLER_150_1213 ();
 FILLCELL_X32 FILLER_150_1250 ();
 FILLCELL_X32 FILLER_150_1282 ();
 FILLCELL_X32 FILLER_150_1314 ();
 FILLCELL_X32 FILLER_150_1346 ();
 FILLCELL_X16 FILLER_150_1378 ();
 FILLCELL_X2 FILLER_150_1394 ();
 FILLCELL_X1 FILLER_150_1396 ();
 FILLCELL_X4 FILLER_150_1429 ();
 FILLCELL_X4 FILLER_150_1445 ();
 FILLCELL_X2 FILLER_150_1462 ();
 FILLCELL_X4 FILLER_150_1476 ();
 FILLCELL_X1 FILLER_150_1480 ();
 FILLCELL_X4 FILLER_150_1484 ();
 FILLCELL_X1 FILLER_150_1488 ();
 FILLCELL_X16 FILLER_150_1498 ();
 FILLCELL_X2 FILLER_150_1514 ();
 FILLCELL_X2 FILLER_150_1527 ();
 FILLCELL_X1 FILLER_150_1529 ();
 FILLCELL_X32 FILLER_150_1567 ();
 FILLCELL_X32 FILLER_150_1599 ();
 FILLCELL_X16 FILLER_150_1631 ();
 FILLCELL_X4 FILLER_150_1647 ();
 FILLCELL_X16 FILLER_151_1 ();
 FILLCELL_X8 FILLER_151_17 ();
 FILLCELL_X4 FILLER_151_25 ();
 FILLCELL_X1 FILLER_151_29 ();
 FILLCELL_X2 FILLER_151_77 ();
 FILLCELL_X1 FILLER_151_86 ();
 FILLCELL_X4 FILLER_151_96 ();
 FILLCELL_X1 FILLER_151_100 ();
 FILLCELL_X8 FILLER_151_110 ();
 FILLCELL_X2 FILLER_151_118 ();
 FILLCELL_X1 FILLER_151_120 ();
 FILLCELL_X1 FILLER_151_141 ();
 FILLCELL_X2 FILLER_151_162 ();
 FILLCELL_X1 FILLER_151_164 ();
 FILLCELL_X4 FILLER_151_175 ();
 FILLCELL_X1 FILLER_151_190 ();
 FILLCELL_X1 FILLER_151_193 ();
 FILLCELL_X2 FILLER_151_211 ();
 FILLCELL_X4 FILLER_151_216 ();
 FILLCELL_X1 FILLER_151_240 ();
 FILLCELL_X4 FILLER_151_247 ();
 FILLCELL_X1 FILLER_151_251 ();
 FILLCELL_X2 FILLER_151_300 ();
 FILLCELL_X1 FILLER_151_348 ();
 FILLCELL_X1 FILLER_151_378 ();
 FILLCELL_X8 FILLER_151_384 ();
 FILLCELL_X4 FILLER_151_392 ();
 FILLCELL_X2 FILLER_151_396 ();
 FILLCELL_X2 FILLER_151_402 ();
 FILLCELL_X8 FILLER_151_427 ();
 FILLCELL_X2 FILLER_151_435 ();
 FILLCELL_X2 FILLER_151_453 ();
 FILLCELL_X4 FILLER_151_462 ();
 FILLCELL_X1 FILLER_151_491 ();
 FILLCELL_X1 FILLER_151_519 ();
 FILLCELL_X1 FILLER_151_524 ();
 FILLCELL_X1 FILLER_151_528 ();
 FILLCELL_X4 FILLER_151_534 ();
 FILLCELL_X2 FILLER_151_538 ();
 FILLCELL_X1 FILLER_151_540 ();
 FILLCELL_X1 FILLER_151_545 ();
 FILLCELL_X1 FILLER_151_549 ();
 FILLCELL_X2 FILLER_151_591 ();
 FILLCELL_X4 FILLER_151_627 ();
 FILLCELL_X8 FILLER_151_638 ();
 FILLCELL_X1 FILLER_151_646 ();
 FILLCELL_X1 FILLER_151_654 ();
 FILLCELL_X8 FILLER_151_662 ();
 FILLCELL_X4 FILLER_151_670 ();
 FILLCELL_X1 FILLER_151_674 ();
 FILLCELL_X2 FILLER_151_715 ();
 FILLCELL_X8 FILLER_151_737 ();
 FILLCELL_X1 FILLER_151_745 ();
 FILLCELL_X1 FILLER_151_766 ();
 FILLCELL_X8 FILLER_151_794 ();
 FILLCELL_X8 FILLER_151_809 ();
 FILLCELL_X1 FILLER_151_817 ();
 FILLCELL_X1 FILLER_151_825 ();
 FILLCELL_X4 FILLER_151_863 ();
 FILLCELL_X2 FILLER_151_867 ();
 FILLCELL_X1 FILLER_151_869 ();
 FILLCELL_X2 FILLER_151_890 ();
 FILLCELL_X1 FILLER_151_896 ();
 FILLCELL_X16 FILLER_151_906 ();
 FILLCELL_X1 FILLER_151_922 ();
 FILLCELL_X4 FILLER_151_938 ();
 FILLCELL_X1 FILLER_151_942 ();
 FILLCELL_X32 FILLER_151_963 ();
 FILLCELL_X2 FILLER_151_995 ();
 FILLCELL_X1 FILLER_151_997 ();
 FILLCELL_X4 FILLER_151_1018 ();
 FILLCELL_X2 FILLER_151_1022 ();
 FILLCELL_X32 FILLER_151_1044 ();
 FILLCELL_X4 FILLER_151_1076 ();
 FILLCELL_X2 FILLER_151_1080 ();
 FILLCELL_X1 FILLER_151_1082 ();
 FILLCELL_X32 FILLER_151_1088 ();
 FILLCELL_X32 FILLER_151_1120 ();
 FILLCELL_X32 FILLER_151_1152 ();
 FILLCELL_X32 FILLER_151_1184 ();
 FILLCELL_X8 FILLER_151_1216 ();
 FILLCELL_X4 FILLER_151_1224 ();
 FILLCELL_X8 FILLER_151_1234 ();
 FILLCELL_X1 FILLER_151_1242 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X32 FILLER_151_1296 ();
 FILLCELL_X32 FILLER_151_1328 ();
 FILLCELL_X32 FILLER_151_1360 ();
 FILLCELL_X2 FILLER_151_1392 ();
 FILLCELL_X2 FILLER_151_1401 ();
 FILLCELL_X2 FILLER_151_1411 ();
 FILLCELL_X1 FILLER_151_1413 ();
 FILLCELL_X8 FILLER_151_1428 ();
 FILLCELL_X1 FILLER_151_1436 ();
 FILLCELL_X2 FILLER_151_1444 ();
 FILLCELL_X4 FILLER_151_1482 ();
 FILLCELL_X4 FILLER_151_1509 ();
 FILLCELL_X1 FILLER_151_1513 ();
 FILLCELL_X1 FILLER_151_1521 ();
 FILLCELL_X1 FILLER_151_1525 ();
 FILLCELL_X2 FILLER_151_1530 ();
 FILLCELL_X4 FILLER_151_1536 ();
 FILLCELL_X2 FILLER_151_1540 ();
 FILLCELL_X2 FILLER_151_1561 ();
 FILLCELL_X2 FILLER_151_1574 ();
 FILLCELL_X1 FILLER_151_1576 ();
 FILLCELL_X32 FILLER_151_1584 ();
 FILLCELL_X32 FILLER_151_1616 ();
 FILLCELL_X2 FILLER_151_1648 ();
 FILLCELL_X1 FILLER_151_1650 ();
 FILLCELL_X16 FILLER_152_1 ();
 FILLCELL_X4 FILLER_152_17 ();
 FILLCELL_X2 FILLER_152_21 ();
 FILLCELL_X1 FILLER_152_23 ();
 FILLCELL_X2 FILLER_152_44 ();
 FILLCELL_X8 FILLER_152_53 ();
 FILLCELL_X2 FILLER_152_61 ();
 FILLCELL_X8 FILLER_152_70 ();
 FILLCELL_X16 FILLER_152_87 ();
 FILLCELL_X2 FILLER_152_110 ();
 FILLCELL_X1 FILLER_152_112 ();
 FILLCELL_X1 FILLER_152_142 ();
 FILLCELL_X1 FILLER_152_157 ();
 FILLCELL_X2 FILLER_152_178 ();
 FILLCELL_X1 FILLER_152_180 ();
 FILLCELL_X8 FILLER_152_216 ();
 FILLCELL_X4 FILLER_152_224 ();
 FILLCELL_X8 FILLER_152_235 ();
 FILLCELL_X2 FILLER_152_254 ();
 FILLCELL_X1 FILLER_152_263 ();
 FILLCELL_X4 FILLER_152_273 ();
 FILLCELL_X2 FILLER_152_277 ();
 FILLCELL_X1 FILLER_152_279 ();
 FILLCELL_X1 FILLER_152_284 ();
 FILLCELL_X4 FILLER_152_288 ();
 FILLCELL_X1 FILLER_152_292 ();
 FILLCELL_X1 FILLER_152_298 ();
 FILLCELL_X1 FILLER_152_309 ();
 FILLCELL_X8 FILLER_152_313 ();
 FILLCELL_X4 FILLER_152_321 ();
 FILLCELL_X8 FILLER_152_341 ();
 FILLCELL_X1 FILLER_152_353 ();
 FILLCELL_X2 FILLER_152_362 ();
 FILLCELL_X1 FILLER_152_364 ();
 FILLCELL_X4 FILLER_152_368 ();
 FILLCELL_X1 FILLER_152_372 ();
 FILLCELL_X8 FILLER_152_386 ();
 FILLCELL_X1 FILLER_152_394 ();
 FILLCELL_X1 FILLER_152_418 ();
 FILLCELL_X2 FILLER_152_423 ();
 FILLCELL_X1 FILLER_152_425 ();
 FILLCELL_X2 FILLER_152_452 ();
 FILLCELL_X1 FILLER_152_454 ();
 FILLCELL_X8 FILLER_152_462 ();
 FILLCELL_X1 FILLER_152_470 ();
 FILLCELL_X4 FILLER_152_485 ();
 FILLCELL_X2 FILLER_152_489 ();
 FILLCELL_X1 FILLER_152_491 ();
 FILLCELL_X2 FILLER_152_503 ();
 FILLCELL_X1 FILLER_152_505 ();
 FILLCELL_X1 FILLER_152_509 ();
 FILLCELL_X1 FILLER_152_514 ();
 FILLCELL_X2 FILLER_152_538 ();
 FILLCELL_X4 FILLER_152_545 ();
 FILLCELL_X1 FILLER_152_564 ();
 FILLCELL_X4 FILLER_152_592 ();
 FILLCELL_X4 FILLER_152_600 ();
 FILLCELL_X4 FILLER_152_619 ();
 FILLCELL_X1 FILLER_152_623 ();
 FILLCELL_X8 FILLER_152_632 ();
 FILLCELL_X1 FILLER_152_647 ();
 FILLCELL_X16 FILLER_152_655 ();
 FILLCELL_X4 FILLER_152_671 ();
 FILLCELL_X16 FILLER_152_689 ();
 FILLCELL_X8 FILLER_152_705 ();
 FILLCELL_X4 FILLER_152_713 ();
 FILLCELL_X4 FILLER_152_724 ();
 FILLCELL_X1 FILLER_152_728 ();
 FILLCELL_X1 FILLER_152_745 ();
 FILLCELL_X4 FILLER_152_758 ();
 FILLCELL_X2 FILLER_152_762 ();
 FILLCELL_X1 FILLER_152_773 ();
 FILLCELL_X1 FILLER_152_796 ();
 FILLCELL_X16 FILLER_152_846 ();
 FILLCELL_X4 FILLER_152_862 ();
 FILLCELL_X2 FILLER_152_866 ();
 FILLCELL_X1 FILLER_152_868 ();
 FILLCELL_X16 FILLER_152_876 ();
 FILLCELL_X4 FILLER_152_892 ();
 FILLCELL_X1 FILLER_152_896 ();
 FILLCELL_X16 FILLER_152_937 ();
 FILLCELL_X8 FILLER_152_953 ();
 FILLCELL_X4 FILLER_152_961 ();
 FILLCELL_X1 FILLER_152_965 ();
 FILLCELL_X2 FILLER_152_970 ();
 FILLCELL_X1 FILLER_152_972 ();
 FILLCELL_X8 FILLER_152_997 ();
 FILLCELL_X2 FILLER_152_1005 ();
 FILLCELL_X1 FILLER_152_1007 ();
 FILLCELL_X4 FILLER_152_1018 ();
 FILLCELL_X1 FILLER_152_1027 ();
 FILLCELL_X2 FILLER_152_1030 ();
 FILLCELL_X2 FILLER_152_1052 ();
 FILLCELL_X32 FILLER_152_1071 ();
 FILLCELL_X32 FILLER_152_1103 ();
 FILLCELL_X32 FILLER_152_1135 ();
 FILLCELL_X32 FILLER_152_1167 ();
 FILLCELL_X32 FILLER_152_1199 ();
 FILLCELL_X32 FILLER_152_1231 ();
 FILLCELL_X32 FILLER_152_1263 ();
 FILLCELL_X32 FILLER_152_1295 ();
 FILLCELL_X32 FILLER_152_1327 ();
 FILLCELL_X32 FILLER_152_1359 ();
 FILLCELL_X2 FILLER_152_1391 ();
 FILLCELL_X1 FILLER_152_1404 ();
 FILLCELL_X2 FILLER_152_1409 ();
 FILLCELL_X4 FILLER_152_1415 ();
 FILLCELL_X2 FILLER_152_1419 ();
 FILLCELL_X1 FILLER_152_1421 ();
 FILLCELL_X2 FILLER_152_1425 ();
 FILLCELL_X1 FILLER_152_1443 ();
 FILLCELL_X1 FILLER_152_1464 ();
 FILLCELL_X1 FILLER_152_1483 ();
 FILLCELL_X2 FILLER_152_1487 ();
 FILLCELL_X1 FILLER_152_1496 ();
 FILLCELL_X2 FILLER_152_1500 ();
 FILLCELL_X8 FILLER_152_1504 ();
 FILLCELL_X2 FILLER_152_1512 ();
 FILLCELL_X1 FILLER_152_1522 ();
 FILLCELL_X1 FILLER_152_1534 ();
 FILLCELL_X2 FILLER_152_1540 ();
 FILLCELL_X32 FILLER_152_1560 ();
 FILLCELL_X32 FILLER_152_1592 ();
 FILLCELL_X16 FILLER_152_1624 ();
 FILLCELL_X8 FILLER_152_1640 ();
 FILLCELL_X2 FILLER_152_1648 ();
 FILLCELL_X1 FILLER_152_1650 ();
 FILLCELL_X8 FILLER_153_1 ();
 FILLCELL_X4 FILLER_153_9 ();
 FILLCELL_X1 FILLER_153_13 ();
 FILLCELL_X4 FILLER_153_41 ();
 FILLCELL_X2 FILLER_153_45 ();
 FILLCELL_X8 FILLER_153_67 ();
 FILLCELL_X2 FILLER_153_75 ();
 FILLCELL_X1 FILLER_153_77 ();
 FILLCELL_X8 FILLER_153_82 ();
 FILLCELL_X4 FILLER_153_90 ();
 FILLCELL_X2 FILLER_153_121 ();
 FILLCELL_X8 FILLER_153_150 ();
 FILLCELL_X2 FILLER_153_158 ();
 FILLCELL_X1 FILLER_153_160 ();
 FILLCELL_X4 FILLER_153_168 ();
 FILLCELL_X2 FILLER_153_172 ();
 FILLCELL_X1 FILLER_153_174 ();
 FILLCELL_X16 FILLER_153_182 ();
 FILLCELL_X2 FILLER_153_198 ();
 FILLCELL_X1 FILLER_153_200 ();
 FILLCELL_X2 FILLER_153_208 ();
 FILLCELL_X1 FILLER_153_210 ();
 FILLCELL_X1 FILLER_153_218 ();
 FILLCELL_X2 FILLER_153_239 ();
 FILLCELL_X4 FILLER_153_267 ();
 FILLCELL_X2 FILLER_153_271 ();
 FILLCELL_X4 FILLER_153_280 ();
 FILLCELL_X1 FILLER_153_284 ();
 FILLCELL_X2 FILLER_153_288 ();
 FILLCELL_X1 FILLER_153_290 ();
 FILLCELL_X4 FILLER_153_296 ();
 FILLCELL_X1 FILLER_153_300 ();
 FILLCELL_X4 FILLER_153_305 ();
 FILLCELL_X4 FILLER_153_316 ();
 FILLCELL_X4 FILLER_153_360 ();
 FILLCELL_X8 FILLER_153_387 ();
 FILLCELL_X1 FILLER_153_395 ();
 FILLCELL_X1 FILLER_153_404 ();
 FILLCELL_X2 FILLER_153_437 ();
 FILLCELL_X1 FILLER_153_443 ();
 FILLCELL_X2 FILLER_153_460 ();
 FILLCELL_X1 FILLER_153_462 ();
 FILLCELL_X1 FILLER_153_488 ();
 FILLCELL_X2 FILLER_153_493 ();
 FILLCELL_X1 FILLER_153_495 ();
 FILLCELL_X2 FILLER_153_499 ();
 FILLCELL_X1 FILLER_153_509 ();
 FILLCELL_X2 FILLER_153_515 ();
 FILLCELL_X1 FILLER_153_517 ();
 FILLCELL_X4 FILLER_153_562 ();
 FILLCELL_X1 FILLER_153_566 ();
 FILLCELL_X1 FILLER_153_594 ();
 FILLCELL_X2 FILLER_153_629 ();
 FILLCELL_X1 FILLER_153_659 ();
 FILLCELL_X8 FILLER_153_694 ();
 FILLCELL_X8 FILLER_153_738 ();
 FILLCELL_X1 FILLER_153_746 ();
 FILLCELL_X8 FILLER_153_749 ();
 FILLCELL_X1 FILLER_153_757 ();
 FILLCELL_X4 FILLER_153_778 ();
 FILLCELL_X16 FILLER_153_791 ();
 FILLCELL_X8 FILLER_153_807 ();
 FILLCELL_X4 FILLER_153_815 ();
 FILLCELL_X1 FILLER_153_819 ();
 FILLCELL_X8 FILLER_153_825 ();
 FILLCELL_X4 FILLER_153_833 ();
 FILLCELL_X1 FILLER_153_837 ();
 FILLCELL_X4 FILLER_153_842 ();
 FILLCELL_X1 FILLER_153_846 ();
 FILLCELL_X32 FILLER_153_860 ();
 FILLCELL_X4 FILLER_153_892 ();
 FILLCELL_X2 FILLER_153_896 ();
 FILLCELL_X2 FILLER_153_944 ();
 FILLCELL_X2 FILLER_153_951 ();
 FILLCELL_X1 FILLER_153_953 ();
 FILLCELL_X2 FILLER_153_1004 ();
 FILLCELL_X4 FILLER_153_1033 ();
 FILLCELL_X1 FILLER_153_1037 ();
 FILLCELL_X2 FILLER_153_1045 ();
 FILLCELL_X4 FILLER_153_1051 ();
 FILLCELL_X2 FILLER_153_1055 ();
 FILLCELL_X4 FILLER_153_1062 ();
 FILLCELL_X2 FILLER_153_1066 ();
 FILLCELL_X1 FILLER_153_1068 ();
 FILLCELL_X32 FILLER_153_1096 ();
 FILLCELL_X32 FILLER_153_1128 ();
 FILLCELL_X32 FILLER_153_1160 ();
 FILLCELL_X32 FILLER_153_1192 ();
 FILLCELL_X32 FILLER_153_1224 ();
 FILLCELL_X4 FILLER_153_1256 ();
 FILLCELL_X2 FILLER_153_1260 ();
 FILLCELL_X1 FILLER_153_1262 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X32 FILLER_153_1296 ();
 FILLCELL_X32 FILLER_153_1328 ();
 FILLCELL_X8 FILLER_153_1360 ();
 FILLCELL_X2 FILLER_153_1368 ();
 FILLCELL_X4 FILLER_153_1405 ();
 FILLCELL_X2 FILLER_153_1409 ();
 FILLCELL_X16 FILLER_153_1415 ();
 FILLCELL_X8 FILLER_153_1431 ();
 FILLCELL_X1 FILLER_153_1439 ();
 FILLCELL_X1 FILLER_153_1446 ();
 FILLCELL_X8 FILLER_153_1451 ();
 FILLCELL_X4 FILLER_153_1459 ();
 FILLCELL_X2 FILLER_153_1463 ();
 FILLCELL_X1 FILLER_153_1465 ();
 FILLCELL_X8 FILLER_153_1475 ();
 FILLCELL_X2 FILLER_153_1483 ();
 FILLCELL_X1 FILLER_153_1488 ();
 FILLCELL_X1 FILLER_153_1493 ();
 FILLCELL_X2 FILLER_153_1500 ();
 FILLCELL_X16 FILLER_153_1509 ();
 FILLCELL_X4 FILLER_153_1525 ();
 FILLCELL_X1 FILLER_153_1529 ();
 FILLCELL_X2 FILLER_153_1533 ();
 FILLCELL_X4 FILLER_153_1552 ();
 FILLCELL_X1 FILLER_153_1556 ();
 FILLCELL_X2 FILLER_153_1564 ();
 FILLCELL_X32 FILLER_153_1591 ();
 FILLCELL_X16 FILLER_153_1623 ();
 FILLCELL_X8 FILLER_153_1639 ();
 FILLCELL_X4 FILLER_153_1647 ();
 FILLCELL_X16 FILLER_154_1 ();
 FILLCELL_X2 FILLER_154_17 ();
 FILLCELL_X4 FILLER_154_58 ();
 FILLCELL_X2 FILLER_154_62 ();
 FILLCELL_X2 FILLER_154_100 ();
 FILLCELL_X1 FILLER_154_102 ();
 FILLCELL_X2 FILLER_154_123 ();
 FILLCELL_X1 FILLER_154_125 ();
 FILLCELL_X8 FILLER_154_138 ();
 FILLCELL_X4 FILLER_154_159 ();
 FILLCELL_X1 FILLER_154_170 ();
 FILLCELL_X8 FILLER_154_198 ();
 FILLCELL_X4 FILLER_154_206 ();
 FILLCELL_X2 FILLER_154_210 ();
 FILLCELL_X1 FILLER_154_212 ();
 FILLCELL_X1 FILLER_154_234 ();
 FILLCELL_X2 FILLER_154_242 ();
 FILLCELL_X1 FILLER_154_244 ();
 FILLCELL_X1 FILLER_154_310 ();
 FILLCELL_X16 FILLER_154_336 ();
 FILLCELL_X4 FILLER_154_388 ();
 FILLCELL_X2 FILLER_154_392 ();
 FILLCELL_X1 FILLER_154_394 ();
 FILLCELL_X2 FILLER_154_420 ();
 FILLCELL_X4 FILLER_154_458 ();
 FILLCELL_X1 FILLER_154_462 ();
 FILLCELL_X4 FILLER_154_470 ();
 FILLCELL_X1 FILLER_154_478 ();
 FILLCELL_X2 FILLER_154_506 ();
 FILLCELL_X2 FILLER_154_513 ();
 FILLCELL_X1 FILLER_154_522 ();
 FILLCELL_X2 FILLER_154_572 ();
 FILLCELL_X8 FILLER_154_594 ();
 FILLCELL_X4 FILLER_154_602 ();
 FILLCELL_X1 FILLER_154_630 ();
 FILLCELL_X2 FILLER_154_632 ();
 FILLCELL_X1 FILLER_154_637 ();
 FILLCELL_X8 FILLER_154_645 ();
 FILLCELL_X4 FILLER_154_653 ();
 FILLCELL_X1 FILLER_154_657 ();
 FILLCELL_X8 FILLER_154_663 ();
 FILLCELL_X2 FILLER_154_671 ();
 FILLCELL_X1 FILLER_154_693 ();
 FILLCELL_X1 FILLER_154_719 ();
 FILLCELL_X2 FILLER_154_724 ();
 FILLCELL_X8 FILLER_154_733 ();
 FILLCELL_X4 FILLER_154_741 ();
 FILLCELL_X1 FILLER_154_745 ();
 FILLCELL_X2 FILLER_154_750 ();
 FILLCELL_X2 FILLER_154_757 ();
 FILLCELL_X4 FILLER_154_763 ();
 FILLCELL_X2 FILLER_154_790 ();
 FILLCELL_X2 FILLER_154_812 ();
 FILLCELL_X1 FILLER_154_814 ();
 FILLCELL_X2 FILLER_154_818 ();
 FILLCELL_X4 FILLER_154_825 ();
 FILLCELL_X4 FILLER_154_836 ();
 FILLCELL_X2 FILLER_154_840 ();
 FILLCELL_X1 FILLER_154_842 ();
 FILLCELL_X8 FILLER_154_914 ();
 FILLCELL_X1 FILLER_154_949 ();
 FILLCELL_X16 FILLER_154_1031 ();
 FILLCELL_X4 FILLER_154_1047 ();
 FILLCELL_X2 FILLER_154_1051 ();
 FILLCELL_X1 FILLER_154_1053 ();
 FILLCELL_X1 FILLER_154_1060 ();
 FILLCELL_X16 FILLER_154_1093 ();
 FILLCELL_X8 FILLER_154_1109 ();
 FILLCELL_X4 FILLER_154_1117 ();
 FILLCELL_X2 FILLER_154_1121 ();
 FILLCELL_X32 FILLER_154_1133 ();
 FILLCELL_X32 FILLER_154_1165 ();
 FILLCELL_X32 FILLER_154_1197 ();
 FILLCELL_X32 FILLER_154_1229 ();
 FILLCELL_X32 FILLER_154_1261 ();
 FILLCELL_X32 FILLER_154_1293 ();
 FILLCELL_X32 FILLER_154_1325 ();
 FILLCELL_X16 FILLER_154_1357 ();
 FILLCELL_X4 FILLER_154_1373 ();
 FILLCELL_X2 FILLER_154_1377 ();
 FILLCELL_X1 FILLER_154_1379 ();
 FILLCELL_X1 FILLER_154_1400 ();
 FILLCELL_X4 FILLER_154_1420 ();
 FILLCELL_X2 FILLER_154_1424 ();
 FILLCELL_X1 FILLER_154_1426 ();
 FILLCELL_X8 FILLER_154_1431 ();
 FILLCELL_X1 FILLER_154_1439 ();
 FILLCELL_X4 FILLER_154_1445 ();
 FILLCELL_X8 FILLER_154_1452 ();
 FILLCELL_X4 FILLER_154_1460 ();
 FILLCELL_X4 FILLER_154_1467 ();
 FILLCELL_X1 FILLER_154_1471 ();
 FILLCELL_X8 FILLER_154_1480 ();
 FILLCELL_X1 FILLER_154_1488 ();
 FILLCELL_X2 FILLER_154_1499 ();
 FILLCELL_X1 FILLER_154_1501 ();
 FILLCELL_X4 FILLER_154_1525 ();
 FILLCELL_X2 FILLER_154_1529 ();
 FILLCELL_X32 FILLER_154_1558 ();
 FILLCELL_X32 FILLER_154_1590 ();
 FILLCELL_X16 FILLER_154_1622 ();
 FILLCELL_X8 FILLER_154_1638 ();
 FILLCELL_X4 FILLER_154_1646 ();
 FILLCELL_X1 FILLER_154_1650 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X2 FILLER_155_33 ();
 FILLCELL_X1 FILLER_155_35 ();
 FILLCELL_X1 FILLER_155_63 ();
 FILLCELL_X2 FILLER_155_79 ();
 FILLCELL_X2 FILLER_155_104 ();
 FILLCELL_X2 FILLER_155_126 ();
 FILLCELL_X2 FILLER_155_137 ();
 FILLCELL_X4 FILLER_155_146 ();
 FILLCELL_X2 FILLER_155_170 ();
 FILLCELL_X2 FILLER_155_241 ();
 FILLCELL_X1 FILLER_155_243 ();
 FILLCELL_X8 FILLER_155_247 ();
 FILLCELL_X4 FILLER_155_266 ();
 FILLCELL_X1 FILLER_155_270 ();
 FILLCELL_X4 FILLER_155_338 ();
 FILLCELL_X4 FILLER_155_362 ();
 FILLCELL_X2 FILLER_155_366 ();
 FILLCELL_X1 FILLER_155_372 ();
 FILLCELL_X8 FILLER_155_383 ();
 FILLCELL_X2 FILLER_155_391 ();
 FILLCELL_X16 FILLER_155_416 ();
 FILLCELL_X8 FILLER_155_432 ();
 FILLCELL_X4 FILLER_155_440 ();
 FILLCELL_X16 FILLER_155_461 ();
 FILLCELL_X8 FILLER_155_477 ();
 FILLCELL_X4 FILLER_155_485 ();
 FILLCELL_X1 FILLER_155_542 ();
 FILLCELL_X1 FILLER_155_550 ();
 FILLCELL_X2 FILLER_155_574 ();
 FILLCELL_X1 FILLER_155_576 ();
 FILLCELL_X2 FILLER_155_581 ();
 FILLCELL_X8 FILLER_155_586 ();
 FILLCELL_X4 FILLER_155_594 ();
 FILLCELL_X1 FILLER_155_598 ();
 FILLCELL_X4 FILLER_155_606 ();
 FILLCELL_X2 FILLER_155_610 ();
 FILLCELL_X1 FILLER_155_612 ();
 FILLCELL_X4 FILLER_155_660 ();
 FILLCELL_X4 FILLER_155_669 ();
 FILLCELL_X1 FILLER_155_673 ();
 FILLCELL_X4 FILLER_155_681 ();
 FILLCELL_X4 FILLER_155_705 ();
 FILLCELL_X2 FILLER_155_709 ();
 FILLCELL_X1 FILLER_155_743 ();
 FILLCELL_X8 FILLER_155_767 ();
 FILLCELL_X1 FILLER_155_775 ();
 FILLCELL_X4 FILLER_155_783 ();
 FILLCELL_X2 FILLER_155_787 ();
 FILLCELL_X1 FILLER_155_789 ();
 FILLCELL_X4 FILLER_155_797 ();
 FILLCELL_X2 FILLER_155_825 ();
 FILLCELL_X4 FILLER_155_847 ();
 FILLCELL_X2 FILLER_155_851 ();
 FILLCELL_X1 FILLER_155_853 ();
 FILLCELL_X8 FILLER_155_874 ();
 FILLCELL_X2 FILLER_155_882 ();
 FILLCELL_X1 FILLER_155_884 ();
 FILLCELL_X4 FILLER_155_930 ();
 FILLCELL_X2 FILLER_155_941 ();
 FILLCELL_X2 FILLER_155_952 ();
 FILLCELL_X2 FILLER_155_961 ();
 FILLCELL_X2 FILLER_155_970 ();
 FILLCELL_X1 FILLER_155_972 ();
 FILLCELL_X4 FILLER_155_982 ();
 FILLCELL_X1 FILLER_155_990 ();
 FILLCELL_X2 FILLER_155_1000 ();
 FILLCELL_X1 FILLER_155_1009 ();
 FILLCELL_X2 FILLER_155_1030 ();
 FILLCELL_X4 FILLER_155_1039 ();
 FILLCELL_X2 FILLER_155_1043 ();
 FILLCELL_X2 FILLER_155_1072 ();
 FILLCELL_X32 FILLER_155_1094 ();
 FILLCELL_X32 FILLER_155_1126 ();
 FILLCELL_X32 FILLER_155_1158 ();
 FILLCELL_X32 FILLER_155_1190 ();
 FILLCELL_X32 FILLER_155_1222 ();
 FILLCELL_X8 FILLER_155_1254 ();
 FILLCELL_X1 FILLER_155_1262 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X32 FILLER_155_1296 ();
 FILLCELL_X32 FILLER_155_1328 ();
 FILLCELL_X32 FILLER_155_1360 ();
 FILLCELL_X8 FILLER_155_1392 ();
 FILLCELL_X4 FILLER_155_1420 ();
 FILLCELL_X2 FILLER_155_1424 ();
 FILLCELL_X1 FILLER_155_1471 ();
 FILLCELL_X1 FILLER_155_1480 ();
 FILLCELL_X2 FILLER_155_1497 ();
 FILLCELL_X1 FILLER_155_1499 ();
 FILLCELL_X8 FILLER_155_1506 ();
 FILLCELL_X1 FILLER_155_1514 ();
 FILLCELL_X8 FILLER_155_1520 ();
 FILLCELL_X4 FILLER_155_1528 ();
 FILLCELL_X2 FILLER_155_1532 ();
 FILLCELL_X1 FILLER_155_1534 ();
 FILLCELL_X2 FILLER_155_1553 ();
 FILLCELL_X32 FILLER_155_1558 ();
 FILLCELL_X32 FILLER_155_1590 ();
 FILLCELL_X16 FILLER_155_1622 ();
 FILLCELL_X8 FILLER_155_1638 ();
 FILLCELL_X4 FILLER_155_1646 ();
 FILLCELL_X1 FILLER_155_1650 ();
 FILLCELL_X16 FILLER_156_1 ();
 FILLCELL_X8 FILLER_156_17 ();
 FILLCELL_X4 FILLER_156_25 ();
 FILLCELL_X1 FILLER_156_29 ();
 FILLCELL_X2 FILLER_156_50 ();
 FILLCELL_X2 FILLER_156_59 ();
 FILLCELL_X1 FILLER_156_61 ();
 FILLCELL_X8 FILLER_156_75 ();
 FILLCELL_X1 FILLER_156_83 ();
 FILLCELL_X4 FILLER_156_97 ();
 FILLCELL_X4 FILLER_156_108 ();
 FILLCELL_X2 FILLER_156_112 ();
 FILLCELL_X1 FILLER_156_176 ();
 FILLCELL_X2 FILLER_156_184 ();
 FILLCELL_X2 FILLER_156_203 ();
 FILLCELL_X1 FILLER_156_205 ();
 FILLCELL_X1 FILLER_156_213 ();
 FILLCELL_X1 FILLER_156_221 ();
 FILLCELL_X2 FILLER_156_255 ();
 FILLCELL_X2 FILLER_156_261 ();
 FILLCELL_X8 FILLER_156_306 ();
 FILLCELL_X4 FILLER_156_337 ();
 FILLCELL_X2 FILLER_156_341 ();
 FILLCELL_X8 FILLER_156_350 ();
 FILLCELL_X2 FILLER_156_358 ();
 FILLCELL_X2 FILLER_156_385 ();
 FILLCELL_X1 FILLER_156_405 ();
 FILLCELL_X2 FILLER_156_442 ();
 FILLCELL_X2 FILLER_156_464 ();
 FILLCELL_X1 FILLER_156_466 ();
 FILLCELL_X4 FILLER_156_485 ();
 FILLCELL_X8 FILLER_156_506 ();
 FILLCELL_X2 FILLER_156_514 ();
 FILLCELL_X8 FILLER_156_534 ();
 FILLCELL_X2 FILLER_156_542 ();
 FILLCELL_X1 FILLER_156_544 ();
 FILLCELL_X1 FILLER_156_574 ();
 FILLCELL_X1 FILLER_156_599 ();
 FILLCELL_X8 FILLER_156_607 ();
 FILLCELL_X2 FILLER_156_615 ();
 FILLCELL_X1 FILLER_156_630 ();
 FILLCELL_X1 FILLER_156_639 ();
 FILLCELL_X2 FILLER_156_669 ();
 FILLCELL_X1 FILLER_156_698 ();
 FILLCELL_X8 FILLER_156_719 ();
 FILLCELL_X2 FILLER_156_727 ();
 FILLCELL_X8 FILLER_156_736 ();
 FILLCELL_X2 FILLER_156_744 ();
 FILLCELL_X1 FILLER_156_753 ();
 FILLCELL_X8 FILLER_156_791 ();
 FILLCELL_X4 FILLER_156_799 ();
 FILLCELL_X2 FILLER_156_803 ();
 FILLCELL_X2 FILLER_156_844 ();
 FILLCELL_X1 FILLER_156_846 ();
 FILLCELL_X8 FILLER_156_859 ();
 FILLCELL_X4 FILLER_156_875 ();
 FILLCELL_X1 FILLER_156_879 ();
 FILLCELL_X1 FILLER_156_889 ();
 FILLCELL_X1 FILLER_156_897 ();
 FILLCELL_X2 FILLER_156_907 ();
 FILLCELL_X1 FILLER_156_916 ();
 FILLCELL_X2 FILLER_156_921 ();
 FILLCELL_X2 FILLER_156_928 ();
 FILLCELL_X2 FILLER_156_937 ();
 FILLCELL_X4 FILLER_156_959 ();
 FILLCELL_X2 FILLER_156_963 ();
 FILLCELL_X1 FILLER_156_965 ();
 FILLCELL_X8 FILLER_156_1021 ();
 FILLCELL_X2 FILLER_156_1054 ();
 FILLCELL_X1 FILLER_156_1056 ();
 FILLCELL_X2 FILLER_156_1069 ();
 FILLCELL_X1 FILLER_156_1071 ();
 FILLCELL_X32 FILLER_156_1079 ();
 FILLCELL_X32 FILLER_156_1111 ();
 FILLCELL_X32 FILLER_156_1143 ();
 FILLCELL_X32 FILLER_156_1175 ();
 FILLCELL_X32 FILLER_156_1207 ();
 FILLCELL_X32 FILLER_156_1239 ();
 FILLCELL_X32 FILLER_156_1271 ();
 FILLCELL_X32 FILLER_156_1303 ();
 FILLCELL_X32 FILLER_156_1335 ();
 FILLCELL_X16 FILLER_156_1367 ();
 FILLCELL_X8 FILLER_156_1383 ();
 FILLCELL_X1 FILLER_156_1391 ();
 FILLCELL_X1 FILLER_156_1405 ();
 FILLCELL_X2 FILLER_156_1410 ();
 FILLCELL_X2 FILLER_156_1415 ();
 FILLCELL_X2 FILLER_156_1435 ();
 FILLCELL_X1 FILLER_156_1437 ();
 FILLCELL_X8 FILLER_156_1442 ();
 FILLCELL_X1 FILLER_156_1464 ();
 FILLCELL_X2 FILLER_156_1476 ();
 FILLCELL_X1 FILLER_156_1478 ();
 FILLCELL_X4 FILLER_156_1482 ();
 FILLCELL_X1 FILLER_156_1486 ();
 FILLCELL_X4 FILLER_156_1491 ();
 FILLCELL_X2 FILLER_156_1495 ();
 FILLCELL_X8 FILLER_156_1522 ();
 FILLCELL_X4 FILLER_156_1530 ();
 FILLCELL_X4 FILLER_156_1551 ();
 FILLCELL_X1 FILLER_156_1555 ();
 FILLCELL_X32 FILLER_156_1572 ();
 FILLCELL_X32 FILLER_156_1604 ();
 FILLCELL_X8 FILLER_156_1636 ();
 FILLCELL_X4 FILLER_156_1644 ();
 FILLCELL_X2 FILLER_156_1648 ();
 FILLCELL_X1 FILLER_156_1650 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X4 FILLER_157_33 ();
 FILLCELL_X2 FILLER_157_64 ();
 FILLCELL_X8 FILLER_157_98 ();
 FILLCELL_X2 FILLER_157_106 ();
 FILLCELL_X1 FILLER_157_108 ();
 FILLCELL_X1 FILLER_157_129 ();
 FILLCELL_X2 FILLER_157_137 ();
 FILLCELL_X1 FILLER_157_139 ();
 FILLCELL_X1 FILLER_157_151 ();
 FILLCELL_X1 FILLER_157_161 ();
 FILLCELL_X1 FILLER_157_169 ();
 FILLCELL_X2 FILLER_157_190 ();
 FILLCELL_X8 FILLER_157_199 ();
 FILLCELL_X2 FILLER_157_207 ();
 FILLCELL_X1 FILLER_157_209 ();
 FILLCELL_X4 FILLER_157_233 ();
 FILLCELL_X1 FILLER_157_237 ();
 FILLCELL_X4 FILLER_157_279 ();
 FILLCELL_X2 FILLER_157_286 ();
 FILLCELL_X8 FILLER_157_312 ();
 FILLCELL_X2 FILLER_157_320 ();
 FILLCELL_X1 FILLER_157_326 ();
 FILLCELL_X1 FILLER_157_339 ();
 FILLCELL_X1 FILLER_157_360 ();
 FILLCELL_X1 FILLER_157_365 ();
 FILLCELL_X1 FILLER_157_406 ();
 FILLCELL_X4 FILLER_157_427 ();
 FILLCELL_X8 FILLER_157_434 ();
 FILLCELL_X1 FILLER_157_442 ();
 FILLCELL_X2 FILLER_157_450 ();
 FILLCELL_X8 FILLER_157_456 ();
 FILLCELL_X1 FILLER_157_464 ();
 FILLCELL_X1 FILLER_157_489 ();
 FILLCELL_X2 FILLER_157_514 ();
 FILLCELL_X1 FILLER_157_516 ();
 FILLCELL_X1 FILLER_157_542 ();
 FILLCELL_X4 FILLER_157_550 ();
 FILLCELL_X2 FILLER_157_554 ();
 FILLCELL_X4 FILLER_157_563 ();
 FILLCELL_X1 FILLER_157_567 ();
 FILLCELL_X2 FILLER_157_574 ();
 FILLCELL_X1 FILLER_157_576 ();
 FILLCELL_X8 FILLER_157_611 ();
 FILLCELL_X2 FILLER_157_619 ();
 FILLCELL_X1 FILLER_157_621 ();
 FILLCELL_X1 FILLER_157_642 ();
 FILLCELL_X8 FILLER_157_677 ();
 FILLCELL_X4 FILLER_157_685 ();
 FILLCELL_X2 FILLER_157_689 ();
 FILLCELL_X1 FILLER_157_691 ();
 FILLCELL_X2 FILLER_157_719 ();
 FILLCELL_X1 FILLER_157_721 ();
 FILLCELL_X4 FILLER_157_742 ();
 FILLCELL_X4 FILLER_157_786 ();
 FILLCELL_X2 FILLER_157_790 ();
 FILLCELL_X1 FILLER_157_792 ();
 FILLCELL_X4 FILLER_157_800 ();
 FILLCELL_X2 FILLER_157_804 ();
 FILLCELL_X2 FILLER_157_818 ();
 FILLCELL_X16 FILLER_157_822 ();
 FILLCELL_X4 FILLER_157_838 ();
 FILLCELL_X2 FILLER_157_842 ();
 FILLCELL_X1 FILLER_157_844 ();
 FILLCELL_X2 FILLER_157_852 ();
 FILLCELL_X4 FILLER_157_899 ();
 FILLCELL_X1 FILLER_157_903 ();
 FILLCELL_X4 FILLER_157_956 ();
 FILLCELL_X2 FILLER_157_960 ();
 FILLCELL_X16 FILLER_157_998 ();
 FILLCELL_X1 FILLER_157_1014 ();
 FILLCELL_X2 FILLER_157_1037 ();
 FILLCELL_X8 FILLER_157_1044 ();
 FILLCELL_X8 FILLER_157_1061 ();
 FILLCELL_X2 FILLER_157_1069 ();
 FILLCELL_X1 FILLER_157_1071 ();
 FILLCELL_X32 FILLER_157_1092 ();
 FILLCELL_X32 FILLER_157_1124 ();
 FILLCELL_X32 FILLER_157_1156 ();
 FILLCELL_X32 FILLER_157_1188 ();
 FILLCELL_X32 FILLER_157_1220 ();
 FILLCELL_X8 FILLER_157_1252 ();
 FILLCELL_X2 FILLER_157_1260 ();
 FILLCELL_X1 FILLER_157_1262 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X32 FILLER_157_1296 ();
 FILLCELL_X32 FILLER_157_1328 ();
 FILLCELL_X16 FILLER_157_1360 ();
 FILLCELL_X8 FILLER_157_1376 ();
 FILLCELL_X2 FILLER_157_1384 ();
 FILLCELL_X1 FILLER_157_1386 ();
 FILLCELL_X1 FILLER_157_1435 ();
 FILLCELL_X1 FILLER_157_1444 ();
 FILLCELL_X2 FILLER_157_1450 ();
 FILLCELL_X8 FILLER_157_1459 ();
 FILLCELL_X1 FILLER_157_1467 ();
 FILLCELL_X8 FILLER_157_1486 ();
 FILLCELL_X8 FILLER_157_1503 ();
 FILLCELL_X4 FILLER_157_1511 ();
 FILLCELL_X2 FILLER_157_1519 ();
 FILLCELL_X4 FILLER_157_1538 ();
 FILLCELL_X1 FILLER_157_1558 ();
 FILLCELL_X32 FILLER_157_1566 ();
 FILLCELL_X32 FILLER_157_1598 ();
 FILLCELL_X16 FILLER_157_1630 ();
 FILLCELL_X4 FILLER_157_1646 ();
 FILLCELL_X1 FILLER_157_1650 ();
 FILLCELL_X16 FILLER_158_1 ();
 FILLCELL_X8 FILLER_158_17 ();
 FILLCELL_X2 FILLER_158_74 ();
 FILLCELL_X4 FILLER_158_96 ();
 FILLCELL_X2 FILLER_158_100 ();
 FILLCELL_X1 FILLER_158_102 ();
 FILLCELL_X8 FILLER_158_116 ();
 FILLCELL_X1 FILLER_158_124 ();
 FILLCELL_X2 FILLER_158_145 ();
 FILLCELL_X4 FILLER_158_156 ();
 FILLCELL_X2 FILLER_158_160 ();
 FILLCELL_X16 FILLER_158_203 ();
 FILLCELL_X4 FILLER_158_219 ();
 FILLCELL_X2 FILLER_158_223 ();
 FILLCELL_X2 FILLER_158_245 ();
 FILLCELL_X2 FILLER_158_250 ();
 FILLCELL_X1 FILLER_158_252 ();
 FILLCELL_X1 FILLER_158_282 ();
 FILLCELL_X2 FILLER_158_298 ();
 FILLCELL_X16 FILLER_158_307 ();
 FILLCELL_X4 FILLER_158_323 ();
 FILLCELL_X2 FILLER_158_327 ();
 FILLCELL_X1 FILLER_158_329 ();
 FILLCELL_X2 FILLER_158_350 ();
 FILLCELL_X1 FILLER_158_352 ();
 FILLCELL_X8 FILLER_158_356 ();
 FILLCELL_X2 FILLER_158_364 ();
 FILLCELL_X1 FILLER_158_366 ();
 FILLCELL_X2 FILLER_158_371 ();
 FILLCELL_X1 FILLER_158_373 ();
 FILLCELL_X1 FILLER_158_377 ();
 FILLCELL_X2 FILLER_158_383 ();
 FILLCELL_X8 FILLER_158_388 ();
 FILLCELL_X4 FILLER_158_396 ();
 FILLCELL_X1 FILLER_158_404 ();
 FILLCELL_X4 FILLER_158_408 ();
 FILLCELL_X2 FILLER_158_416 ();
 FILLCELL_X1 FILLER_158_418 ();
 FILLCELL_X4 FILLER_158_426 ();
 FILLCELL_X2 FILLER_158_430 ();
 FILLCELL_X1 FILLER_158_432 ();
 FILLCELL_X4 FILLER_158_453 ();
 FILLCELL_X2 FILLER_158_477 ();
 FILLCELL_X1 FILLER_158_502 ();
 FILLCELL_X2 FILLER_158_511 ();
 FILLCELL_X1 FILLER_158_536 ();
 FILLCELL_X4 FILLER_158_557 ();
 FILLCELL_X2 FILLER_158_561 ();
 FILLCELL_X1 FILLER_158_563 ();
 FILLCELL_X4 FILLER_158_584 ();
 FILLCELL_X8 FILLER_158_594 ();
 FILLCELL_X1 FILLER_158_602 ();
 FILLCELL_X2 FILLER_158_610 ();
 FILLCELL_X2 FILLER_158_619 ();
 FILLCELL_X2 FILLER_158_628 ();
 FILLCELL_X1 FILLER_158_630 ();
 FILLCELL_X8 FILLER_158_632 ();
 FILLCELL_X1 FILLER_158_640 ();
 FILLCELL_X1 FILLER_158_648 ();
 FILLCELL_X4 FILLER_158_664 ();
 FILLCELL_X2 FILLER_158_668 ();
 FILLCELL_X8 FILLER_158_675 ();
 FILLCELL_X1 FILLER_158_683 ();
 FILLCELL_X2 FILLER_158_698 ();
 FILLCELL_X1 FILLER_158_703 ();
 FILLCELL_X8 FILLER_158_711 ();
 FILLCELL_X2 FILLER_158_719 ();
 FILLCELL_X1 FILLER_158_721 ();
 FILLCELL_X2 FILLER_158_742 ();
 FILLCELL_X1 FILLER_158_744 ();
 FILLCELL_X2 FILLER_158_750 ();
 FILLCELL_X1 FILLER_158_752 ();
 FILLCELL_X2 FILLER_158_759 ();
 FILLCELL_X1 FILLER_158_761 ();
 FILLCELL_X4 FILLER_158_770 ();
 FILLCELL_X2 FILLER_158_774 ();
 FILLCELL_X2 FILLER_158_783 ();
 FILLCELL_X4 FILLER_158_825 ();
 FILLCELL_X2 FILLER_158_829 ();
 FILLCELL_X8 FILLER_158_833 ();
 FILLCELL_X4 FILLER_158_841 ();
 FILLCELL_X2 FILLER_158_852 ();
 FILLCELL_X1 FILLER_158_854 ();
 FILLCELL_X16 FILLER_158_860 ();
 FILLCELL_X4 FILLER_158_876 ();
 FILLCELL_X8 FILLER_158_900 ();
 FILLCELL_X1 FILLER_158_908 ();
 FILLCELL_X1 FILLER_158_916 ();
 FILLCELL_X32 FILLER_158_936 ();
 FILLCELL_X4 FILLER_158_968 ();
 FILLCELL_X2 FILLER_158_972 ();
 FILLCELL_X1 FILLER_158_974 ();
 FILLCELL_X4 FILLER_158_1002 ();
 FILLCELL_X8 FILLER_158_1018 ();
 FILLCELL_X2 FILLER_158_1053 ();
 FILLCELL_X4 FILLER_158_1062 ();
 FILLCELL_X2 FILLER_158_1066 ();
 FILLCELL_X32 FILLER_158_1088 ();
 FILLCELL_X32 FILLER_158_1120 ();
 FILLCELL_X16 FILLER_158_1152 ();
 FILLCELL_X8 FILLER_158_1168 ();
 FILLCELL_X4 FILLER_158_1176 ();
 FILLCELL_X2 FILLER_158_1180 ();
 FILLCELL_X32 FILLER_158_1191 ();
 FILLCELL_X32 FILLER_158_1223 ();
 FILLCELL_X32 FILLER_158_1255 ();
 FILLCELL_X32 FILLER_158_1287 ();
 FILLCELL_X32 FILLER_158_1319 ();
 FILLCELL_X32 FILLER_158_1351 ();
 FILLCELL_X8 FILLER_158_1383 ();
 FILLCELL_X1 FILLER_158_1403 ();
 FILLCELL_X4 FILLER_158_1416 ();
 FILLCELL_X1 FILLER_158_1420 ();
 FILLCELL_X8 FILLER_158_1427 ();
 FILLCELL_X2 FILLER_158_1435 ();
 FILLCELL_X1 FILLER_158_1437 ();
 FILLCELL_X8 FILLER_158_1441 ();
 FILLCELL_X1 FILLER_158_1449 ();
 FILLCELL_X2 FILLER_158_1458 ();
 FILLCELL_X4 FILLER_158_1476 ();
 FILLCELL_X2 FILLER_158_1480 ();
 FILLCELL_X4 FILLER_158_1486 ();
 FILLCELL_X4 FILLER_158_1508 ();
 FILLCELL_X1 FILLER_158_1512 ();
 FILLCELL_X4 FILLER_158_1522 ();
 FILLCELL_X4 FILLER_158_1539 ();
 FILLCELL_X2 FILLER_158_1543 ();
 FILLCELL_X1 FILLER_158_1545 ();
 FILLCELL_X4 FILLER_158_1551 ();
 FILLCELL_X1 FILLER_158_1555 ();
 FILLCELL_X32 FILLER_158_1563 ();
 FILLCELL_X32 FILLER_158_1595 ();
 FILLCELL_X16 FILLER_158_1627 ();
 FILLCELL_X8 FILLER_158_1643 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X8 FILLER_159_33 ();
 FILLCELL_X1 FILLER_159_41 ();
 FILLCELL_X8 FILLER_159_65 ();
 FILLCELL_X1 FILLER_159_80 ();
 FILLCELL_X8 FILLER_159_90 ();
 FILLCELL_X4 FILLER_159_98 ();
 FILLCELL_X1 FILLER_159_102 ();
 FILLCELL_X4 FILLER_159_132 ();
 FILLCELL_X2 FILLER_159_136 ();
 FILLCELL_X1 FILLER_159_138 ();
 FILLCELL_X2 FILLER_159_198 ();
 FILLCELL_X1 FILLER_159_200 ();
 FILLCELL_X8 FILLER_159_215 ();
 FILLCELL_X8 FILLER_159_237 ();
 FILLCELL_X4 FILLER_159_245 ();
 FILLCELL_X2 FILLER_159_256 ();
 FILLCELL_X4 FILLER_159_299 ();
 FILLCELL_X2 FILLER_159_303 ();
 FILLCELL_X1 FILLER_159_309 ();
 FILLCELL_X4 FILLER_159_327 ();
 FILLCELL_X2 FILLER_159_331 ();
 FILLCELL_X1 FILLER_159_333 ();
 FILLCELL_X8 FILLER_159_363 ();
 FILLCELL_X4 FILLER_159_371 ();
 FILLCELL_X1 FILLER_159_375 ();
 FILLCELL_X8 FILLER_159_385 ();
 FILLCELL_X4 FILLER_159_393 ();
 FILLCELL_X2 FILLER_159_397 ();
 FILLCELL_X1 FILLER_159_399 ();
 FILLCELL_X1 FILLER_159_404 ();
 FILLCELL_X8 FILLER_159_408 ();
 FILLCELL_X8 FILLER_159_443 ();
 FILLCELL_X1 FILLER_159_458 ();
 FILLCELL_X1 FILLER_159_466 ();
 FILLCELL_X4 FILLER_159_470 ();
 FILLCELL_X1 FILLER_159_481 ();
 FILLCELL_X1 FILLER_159_486 ();
 FILLCELL_X2 FILLER_159_491 ();
 FILLCELL_X1 FILLER_159_498 ();
 FILLCELL_X2 FILLER_159_505 ();
 FILLCELL_X1 FILLER_159_517 ();
 FILLCELL_X2 FILLER_159_522 ();
 FILLCELL_X1 FILLER_159_524 ();
 FILLCELL_X4 FILLER_159_528 ();
 FILLCELL_X2 FILLER_159_532 ();
 FILLCELL_X4 FILLER_159_541 ();
 FILLCELL_X1 FILLER_159_549 ();
 FILLCELL_X4 FILLER_159_553 ();
 FILLCELL_X2 FILLER_159_557 ();
 FILLCELL_X1 FILLER_159_559 ();
 FILLCELL_X2 FILLER_159_599 ();
 FILLCELL_X4 FILLER_159_628 ();
 FILLCELL_X8 FILLER_159_657 ();
 FILLCELL_X4 FILLER_159_665 ();
 FILLCELL_X1 FILLER_159_669 ();
 FILLCELL_X8 FILLER_159_677 ();
 FILLCELL_X4 FILLER_159_685 ();
 FILLCELL_X1 FILLER_159_689 ();
 FILLCELL_X8 FILLER_159_715 ();
 FILLCELL_X4 FILLER_159_723 ();
 FILLCELL_X2 FILLER_159_727 ();
 FILLCELL_X4 FILLER_159_750 ();
 FILLCELL_X4 FILLER_159_777 ();
 FILLCELL_X2 FILLER_159_781 ();
 FILLCELL_X1 FILLER_159_783 ();
 FILLCELL_X4 FILLER_159_804 ();
 FILLCELL_X8 FILLER_159_868 ();
 FILLCELL_X4 FILLER_159_876 ();
 FILLCELL_X1 FILLER_159_880 ();
 FILLCELL_X16 FILLER_159_897 ();
 FILLCELL_X2 FILLER_159_913 ();
 FILLCELL_X1 FILLER_159_920 ();
 FILLCELL_X1 FILLER_159_946 ();
 FILLCELL_X4 FILLER_159_974 ();
 FILLCELL_X2 FILLER_159_987 ();
 FILLCELL_X1 FILLER_159_989 ();
 FILLCELL_X2 FILLER_159_999 ();
 FILLCELL_X4 FILLER_159_1021 ();
 FILLCELL_X4 FILLER_159_1045 ();
 FILLCELL_X4 FILLER_159_1054 ();
 FILLCELL_X8 FILLER_159_1078 ();
 FILLCELL_X1 FILLER_159_1086 ();
 FILLCELL_X32 FILLER_159_1097 ();
 FILLCELL_X32 FILLER_159_1129 ();
 FILLCELL_X32 FILLER_159_1161 ();
 FILLCELL_X32 FILLER_159_1193 ();
 FILLCELL_X32 FILLER_159_1225 ();
 FILLCELL_X4 FILLER_159_1257 ();
 FILLCELL_X2 FILLER_159_1261 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X32 FILLER_159_1296 ();
 FILLCELL_X32 FILLER_159_1328 ();
 FILLCELL_X32 FILLER_159_1360 ();
 FILLCELL_X8 FILLER_159_1392 ();
 FILLCELL_X2 FILLER_159_1400 ();
 FILLCELL_X1 FILLER_159_1407 ();
 FILLCELL_X2 FILLER_159_1449 ();
 FILLCELL_X1 FILLER_159_1451 ();
 FILLCELL_X2 FILLER_159_1459 ();
 FILLCELL_X1 FILLER_159_1461 ();
 FILLCELL_X1 FILLER_159_1475 ();
 FILLCELL_X1 FILLER_159_1486 ();
 FILLCELL_X1 FILLER_159_1511 ();
 FILLCELL_X2 FILLER_159_1533 ();
 FILLCELL_X8 FILLER_159_1541 ();
 FILLCELL_X1 FILLER_159_1549 ();
 FILLCELL_X32 FILLER_159_1555 ();
 FILLCELL_X32 FILLER_159_1587 ();
 FILLCELL_X32 FILLER_159_1619 ();
 FILLCELL_X16 FILLER_160_1 ();
 FILLCELL_X8 FILLER_160_17 ();
 FILLCELL_X4 FILLER_160_25 ();
 FILLCELL_X1 FILLER_160_29 ();
 FILLCELL_X2 FILLER_160_57 ();
 FILLCELL_X2 FILLER_160_72 ();
 FILLCELL_X1 FILLER_160_74 ();
 FILLCELL_X1 FILLER_160_86 ();
 FILLCELL_X8 FILLER_160_92 ();
 FILLCELL_X4 FILLER_160_100 ();
 FILLCELL_X1 FILLER_160_131 ();
 FILLCELL_X16 FILLER_160_152 ();
 FILLCELL_X1 FILLER_160_168 ();
 FILLCELL_X1 FILLER_160_181 ();
 FILLCELL_X8 FILLER_160_209 ();
 FILLCELL_X4 FILLER_160_217 ();
 FILLCELL_X2 FILLER_160_221 ();
 FILLCELL_X4 FILLER_160_257 ();
 FILLCELL_X1 FILLER_160_261 ();
 FILLCELL_X4 FILLER_160_269 ();
 FILLCELL_X2 FILLER_160_273 ();
 FILLCELL_X1 FILLER_160_275 ();
 FILLCELL_X1 FILLER_160_320 ();
 FILLCELL_X2 FILLER_160_344 ();
 FILLCELL_X4 FILLER_160_356 ();
 FILLCELL_X2 FILLER_160_367 ();
 FILLCELL_X4 FILLER_160_392 ();
 FILLCELL_X1 FILLER_160_396 ();
 FILLCELL_X1 FILLER_160_417 ();
 FILLCELL_X8 FILLER_160_421 ();
 FILLCELL_X4 FILLER_160_429 ();
 FILLCELL_X2 FILLER_160_457 ();
 FILLCELL_X1 FILLER_160_459 ();
 FILLCELL_X4 FILLER_160_471 ();
 FILLCELL_X4 FILLER_160_518 ();
 FILLCELL_X8 FILLER_160_611 ();
 FILLCELL_X1 FILLER_160_619 ();
 FILLCELL_X4 FILLER_160_627 ();
 FILLCELL_X4 FILLER_160_632 ();
 FILLCELL_X4 FILLER_160_656 ();
 FILLCELL_X1 FILLER_160_684 ();
 FILLCELL_X2 FILLER_160_701 ();
 FILLCELL_X4 FILLER_160_710 ();
 FILLCELL_X1 FILLER_160_734 ();
 FILLCELL_X1 FILLER_160_740 ();
 FILLCELL_X1 FILLER_160_765 ();
 FILLCELL_X4 FILLER_160_786 ();
 FILLCELL_X1 FILLER_160_790 ();
 FILLCELL_X2 FILLER_160_798 ();
 FILLCELL_X4 FILLER_160_804 ();
 FILLCELL_X1 FILLER_160_816 ();
 FILLCELL_X1 FILLER_160_820 ();
 FILLCELL_X4 FILLER_160_828 ();
 FILLCELL_X2 FILLER_160_832 ();
 FILLCELL_X2 FILLER_160_839 ();
 FILLCELL_X1 FILLER_160_841 ();
 FILLCELL_X4 FILLER_160_845 ();
 FILLCELL_X1 FILLER_160_849 ();
 FILLCELL_X2 FILLER_160_889 ();
 FILLCELL_X1 FILLER_160_891 ();
 FILLCELL_X4 FILLER_160_912 ();
 FILLCELL_X2 FILLER_160_916 ();
 FILLCELL_X8 FILLER_160_942 ();
 FILLCELL_X2 FILLER_160_950 ();
 FILLCELL_X1 FILLER_160_952 ();
 FILLCELL_X2 FILLER_160_1018 ();
 FILLCELL_X4 FILLER_160_1034 ();
 FILLCELL_X2 FILLER_160_1038 ();
 FILLCELL_X1 FILLER_160_1040 ();
 FILLCELL_X4 FILLER_160_1054 ();
 FILLCELL_X32 FILLER_160_1072 ();
 FILLCELL_X32 FILLER_160_1104 ();
 FILLCELL_X32 FILLER_160_1136 ();
 FILLCELL_X32 FILLER_160_1168 ();
 FILLCELL_X32 FILLER_160_1200 ();
 FILLCELL_X32 FILLER_160_1232 ();
 FILLCELL_X32 FILLER_160_1264 ();
 FILLCELL_X32 FILLER_160_1296 ();
 FILLCELL_X32 FILLER_160_1328 ();
 FILLCELL_X32 FILLER_160_1360 ();
 FILLCELL_X8 FILLER_160_1392 ();
 FILLCELL_X4 FILLER_160_1400 ();
 FILLCELL_X2 FILLER_160_1404 ();
 FILLCELL_X1 FILLER_160_1406 ();
 FILLCELL_X4 FILLER_160_1425 ();
 FILLCELL_X4 FILLER_160_1432 ();
 FILLCELL_X4 FILLER_160_1440 ();
 FILLCELL_X2 FILLER_160_1444 ();
 FILLCELL_X1 FILLER_160_1450 ();
 FILLCELL_X1 FILLER_160_1455 ();
 FILLCELL_X2 FILLER_160_1465 ();
 FILLCELL_X1 FILLER_160_1467 ();
 FILLCELL_X4 FILLER_160_1479 ();
 FILLCELL_X1 FILLER_160_1483 ();
 FILLCELL_X1 FILLER_160_1488 ();
 FILLCELL_X1 FILLER_160_1493 ();
 FILLCELL_X2 FILLER_160_1520 ();
 FILLCELL_X1 FILLER_160_1522 ();
 FILLCELL_X2 FILLER_160_1528 ();
 FILLCELL_X1 FILLER_160_1530 ();
 FILLCELL_X4 FILLER_160_1541 ();
 FILLCELL_X1 FILLER_160_1545 ();
 FILLCELL_X4 FILLER_160_1553 ();
 FILLCELL_X2 FILLER_160_1557 ();
 FILLCELL_X32 FILLER_160_1566 ();
 FILLCELL_X32 FILLER_160_1598 ();
 FILLCELL_X16 FILLER_160_1630 ();
 FILLCELL_X4 FILLER_160_1646 ();
 FILLCELL_X1 FILLER_160_1650 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X1 FILLER_161_33 ();
 FILLCELL_X8 FILLER_161_42 ();
 FILLCELL_X2 FILLER_161_50 ();
 FILLCELL_X1 FILLER_161_52 ();
 FILLCELL_X4 FILLER_161_60 ();
 FILLCELL_X16 FILLER_161_93 ();
 FILLCELL_X8 FILLER_161_109 ();
 FILLCELL_X4 FILLER_161_117 ();
 FILLCELL_X1 FILLER_161_121 ();
 FILLCELL_X4 FILLER_161_142 ();
 FILLCELL_X1 FILLER_161_146 ();
 FILLCELL_X2 FILLER_161_154 ();
 FILLCELL_X1 FILLER_161_156 ();
 FILLCELL_X1 FILLER_161_177 ();
 FILLCELL_X4 FILLER_161_198 ();
 FILLCELL_X2 FILLER_161_202 ();
 FILLCELL_X16 FILLER_161_211 ();
 FILLCELL_X2 FILLER_161_227 ();
 FILLCELL_X1 FILLER_161_229 ();
 FILLCELL_X4 FILLER_161_237 ();
 FILLCELL_X2 FILLER_161_241 ();
 FILLCELL_X1 FILLER_161_243 ();
 FILLCELL_X1 FILLER_161_247 ();
 FILLCELL_X2 FILLER_161_273 ();
 FILLCELL_X4 FILLER_161_282 ();
 FILLCELL_X1 FILLER_161_350 ();
 FILLCELL_X2 FILLER_161_380 ();
 FILLCELL_X2 FILLER_161_385 ();
 FILLCELL_X4 FILLER_161_395 ();
 FILLCELL_X1 FILLER_161_443 ();
 FILLCELL_X1 FILLER_161_451 ();
 FILLCELL_X8 FILLER_161_456 ();
 FILLCELL_X1 FILLER_161_464 ();
 FILLCELL_X1 FILLER_161_485 ();
 FILLCELL_X1 FILLER_161_490 ();
 FILLCELL_X1 FILLER_161_544 ();
 FILLCELL_X8 FILLER_161_585 ();
 FILLCELL_X1 FILLER_161_593 ();
 FILLCELL_X2 FILLER_161_601 ();
 FILLCELL_X1 FILLER_161_603 ();
 FILLCELL_X1 FILLER_161_615 ();
 FILLCELL_X1 FILLER_161_619 ();
 FILLCELL_X2 FILLER_161_652 ();
 FILLCELL_X1 FILLER_161_654 ();
 FILLCELL_X2 FILLER_161_698 ();
 FILLCELL_X1 FILLER_161_700 ();
 FILLCELL_X1 FILLER_161_721 ();
 FILLCELL_X4 FILLER_161_742 ();
 FILLCELL_X2 FILLER_161_746 ();
 FILLCELL_X1 FILLER_161_751 ();
 FILLCELL_X2 FILLER_161_784 ();
 FILLCELL_X8 FILLER_161_806 ();
 FILLCELL_X2 FILLER_161_814 ();
 FILLCELL_X8 FILLER_161_840 ();
 FILLCELL_X2 FILLER_161_848 ();
 FILLCELL_X1 FILLER_161_850 ();
 FILLCELL_X16 FILLER_161_862 ();
 FILLCELL_X2 FILLER_161_898 ();
 FILLCELL_X1 FILLER_161_900 ();
 FILLCELL_X4 FILLER_161_908 ();
 FILLCELL_X1 FILLER_161_912 ();
 FILLCELL_X1 FILLER_161_933 ();
 FILLCELL_X32 FILLER_161_961 ();
 FILLCELL_X4 FILLER_161_993 ();
 FILLCELL_X2 FILLER_161_997 ();
 FILLCELL_X8 FILLER_161_1002 ();
 FILLCELL_X4 FILLER_161_1010 ();
 FILLCELL_X2 FILLER_161_1014 ();
 FILLCELL_X1 FILLER_161_1036 ();
 FILLCELL_X2 FILLER_161_1044 ();
 FILLCELL_X2 FILLER_161_1082 ();
 FILLCELL_X1 FILLER_161_1084 ();
 FILLCELL_X32 FILLER_161_1105 ();
 FILLCELL_X32 FILLER_161_1137 ();
 FILLCELL_X32 FILLER_161_1169 ();
 FILLCELL_X32 FILLER_161_1201 ();
 FILLCELL_X16 FILLER_161_1233 ();
 FILLCELL_X8 FILLER_161_1249 ();
 FILLCELL_X4 FILLER_161_1257 ();
 FILLCELL_X2 FILLER_161_1261 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_161_1328 ();
 FILLCELL_X32 FILLER_161_1360 ();
 FILLCELL_X16 FILLER_161_1392 ();
 FILLCELL_X4 FILLER_161_1408 ();
 FILLCELL_X2 FILLER_161_1412 ();
 FILLCELL_X1 FILLER_161_1414 ();
 FILLCELL_X16 FILLER_161_1420 ();
 FILLCELL_X8 FILLER_161_1436 ();
 FILLCELL_X2 FILLER_161_1444 ();
 FILLCELL_X4 FILLER_161_1450 ();
 FILLCELL_X2 FILLER_161_1454 ();
 FILLCELL_X1 FILLER_161_1456 ();
 FILLCELL_X8 FILLER_161_1464 ();
 FILLCELL_X2 FILLER_161_1472 ();
 FILLCELL_X1 FILLER_161_1474 ();
 FILLCELL_X2 FILLER_161_1479 ();
 FILLCELL_X4 FILLER_161_1507 ();
 FILLCELL_X1 FILLER_161_1511 ();
 FILLCELL_X4 FILLER_161_1516 ();
 FILLCELL_X32 FILLER_161_1527 ();
 FILLCELL_X32 FILLER_161_1559 ();
 FILLCELL_X32 FILLER_161_1591 ();
 FILLCELL_X16 FILLER_161_1623 ();
 FILLCELL_X8 FILLER_161_1639 ();
 FILLCELL_X4 FILLER_161_1647 ();
 FILLCELL_X16 FILLER_162_1 ();
 FILLCELL_X8 FILLER_162_17 ();
 FILLCELL_X1 FILLER_162_25 ();
 FILLCELL_X8 FILLER_162_66 ();
 FILLCELL_X1 FILLER_162_74 ();
 FILLCELL_X4 FILLER_162_95 ();
 FILLCELL_X1 FILLER_162_99 ();
 FILLCELL_X16 FILLER_162_104 ();
 FILLCELL_X4 FILLER_162_120 ();
 FILLCELL_X2 FILLER_162_124 ();
 FILLCELL_X1 FILLER_162_126 ();
 FILLCELL_X1 FILLER_162_182 ();
 FILLCELL_X2 FILLER_162_223 ();
 FILLCELL_X1 FILLER_162_225 ();
 FILLCELL_X2 FILLER_162_239 ();
 FILLCELL_X2 FILLER_162_264 ();
 FILLCELL_X1 FILLER_162_266 ();
 FILLCELL_X16 FILLER_162_276 ();
 FILLCELL_X8 FILLER_162_292 ();
 FILLCELL_X4 FILLER_162_303 ();
 FILLCELL_X1 FILLER_162_307 ();
 FILLCELL_X4 FILLER_162_312 ();
 FILLCELL_X2 FILLER_162_316 ();
 FILLCELL_X1 FILLER_162_318 ();
 FILLCELL_X8 FILLER_162_322 ();
 FILLCELL_X4 FILLER_162_330 ();
 FILLCELL_X2 FILLER_162_334 ();
 FILLCELL_X1 FILLER_162_336 ();
 FILLCELL_X2 FILLER_162_345 ();
 FILLCELL_X1 FILLER_162_350 ();
 FILLCELL_X8 FILLER_162_360 ();
 FILLCELL_X4 FILLER_162_368 ();
 FILLCELL_X1 FILLER_162_392 ();
 FILLCELL_X4 FILLER_162_396 ();
 FILLCELL_X1 FILLER_162_400 ();
 FILLCELL_X8 FILLER_162_421 ();
 FILLCELL_X2 FILLER_162_429 ();
 FILLCELL_X1 FILLER_162_431 ();
 FILLCELL_X16 FILLER_162_452 ();
 FILLCELL_X2 FILLER_162_468 ();
 FILLCELL_X1 FILLER_162_482 ();
 FILLCELL_X1 FILLER_162_503 ();
 FILLCELL_X2 FILLER_162_512 ();
 FILLCELL_X1 FILLER_162_514 ();
 FILLCELL_X8 FILLER_162_538 ();
 FILLCELL_X2 FILLER_162_546 ();
 FILLCELL_X1 FILLER_162_548 ();
 FILLCELL_X2 FILLER_162_564 ();
 FILLCELL_X16 FILLER_162_580 ();
 FILLCELL_X8 FILLER_162_596 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X4 FILLER_162_632 ();
 FILLCELL_X1 FILLER_162_639 ();
 FILLCELL_X2 FILLER_162_651 ();
 FILLCELL_X1 FILLER_162_653 ();
 FILLCELL_X4 FILLER_162_659 ();
 FILLCELL_X2 FILLER_162_663 ();
 FILLCELL_X1 FILLER_162_665 ();
 FILLCELL_X8 FILLER_162_669 ();
 FILLCELL_X1 FILLER_162_677 ();
 FILLCELL_X4 FILLER_162_685 ();
 FILLCELL_X2 FILLER_162_693 ();
 FILLCELL_X1 FILLER_162_695 ();
 FILLCELL_X8 FILLER_162_701 ();
 FILLCELL_X4 FILLER_162_709 ();
 FILLCELL_X1 FILLER_162_713 ();
 FILLCELL_X4 FILLER_162_741 ();
 FILLCELL_X1 FILLER_162_745 ();
 FILLCELL_X1 FILLER_162_766 ();
 FILLCELL_X2 FILLER_162_771 ();
 FILLCELL_X8 FILLER_162_785 ();
 FILLCELL_X4 FILLER_162_793 ();
 FILLCELL_X2 FILLER_162_801 ();
 FILLCELL_X8 FILLER_162_806 ();
 FILLCELL_X4 FILLER_162_814 ();
 FILLCELL_X1 FILLER_162_818 ();
 FILLCELL_X8 FILLER_162_824 ();
 FILLCELL_X8 FILLER_162_834 ();
 FILLCELL_X4 FILLER_162_842 ();
 FILLCELL_X2 FILLER_162_846 ();
 FILLCELL_X1 FILLER_162_848 ();
 FILLCELL_X2 FILLER_162_871 ();
 FILLCELL_X1 FILLER_162_873 ();
 FILLCELL_X8 FILLER_162_905 ();
 FILLCELL_X4 FILLER_162_913 ();
 FILLCELL_X4 FILLER_162_924 ();
 FILLCELL_X4 FILLER_162_931 ();
 FILLCELL_X2 FILLER_162_935 ();
 FILLCELL_X1 FILLER_162_937 ();
 FILLCELL_X2 FILLER_162_965 ();
 FILLCELL_X1 FILLER_162_997 ();
 FILLCELL_X4 FILLER_162_1044 ();
 FILLCELL_X8 FILLER_162_1073 ();
 FILLCELL_X4 FILLER_162_1081 ();
 FILLCELL_X1 FILLER_162_1085 ();
 FILLCELL_X4 FILLER_162_1096 ();
 FILLCELL_X32 FILLER_162_1110 ();
 FILLCELL_X32 FILLER_162_1142 ();
 FILLCELL_X1 FILLER_162_1174 ();
 FILLCELL_X32 FILLER_162_1195 ();
 FILLCELL_X32 FILLER_162_1227 ();
 FILLCELL_X32 FILLER_162_1259 ();
 FILLCELL_X32 FILLER_162_1291 ();
 FILLCELL_X32 FILLER_162_1323 ();
 FILLCELL_X32 FILLER_162_1355 ();
 FILLCELL_X32 FILLER_162_1387 ();
 FILLCELL_X32 FILLER_162_1419 ();
 FILLCELL_X32 FILLER_162_1451 ();
 FILLCELL_X32 FILLER_162_1483 ();
 FILLCELL_X32 FILLER_162_1515 ();
 FILLCELL_X32 FILLER_162_1547 ();
 FILLCELL_X32 FILLER_162_1579 ();
 FILLCELL_X32 FILLER_162_1611 ();
 FILLCELL_X8 FILLER_162_1643 ();
 FILLCELL_X16 FILLER_163_1 ();
 FILLCELL_X4 FILLER_163_17 ();
 FILLCELL_X2 FILLER_163_21 ();
 FILLCELL_X1 FILLER_163_23 ();
 FILLCELL_X4 FILLER_163_71 ();
 FILLCELL_X2 FILLER_163_75 ();
 FILLCELL_X1 FILLER_163_82 ();
 FILLCELL_X1 FILLER_163_127 ();
 FILLCELL_X1 FILLER_163_138 ();
 FILLCELL_X4 FILLER_163_196 ();
 FILLCELL_X2 FILLER_163_200 ();
 FILLCELL_X2 FILLER_163_242 ();
 FILLCELL_X8 FILLER_163_251 ();
 FILLCELL_X2 FILLER_163_259 ();
 FILLCELL_X4 FILLER_163_268 ();
 FILLCELL_X1 FILLER_163_272 ();
 FILLCELL_X2 FILLER_163_287 ();
 FILLCELL_X1 FILLER_163_289 ();
 FILLCELL_X2 FILLER_163_294 ();
 FILLCELL_X1 FILLER_163_296 ();
 FILLCELL_X2 FILLER_163_300 ();
 FILLCELL_X1 FILLER_163_302 ();
 FILLCELL_X2 FILLER_163_355 ();
 FILLCELL_X8 FILLER_163_384 ();
 FILLCELL_X4 FILLER_163_392 ();
 FILLCELL_X2 FILLER_163_396 ();
 FILLCELL_X8 FILLER_163_421 ();
 FILLCELL_X2 FILLER_163_449 ();
 FILLCELL_X8 FILLER_163_455 ();
 FILLCELL_X2 FILLER_163_463 ();
 FILLCELL_X1 FILLER_163_465 ();
 FILLCELL_X1 FILLER_163_495 ();
 FILLCELL_X2 FILLER_163_500 ();
 FILLCELL_X1 FILLER_163_502 ();
 FILLCELL_X8 FILLER_163_506 ();
 FILLCELL_X2 FILLER_163_514 ();
 FILLCELL_X1 FILLER_163_516 ();
 FILLCELL_X8 FILLER_163_546 ();
 FILLCELL_X1 FILLER_163_554 ();
 FILLCELL_X8 FILLER_163_583 ();
 FILLCELL_X4 FILLER_163_591 ();
 FILLCELL_X1 FILLER_163_595 ();
 FILLCELL_X8 FILLER_163_616 ();
 FILLCELL_X4 FILLER_163_624 ();
 FILLCELL_X2 FILLER_163_628 ();
 FILLCELL_X1 FILLER_163_630 ();
 FILLCELL_X1 FILLER_163_635 ();
 FILLCELL_X1 FILLER_163_656 ();
 FILLCELL_X1 FILLER_163_660 ();
 FILLCELL_X4 FILLER_163_696 ();
 FILLCELL_X2 FILLER_163_700 ();
 FILLCELL_X1 FILLER_163_702 ();
 FILLCELL_X8 FILLER_163_710 ();
 FILLCELL_X2 FILLER_163_743 ();
 FILLCELL_X1 FILLER_163_745 ();
 FILLCELL_X4 FILLER_163_765 ();
 FILLCELL_X2 FILLER_163_769 ();
 FILLCELL_X4 FILLER_163_778 ();
 FILLCELL_X2 FILLER_163_816 ();
 FILLCELL_X8 FILLER_163_838 ();
 FILLCELL_X2 FILLER_163_878 ();
 FILLCELL_X4 FILLER_163_907 ();
 FILLCELL_X1 FILLER_163_911 ();
 FILLCELL_X4 FILLER_163_925 ();
 FILLCELL_X4 FILLER_163_936 ();
 FILLCELL_X8 FILLER_163_947 ();
 FILLCELL_X4 FILLER_163_955 ();
 FILLCELL_X2 FILLER_163_959 ();
 FILLCELL_X1 FILLER_163_961 ();
 FILLCELL_X1 FILLER_163_979 ();
 FILLCELL_X1 FILLER_163_984 ();
 FILLCELL_X1 FILLER_163_1003 ();
 FILLCELL_X4 FILLER_163_1007 ();
 FILLCELL_X2 FILLER_163_1018 ();
 FILLCELL_X8 FILLER_163_1040 ();
 FILLCELL_X1 FILLER_163_1048 ();
 FILLCELL_X16 FILLER_163_1066 ();
 FILLCELL_X2 FILLER_163_1082 ();
 FILLCELL_X1 FILLER_163_1084 ();
 FILLCELL_X32 FILLER_163_1112 ();
 FILLCELL_X32 FILLER_163_1144 ();
 FILLCELL_X8 FILLER_163_1176 ();
 FILLCELL_X2 FILLER_163_1184 ();
 FILLCELL_X1 FILLER_163_1186 ();
 FILLCELL_X32 FILLER_163_1191 ();
 FILLCELL_X32 FILLER_163_1223 ();
 FILLCELL_X8 FILLER_163_1255 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X32 FILLER_163_1296 ();
 FILLCELL_X32 FILLER_163_1328 ();
 FILLCELL_X32 FILLER_163_1360 ();
 FILLCELL_X32 FILLER_163_1392 ();
 FILLCELL_X32 FILLER_163_1424 ();
 FILLCELL_X32 FILLER_163_1456 ();
 FILLCELL_X32 FILLER_163_1488 ();
 FILLCELL_X32 FILLER_163_1520 ();
 FILLCELL_X32 FILLER_163_1552 ();
 FILLCELL_X32 FILLER_163_1584 ();
 FILLCELL_X32 FILLER_163_1616 ();
 FILLCELL_X2 FILLER_163_1648 ();
 FILLCELL_X1 FILLER_163_1650 ();
 FILLCELL_X16 FILLER_164_1 ();
 FILLCELL_X8 FILLER_164_17 ();
 FILLCELL_X4 FILLER_164_25 ();
 FILLCELL_X1 FILLER_164_36 ();
 FILLCELL_X8 FILLER_164_44 ();
 FILLCELL_X2 FILLER_164_52 ();
 FILLCELL_X1 FILLER_164_54 ();
 FILLCELL_X2 FILLER_164_75 ();
 FILLCELL_X1 FILLER_164_77 ();
 FILLCELL_X2 FILLER_164_85 ();
 FILLCELL_X1 FILLER_164_97 ();
 FILLCELL_X2 FILLER_164_125 ();
 FILLCELL_X1 FILLER_164_127 ();
 FILLCELL_X2 FILLER_164_152 ();
 FILLCELL_X16 FILLER_164_194 ();
 FILLCELL_X8 FILLER_164_210 ();
 FILLCELL_X2 FILLER_164_218 ();
 FILLCELL_X1 FILLER_164_220 ();
 FILLCELL_X1 FILLER_164_241 ();
 FILLCELL_X1 FILLER_164_246 ();
 FILLCELL_X1 FILLER_164_250 ();
 FILLCELL_X2 FILLER_164_255 ();
 FILLCELL_X4 FILLER_164_260 ();
 FILLCELL_X4 FILLER_164_309 ();
 FILLCELL_X2 FILLER_164_313 ();
 FILLCELL_X1 FILLER_164_340 ();
 FILLCELL_X2 FILLER_164_355 ();
 FILLCELL_X4 FILLER_164_364 ();
 FILLCELL_X1 FILLER_164_368 ();
 FILLCELL_X4 FILLER_164_393 ();
 FILLCELL_X1 FILLER_164_397 ();
 FILLCELL_X2 FILLER_164_443 ();
 FILLCELL_X2 FILLER_164_472 ();
 FILLCELL_X1 FILLER_164_474 ();
 FILLCELL_X4 FILLER_164_478 ();
 FILLCELL_X4 FILLER_164_484 ();
 FILLCELL_X8 FILLER_164_513 ();
 FILLCELL_X4 FILLER_164_521 ();
 FILLCELL_X2 FILLER_164_525 ();
 FILLCELL_X2 FILLER_164_531 ();
 FILLCELL_X2 FILLER_164_536 ();
 FILLCELL_X2 FILLER_164_542 ();
 FILLCELL_X1 FILLER_164_544 ();
 FILLCELL_X2 FILLER_164_562 ();
 FILLCELL_X1 FILLER_164_567 ();
 FILLCELL_X4 FILLER_164_577 ();
 FILLCELL_X8 FILLER_164_584 ();
 FILLCELL_X2 FILLER_164_592 ();
 FILLCELL_X2 FILLER_164_598 ();
 FILLCELL_X1 FILLER_164_600 ();
 FILLCELL_X1 FILLER_164_605 ();
 FILLCELL_X4 FILLER_164_609 ();
 FILLCELL_X8 FILLER_164_620 ();
 FILLCELL_X2 FILLER_164_628 ();
 FILLCELL_X1 FILLER_164_630 ();
 FILLCELL_X4 FILLER_164_636 ();
 FILLCELL_X2 FILLER_164_640 ();
 FILLCELL_X1 FILLER_164_642 ();
 FILLCELL_X8 FILLER_164_650 ();
 FILLCELL_X2 FILLER_164_749 ();
 FILLCELL_X1 FILLER_164_751 ();
 FILLCELL_X2 FILLER_164_792 ();
 FILLCELL_X1 FILLER_164_794 ();
 FILLCELL_X4 FILLER_164_802 ();
 FILLCELL_X2 FILLER_164_806 ();
 FILLCELL_X4 FILLER_164_828 ();
 FILLCELL_X2 FILLER_164_832 ();
 FILLCELL_X8 FILLER_164_847 ();
 FILLCELL_X1 FILLER_164_858 ();
 FILLCELL_X4 FILLER_164_866 ();
 FILLCELL_X1 FILLER_164_900 ();
 FILLCELL_X8 FILLER_164_925 ();
 FILLCELL_X1 FILLER_164_933 ();
 FILLCELL_X1 FILLER_164_994 ();
 FILLCELL_X1 FILLER_164_1026 ();
 FILLCELL_X16 FILLER_164_1054 ();
 FILLCELL_X4 FILLER_164_1070 ();
 FILLCELL_X2 FILLER_164_1074 ();
 FILLCELL_X1 FILLER_164_1076 ();
 FILLCELL_X8 FILLER_164_1082 ();
 FILLCELL_X2 FILLER_164_1095 ();
 FILLCELL_X1 FILLER_164_1097 ();
 FILLCELL_X16 FILLER_164_1105 ();
 FILLCELL_X32 FILLER_164_1131 ();
 FILLCELL_X32 FILLER_164_1163 ();
 FILLCELL_X32 FILLER_164_1195 ();
 FILLCELL_X32 FILLER_164_1227 ();
 FILLCELL_X32 FILLER_164_1259 ();
 FILLCELL_X32 FILLER_164_1291 ();
 FILLCELL_X32 FILLER_164_1323 ();
 FILLCELL_X32 FILLER_164_1355 ();
 FILLCELL_X32 FILLER_164_1387 ();
 FILLCELL_X32 FILLER_164_1419 ();
 FILLCELL_X32 FILLER_164_1451 ();
 FILLCELL_X32 FILLER_164_1483 ();
 FILLCELL_X32 FILLER_164_1515 ();
 FILLCELL_X32 FILLER_164_1547 ();
 FILLCELL_X32 FILLER_164_1579 ();
 FILLCELL_X32 FILLER_164_1611 ();
 FILLCELL_X8 FILLER_164_1643 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X8 FILLER_165_33 ();
 FILLCELL_X2 FILLER_165_41 ();
 FILLCELL_X1 FILLER_165_43 ();
 FILLCELL_X2 FILLER_165_57 ();
 FILLCELL_X2 FILLER_165_66 ();
 FILLCELL_X1 FILLER_165_68 ();
 FILLCELL_X2 FILLER_165_89 ();
 FILLCELL_X1 FILLER_165_91 ();
 FILLCELL_X2 FILLER_165_99 ();
 FILLCELL_X16 FILLER_165_138 ();
 FILLCELL_X2 FILLER_165_154 ();
 FILLCELL_X1 FILLER_165_156 ();
 FILLCELL_X4 FILLER_165_166 ();
 FILLCELL_X1 FILLER_165_170 ();
 FILLCELL_X1 FILLER_165_178 ();
 FILLCELL_X2 FILLER_165_186 ();
 FILLCELL_X8 FILLER_165_192 ();
 FILLCELL_X4 FILLER_165_200 ();
 FILLCELL_X2 FILLER_165_204 ();
 FILLCELL_X1 FILLER_165_206 ();
 FILLCELL_X8 FILLER_165_214 ();
 FILLCELL_X4 FILLER_165_222 ();
 FILLCELL_X2 FILLER_165_307 ();
 FILLCELL_X1 FILLER_165_317 ();
 FILLCELL_X2 FILLER_165_327 ();
 FILLCELL_X2 FILLER_165_335 ();
 FILLCELL_X1 FILLER_165_337 ();
 FILLCELL_X16 FILLER_165_358 ();
 FILLCELL_X4 FILLER_165_377 ();
 FILLCELL_X4 FILLER_165_401 ();
 FILLCELL_X2 FILLER_165_405 ();
 FILLCELL_X1 FILLER_165_407 ();
 FILLCELL_X1 FILLER_165_413 ();
 FILLCELL_X8 FILLER_165_437 ();
 FILLCELL_X2 FILLER_165_445 ();
 FILLCELL_X1 FILLER_165_487 ();
 FILLCELL_X2 FILLER_165_545 ();
 FILLCELL_X4 FILLER_165_567 ();
 FILLCELL_X1 FILLER_165_571 ();
 FILLCELL_X2 FILLER_165_577 ();
 FILLCELL_X1 FILLER_165_583 ();
 FILLCELL_X2 FILLER_165_589 ();
 FILLCELL_X16 FILLER_165_654 ();
 FILLCELL_X1 FILLER_165_670 ();
 FILLCELL_X8 FILLER_165_674 ();
 FILLCELL_X1 FILLER_165_682 ();
 FILLCELL_X2 FILLER_165_687 ();
 FILLCELL_X4 FILLER_165_692 ();
 FILLCELL_X2 FILLER_165_696 ();
 FILLCELL_X16 FILLER_165_717 ();
 FILLCELL_X2 FILLER_165_740 ();
 FILLCELL_X1 FILLER_165_742 ();
 FILLCELL_X2 FILLER_165_748 ();
 FILLCELL_X8 FILLER_165_759 ();
 FILLCELL_X2 FILLER_165_767 ();
 FILLCELL_X2 FILLER_165_796 ();
 FILLCELL_X1 FILLER_165_798 ();
 FILLCELL_X32 FILLER_165_819 ();
 FILLCELL_X1 FILLER_165_851 ();
 FILLCELL_X16 FILLER_165_872 ();
 FILLCELL_X4 FILLER_165_888 ();
 FILLCELL_X1 FILLER_165_892 ();
 FILLCELL_X4 FILLER_165_900 ();
 FILLCELL_X2 FILLER_165_921 ();
 FILLCELL_X1 FILLER_165_923 ();
 FILLCELL_X16 FILLER_165_937 ();
 FILLCELL_X8 FILLER_165_953 ();
 FILLCELL_X2 FILLER_165_961 ();
 FILLCELL_X16 FILLER_165_986 ();
 FILLCELL_X1 FILLER_165_1002 ();
 FILLCELL_X2 FILLER_165_1008 ();
 FILLCELL_X1 FILLER_165_1012 ();
 FILLCELL_X4 FILLER_165_1043 ();
 FILLCELL_X1 FILLER_165_1047 ();
 FILLCELL_X8 FILLER_165_1071 ();
 FILLCELL_X4 FILLER_165_1079 ();
 FILLCELL_X1 FILLER_165_1083 ();
 FILLCELL_X32 FILLER_165_1093 ();
 FILLCELL_X32 FILLER_165_1125 ();
 FILLCELL_X32 FILLER_165_1157 ();
 FILLCELL_X32 FILLER_165_1189 ();
 FILLCELL_X32 FILLER_165_1221 ();
 FILLCELL_X8 FILLER_165_1253 ();
 FILLCELL_X2 FILLER_165_1261 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_165_1328 ();
 FILLCELL_X32 FILLER_165_1360 ();
 FILLCELL_X32 FILLER_165_1392 ();
 FILLCELL_X32 FILLER_165_1424 ();
 FILLCELL_X32 FILLER_165_1456 ();
 FILLCELL_X32 FILLER_165_1488 ();
 FILLCELL_X32 FILLER_165_1520 ();
 FILLCELL_X32 FILLER_165_1552 ();
 FILLCELL_X32 FILLER_165_1584 ();
 FILLCELL_X32 FILLER_165_1616 ();
 FILLCELL_X2 FILLER_165_1648 ();
 FILLCELL_X1 FILLER_165_1650 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X16 FILLER_166_33 ();
 FILLCELL_X8 FILLER_166_49 ();
 FILLCELL_X2 FILLER_166_57 ();
 FILLCELL_X4 FILLER_166_86 ();
 FILLCELL_X2 FILLER_166_90 ();
 FILLCELL_X1 FILLER_166_92 ();
 FILLCELL_X8 FILLER_166_147 ();
 FILLCELL_X1 FILLER_166_155 ();
 FILLCELL_X4 FILLER_166_173 ();
 FILLCELL_X2 FILLER_166_177 ();
 FILLCELL_X8 FILLER_166_226 ();
 FILLCELL_X2 FILLER_166_234 ();
 FILLCELL_X1 FILLER_166_236 ();
 FILLCELL_X1 FILLER_166_257 ();
 FILLCELL_X4 FILLER_166_285 ();
 FILLCELL_X2 FILLER_166_289 ();
 FILLCELL_X2 FILLER_166_315 ();
 FILLCELL_X4 FILLER_166_342 ();
 FILLCELL_X16 FILLER_166_351 ();
 FILLCELL_X4 FILLER_166_367 ();
 FILLCELL_X1 FILLER_166_371 ();
 FILLCELL_X2 FILLER_166_377 ();
 FILLCELL_X4 FILLER_166_381 ();
 FILLCELL_X1 FILLER_166_385 ();
 FILLCELL_X8 FILLER_166_390 ();
 FILLCELL_X2 FILLER_166_405 ();
 FILLCELL_X4 FILLER_166_415 ();
 FILLCELL_X1 FILLER_166_423 ();
 FILLCELL_X4 FILLER_166_444 ();
 FILLCELL_X2 FILLER_166_448 ();
 FILLCELL_X1 FILLER_166_450 ();
 FILLCELL_X1 FILLER_166_458 ();
 FILLCELL_X16 FILLER_166_476 ();
 FILLCELL_X4 FILLER_166_492 ();
 FILLCELL_X1 FILLER_166_496 ();
 FILLCELL_X4 FILLER_166_504 ();
 FILLCELL_X1 FILLER_166_508 ();
 FILLCELL_X4 FILLER_166_533 ();
 FILLCELL_X2 FILLER_166_537 ();
 FILLCELL_X8 FILLER_166_544 ();
 FILLCELL_X2 FILLER_166_601 ();
 FILLCELL_X1 FILLER_166_603 ();
 FILLCELL_X1 FILLER_166_611 ();
 FILLCELL_X16 FILLER_166_615 ();
 FILLCELL_X1 FILLER_166_632 ();
 FILLCELL_X2 FILLER_166_699 ();
 FILLCELL_X1 FILLER_166_701 ();
 FILLCELL_X4 FILLER_166_722 ();
 FILLCELL_X1 FILLER_166_726 ();
 FILLCELL_X2 FILLER_166_747 ();
 FILLCELL_X4 FILLER_166_753 ();
 FILLCELL_X1 FILLER_166_757 ();
 FILLCELL_X8 FILLER_166_763 ();
 FILLCELL_X2 FILLER_166_771 ();
 FILLCELL_X8 FILLER_166_792 ();
 FILLCELL_X4 FILLER_166_800 ();
 FILLCELL_X1 FILLER_166_804 ();
 FILLCELL_X4 FILLER_166_845 ();
 FILLCELL_X1 FILLER_166_849 ();
 FILLCELL_X2 FILLER_166_855 ();
 FILLCELL_X8 FILLER_166_904 ();
 FILLCELL_X2 FILLER_166_912 ();
 FILLCELL_X1 FILLER_166_914 ();
 FILLCELL_X2 FILLER_166_923 ();
 FILLCELL_X1 FILLER_166_925 ();
 FILLCELL_X16 FILLER_166_933 ();
 FILLCELL_X2 FILLER_166_949 ();
 FILLCELL_X2 FILLER_166_964 ();
 FILLCELL_X1 FILLER_166_966 ();
 FILLCELL_X8 FILLER_166_972 ();
 FILLCELL_X1 FILLER_166_984 ();
 FILLCELL_X2 FILLER_166_1005 ();
 FILLCELL_X2 FILLER_166_1039 ();
 FILLCELL_X1 FILLER_166_1041 ();
 FILLCELL_X8 FILLER_166_1073 ();
 FILLCELL_X2 FILLER_166_1081 ();
 FILLCELL_X32 FILLER_166_1103 ();
 FILLCELL_X32 FILLER_166_1135 ();
 FILLCELL_X32 FILLER_166_1167 ();
 FILLCELL_X32 FILLER_166_1199 ();
 FILLCELL_X32 FILLER_166_1231 ();
 FILLCELL_X32 FILLER_166_1263 ();
 FILLCELL_X32 FILLER_166_1295 ();
 FILLCELL_X32 FILLER_166_1327 ();
 FILLCELL_X32 FILLER_166_1359 ();
 FILLCELL_X32 FILLER_166_1391 ();
 FILLCELL_X32 FILLER_166_1423 ();
 FILLCELL_X32 FILLER_166_1455 ();
 FILLCELL_X32 FILLER_166_1487 ();
 FILLCELL_X32 FILLER_166_1519 ();
 FILLCELL_X32 FILLER_166_1551 ();
 FILLCELL_X32 FILLER_166_1583 ();
 FILLCELL_X32 FILLER_166_1615 ();
 FILLCELL_X4 FILLER_166_1647 ();
 FILLCELL_X16 FILLER_167_1 ();
 FILLCELL_X8 FILLER_167_17 ();
 FILLCELL_X32 FILLER_167_45 ();
 FILLCELL_X16 FILLER_167_77 ();
 FILLCELL_X2 FILLER_167_93 ();
 FILLCELL_X1 FILLER_167_95 ();
 FILLCELL_X16 FILLER_167_109 ();
 FILLCELL_X4 FILLER_167_125 ();
 FILLCELL_X2 FILLER_167_129 ();
 FILLCELL_X2 FILLER_167_153 ();
 FILLCELL_X1 FILLER_167_180 ();
 FILLCELL_X2 FILLER_167_224 ();
 FILLCELL_X8 FILLER_167_235 ();
 FILLCELL_X1 FILLER_167_250 ();
 FILLCELL_X4 FILLER_167_264 ();
 FILLCELL_X2 FILLER_167_268 ();
 FILLCELL_X1 FILLER_167_270 ();
 FILLCELL_X1 FILLER_167_291 ();
 FILLCELL_X1 FILLER_167_299 ();
 FILLCELL_X1 FILLER_167_305 ();
 FILLCELL_X8 FILLER_167_311 ();
 FILLCELL_X4 FILLER_167_322 ();
 FILLCELL_X1 FILLER_167_326 ();
 FILLCELL_X8 FILLER_167_351 ();
 FILLCELL_X2 FILLER_167_359 ();
 FILLCELL_X1 FILLER_167_361 ();
 FILLCELL_X8 FILLER_167_382 ();
 FILLCELL_X1 FILLER_167_390 ();
 FILLCELL_X1 FILLER_167_411 ();
 FILLCELL_X1 FILLER_167_434 ();
 FILLCELL_X8 FILLER_167_438 ();
 FILLCELL_X4 FILLER_167_446 ();
 FILLCELL_X2 FILLER_167_450 ();
 FILLCELL_X1 FILLER_167_452 ();
 FILLCELL_X4 FILLER_167_457 ();
 FILLCELL_X1 FILLER_167_461 ();
 FILLCELL_X2 FILLER_167_465 ();
 FILLCELL_X4 FILLER_167_490 ();
 FILLCELL_X16 FILLER_167_501 ();
 FILLCELL_X2 FILLER_167_517 ();
 FILLCELL_X2 FILLER_167_531 ();
 FILLCELL_X4 FILLER_167_596 ();
 FILLCELL_X2 FILLER_167_600 ();
 FILLCELL_X2 FILLER_167_671 ();
 FILLCELL_X2 FILLER_167_677 ();
 FILLCELL_X1 FILLER_167_679 ();
 FILLCELL_X8 FILLER_167_683 ();
 FILLCELL_X4 FILLER_167_691 ();
 FILLCELL_X2 FILLER_167_695 ();
 FILLCELL_X2 FILLER_167_716 ();
 FILLCELL_X1 FILLER_167_718 ();
 FILLCELL_X16 FILLER_167_739 ();
 FILLCELL_X1 FILLER_167_755 ();
 FILLCELL_X8 FILLER_167_776 ();
 FILLCELL_X4 FILLER_167_784 ();
 FILLCELL_X2 FILLER_167_788 ();
 FILLCELL_X1 FILLER_167_790 ();
 FILLCELL_X8 FILLER_167_818 ();
 FILLCELL_X2 FILLER_167_826 ();
 FILLCELL_X1 FILLER_167_828 ();
 FILLCELL_X8 FILLER_167_884 ();
 FILLCELL_X2 FILLER_167_892 ();
 FILLCELL_X1 FILLER_167_894 ();
 FILLCELL_X8 FILLER_167_899 ();
 FILLCELL_X4 FILLER_167_907 ();
 FILLCELL_X1 FILLER_167_911 ();
 FILLCELL_X1 FILLER_167_990 ();
 FILLCELL_X16 FILLER_167_994 ();
 FILLCELL_X4 FILLER_167_1010 ();
 FILLCELL_X2 FILLER_167_1014 ();
 FILLCELL_X1 FILLER_167_1030 ();
 FILLCELL_X2 FILLER_167_1056 ();
 FILLCELL_X1 FILLER_167_1058 ();
 FILLCELL_X8 FILLER_167_1066 ();
 FILLCELL_X8 FILLER_167_1077 ();
 FILLCELL_X4 FILLER_167_1085 ();
 FILLCELL_X1 FILLER_167_1089 ();
 FILLCELL_X32 FILLER_167_1097 ();
 FILLCELL_X32 FILLER_167_1129 ();
 FILLCELL_X32 FILLER_167_1161 ();
 FILLCELL_X32 FILLER_167_1193 ();
 FILLCELL_X32 FILLER_167_1225 ();
 FILLCELL_X4 FILLER_167_1257 ();
 FILLCELL_X2 FILLER_167_1261 ();
 FILLCELL_X32 FILLER_167_1264 ();
 FILLCELL_X32 FILLER_167_1296 ();
 FILLCELL_X32 FILLER_167_1328 ();
 FILLCELL_X32 FILLER_167_1360 ();
 FILLCELL_X32 FILLER_167_1392 ();
 FILLCELL_X32 FILLER_167_1424 ();
 FILLCELL_X32 FILLER_167_1456 ();
 FILLCELL_X32 FILLER_167_1488 ();
 FILLCELL_X32 FILLER_167_1520 ();
 FILLCELL_X32 FILLER_167_1552 ();
 FILLCELL_X32 FILLER_167_1584 ();
 FILLCELL_X32 FILLER_167_1616 ();
 FILLCELL_X2 FILLER_167_1648 ();
 FILLCELL_X1 FILLER_167_1650 ();
 FILLCELL_X16 FILLER_168_1 ();
 FILLCELL_X8 FILLER_168_17 ();
 FILLCELL_X4 FILLER_168_25 ();
 FILLCELL_X2 FILLER_168_56 ();
 FILLCELL_X4 FILLER_168_83 ();
 FILLCELL_X8 FILLER_168_105 ();
 FILLCELL_X4 FILLER_168_113 ();
 FILLCELL_X2 FILLER_168_117 ();
 FILLCELL_X2 FILLER_168_132 ();
 FILLCELL_X2 FILLER_168_141 ();
 FILLCELL_X1 FILLER_168_143 ();
 FILLCELL_X2 FILLER_168_164 ();
 FILLCELL_X1 FILLER_168_166 ();
 FILLCELL_X2 FILLER_168_180 ();
 FILLCELL_X1 FILLER_168_189 ();
 FILLCELL_X4 FILLER_168_202 ();
 FILLCELL_X2 FILLER_168_206 ();
 FILLCELL_X1 FILLER_168_208 ();
 FILLCELL_X4 FILLER_168_254 ();
 FILLCELL_X1 FILLER_168_258 ();
 FILLCELL_X1 FILLER_168_286 ();
 FILLCELL_X1 FILLER_168_307 ();
 FILLCELL_X1 FILLER_168_332 ();
 FILLCELL_X8 FILLER_168_343 ();
 FILLCELL_X2 FILLER_168_351 ();
 FILLCELL_X1 FILLER_168_353 ();
 FILLCELL_X2 FILLER_168_377 ();
 FILLCELL_X2 FILLER_168_384 ();
 FILLCELL_X1 FILLER_168_386 ();
 FILLCELL_X1 FILLER_168_404 ();
 FILLCELL_X2 FILLER_168_448 ();
 FILLCELL_X1 FILLER_168_450 ();
 FILLCELL_X1 FILLER_168_522 ();
 FILLCELL_X4 FILLER_168_548 ();
 FILLCELL_X4 FILLER_168_556 ();
 FILLCELL_X2 FILLER_168_560 ();
 FILLCELL_X1 FILLER_168_562 ();
 FILLCELL_X4 FILLER_168_567 ();
 FILLCELL_X1 FILLER_168_574 ();
 FILLCELL_X16 FILLER_168_583 ();
 FILLCELL_X1 FILLER_168_606 ();
 FILLCELL_X2 FILLER_168_615 ();
 FILLCELL_X4 FILLER_168_632 ();
 FILLCELL_X2 FILLER_168_636 ();
 FILLCELL_X1 FILLER_168_638 ();
 FILLCELL_X4 FILLER_168_642 ();
 FILLCELL_X2 FILLER_168_655 ();
 FILLCELL_X4 FILLER_168_684 ();
 FILLCELL_X1 FILLER_168_688 ();
 FILLCELL_X8 FILLER_168_721 ();
 FILLCELL_X2 FILLER_168_729 ();
 FILLCELL_X16 FILLER_168_754 ();
 FILLCELL_X4 FILLER_168_770 ();
 FILLCELL_X2 FILLER_168_774 ();
 FILLCELL_X2 FILLER_168_796 ();
 FILLCELL_X2 FILLER_168_822 ();
 FILLCELL_X2 FILLER_168_831 ();
 FILLCELL_X1 FILLER_168_833 ();
 FILLCELL_X4 FILLER_168_841 ();
 FILLCELL_X1 FILLER_168_845 ();
 FILLCELL_X2 FILLER_168_853 ();
 FILLCELL_X4 FILLER_168_878 ();
 FILLCELL_X1 FILLER_168_882 ();
 FILLCELL_X1 FILLER_168_900 ();
 FILLCELL_X16 FILLER_168_943 ();
 FILLCELL_X2 FILLER_168_959 ();
 FILLCELL_X1 FILLER_168_961 ();
 FILLCELL_X4 FILLER_168_1045 ();
 FILLCELL_X8 FILLER_168_1055 ();
 FILLCELL_X32 FILLER_168_1090 ();
 FILLCELL_X32 FILLER_168_1122 ();
 FILLCELL_X32 FILLER_168_1154 ();
 FILLCELL_X32 FILLER_168_1186 ();
 FILLCELL_X32 FILLER_168_1218 ();
 FILLCELL_X32 FILLER_168_1250 ();
 FILLCELL_X32 FILLER_168_1282 ();
 FILLCELL_X32 FILLER_168_1314 ();
 FILLCELL_X32 FILLER_168_1346 ();
 FILLCELL_X32 FILLER_168_1378 ();
 FILLCELL_X32 FILLER_168_1410 ();
 FILLCELL_X32 FILLER_168_1442 ();
 FILLCELL_X32 FILLER_168_1474 ();
 FILLCELL_X32 FILLER_168_1506 ();
 FILLCELL_X32 FILLER_168_1538 ();
 FILLCELL_X32 FILLER_168_1570 ();
 FILLCELL_X32 FILLER_168_1602 ();
 FILLCELL_X16 FILLER_168_1634 ();
 FILLCELL_X1 FILLER_168_1650 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X4 FILLER_169_33 ();
 FILLCELL_X2 FILLER_169_37 ();
 FILLCELL_X1 FILLER_169_39 ();
 FILLCELL_X4 FILLER_169_47 ();
 FILLCELL_X2 FILLER_169_51 ();
 FILLCELL_X1 FILLER_169_90 ();
 FILLCELL_X4 FILLER_169_111 ();
 FILLCELL_X2 FILLER_169_133 ();
 FILLCELL_X2 FILLER_169_155 ();
 FILLCELL_X4 FILLER_169_184 ();
 FILLCELL_X16 FILLER_169_213 ();
 FILLCELL_X1 FILLER_169_229 ();
 FILLCELL_X2 FILLER_169_243 ();
 FILLCELL_X1 FILLER_169_245 ();
 FILLCELL_X1 FILLER_169_273 ();
 FILLCELL_X4 FILLER_169_281 ();
 FILLCELL_X2 FILLER_169_285 ();
 FILLCELL_X1 FILLER_169_287 ();
 FILLCELL_X2 FILLER_169_302 ();
 FILLCELL_X1 FILLER_169_307 ();
 FILLCELL_X1 FILLER_169_314 ();
 FILLCELL_X2 FILLER_169_319 ();
 FILLCELL_X16 FILLER_169_341 ();
 FILLCELL_X4 FILLER_169_361 ();
 FILLCELL_X1 FILLER_169_368 ();
 FILLCELL_X8 FILLER_169_378 ();
 FILLCELL_X2 FILLER_169_386 ();
 FILLCELL_X1 FILLER_169_415 ();
 FILLCELL_X1 FILLER_169_441 ();
 FILLCELL_X8 FILLER_169_447 ();
 FILLCELL_X4 FILLER_169_455 ();
 FILLCELL_X2 FILLER_169_459 ();
 FILLCELL_X1 FILLER_169_461 ();
 FILLCELL_X2 FILLER_169_482 ();
 FILLCELL_X2 FILLER_169_553 ();
 FILLCELL_X2 FILLER_169_564 ();
 FILLCELL_X2 FILLER_169_586 ();
 FILLCELL_X1 FILLER_169_588 ();
 FILLCELL_X4 FILLER_169_636 ();
 FILLCELL_X2 FILLER_169_660 ();
 FILLCELL_X1 FILLER_169_662 ();
 FILLCELL_X1 FILLER_169_703 ();
 FILLCELL_X1 FILLER_169_706 ();
 FILLCELL_X1 FILLER_169_712 ();
 FILLCELL_X8 FILLER_169_734 ();
 FILLCELL_X4 FILLER_169_742 ();
 FILLCELL_X2 FILLER_169_766 ();
 FILLCELL_X1 FILLER_169_768 ();
 FILLCELL_X1 FILLER_169_788 ();
 FILLCELL_X2 FILLER_169_801 ();
 FILLCELL_X2 FILLER_169_813 ();
 FILLCELL_X1 FILLER_169_815 ();
 FILLCELL_X2 FILLER_169_836 ();
 FILLCELL_X2 FILLER_169_845 ();
 FILLCELL_X2 FILLER_169_860 ();
 FILLCELL_X1 FILLER_169_862 ();
 FILLCELL_X1 FILLER_169_897 ();
 FILLCELL_X4 FILLER_169_927 ();
 FILLCELL_X1 FILLER_169_931 ();
 FILLCELL_X8 FILLER_169_952 ();
 FILLCELL_X4 FILLER_169_960 ();
 FILLCELL_X2 FILLER_169_964 ();
 FILLCELL_X1 FILLER_169_966 ();
 FILLCELL_X16 FILLER_169_974 ();
 FILLCELL_X2 FILLER_169_990 ();
 FILLCELL_X1 FILLER_169_1050 ();
 FILLCELL_X32 FILLER_169_1088 ();
 FILLCELL_X32 FILLER_169_1120 ();
 FILLCELL_X32 FILLER_169_1152 ();
 FILLCELL_X32 FILLER_169_1184 ();
 FILLCELL_X32 FILLER_169_1216 ();
 FILLCELL_X8 FILLER_169_1248 ();
 FILLCELL_X4 FILLER_169_1256 ();
 FILLCELL_X2 FILLER_169_1260 ();
 FILLCELL_X1 FILLER_169_1262 ();
 FILLCELL_X32 FILLER_169_1264 ();
 FILLCELL_X32 FILLER_169_1296 ();
 FILLCELL_X32 FILLER_169_1328 ();
 FILLCELL_X32 FILLER_169_1360 ();
 FILLCELL_X32 FILLER_169_1392 ();
 FILLCELL_X32 FILLER_169_1424 ();
 FILLCELL_X32 FILLER_169_1456 ();
 FILLCELL_X32 FILLER_169_1488 ();
 FILLCELL_X32 FILLER_169_1520 ();
 FILLCELL_X32 FILLER_169_1552 ();
 FILLCELL_X32 FILLER_169_1584 ();
 FILLCELL_X32 FILLER_169_1616 ();
 FILLCELL_X2 FILLER_169_1648 ();
 FILLCELL_X1 FILLER_169_1650 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X8 FILLER_170_33 ();
 FILLCELL_X1 FILLER_170_41 ();
 FILLCELL_X4 FILLER_170_74 ();
 FILLCELL_X2 FILLER_170_78 ();
 FILLCELL_X1 FILLER_170_87 ();
 FILLCELL_X4 FILLER_170_104 ();
 FILLCELL_X2 FILLER_170_108 ();
 FILLCELL_X16 FILLER_170_137 ();
 FILLCELL_X8 FILLER_170_153 ();
 FILLCELL_X2 FILLER_170_161 ();
 FILLCELL_X1 FILLER_170_217 ();
 FILLCELL_X8 FILLER_170_225 ();
 FILLCELL_X4 FILLER_170_233 ();
 FILLCELL_X8 FILLER_170_246 ();
 FILLCELL_X1 FILLER_170_283 ();
 FILLCELL_X1 FILLER_170_304 ();
 FILLCELL_X16 FILLER_170_313 ();
 FILLCELL_X8 FILLER_170_333 ();
 FILLCELL_X2 FILLER_170_341 ();
 FILLCELL_X1 FILLER_170_343 ();
 FILLCELL_X1 FILLER_170_347 ();
 FILLCELL_X2 FILLER_170_373 ();
 FILLCELL_X4 FILLER_170_395 ();
 FILLCELL_X1 FILLER_170_399 ();
 FILLCELL_X2 FILLER_170_404 ();
 FILLCELL_X1 FILLER_170_406 ();
 FILLCELL_X1 FILLER_170_417 ();
 FILLCELL_X1 FILLER_170_425 ();
 FILLCELL_X2 FILLER_170_430 ();
 FILLCELL_X2 FILLER_170_435 ();
 FILLCELL_X1 FILLER_170_437 ();
 FILLCELL_X1 FILLER_170_458 ();
 FILLCELL_X8 FILLER_170_466 ();
 FILLCELL_X4 FILLER_170_478 ();
 FILLCELL_X1 FILLER_170_482 ();
 FILLCELL_X8 FILLER_170_486 ();
 FILLCELL_X2 FILLER_170_494 ();
 FILLCELL_X1 FILLER_170_500 ();
 FILLCELL_X2 FILLER_170_504 ();
 FILLCELL_X8 FILLER_170_510 ();
 FILLCELL_X1 FILLER_170_528 ();
 FILLCELL_X8 FILLER_170_560 ();
 FILLCELL_X2 FILLER_170_568 ();
 FILLCELL_X8 FILLER_170_577 ();
 FILLCELL_X4 FILLER_170_585 ();
 FILLCELL_X1 FILLER_170_612 ();
 FILLCELL_X1 FILLER_170_616 ();
 FILLCELL_X4 FILLER_170_620 ();
 FILLCELL_X8 FILLER_170_632 ();
 FILLCELL_X2 FILLER_170_640 ();
 FILLCELL_X1 FILLER_170_642 ();
 FILLCELL_X16 FILLER_170_648 ();
 FILLCELL_X1 FILLER_170_664 ();
 FILLCELL_X4 FILLER_170_672 ();
 FILLCELL_X2 FILLER_170_676 ();
 FILLCELL_X1 FILLER_170_678 ();
 FILLCELL_X4 FILLER_170_692 ();
 FILLCELL_X1 FILLER_170_696 ();
 FILLCELL_X2 FILLER_170_717 ();
 FILLCELL_X1 FILLER_170_719 ();
 FILLCELL_X2 FILLER_170_740 ();
 FILLCELL_X4 FILLER_170_753 ();
 FILLCELL_X2 FILLER_170_757 ();
 FILLCELL_X4 FILLER_170_766 ();
 FILLCELL_X1 FILLER_170_770 ();
 FILLCELL_X1 FILLER_170_783 ();
 FILLCELL_X4 FILLER_170_811 ();
 FILLCELL_X2 FILLER_170_815 ();
 FILLCELL_X1 FILLER_170_817 ();
 FILLCELL_X8 FILLER_170_830 ();
 FILLCELL_X1 FILLER_170_838 ();
 FILLCELL_X8 FILLER_170_864 ();
 FILLCELL_X4 FILLER_170_872 ();
 FILLCELL_X2 FILLER_170_876 ();
 FILLCELL_X1 FILLER_170_878 ();
 FILLCELL_X2 FILLER_170_909 ();
 FILLCELL_X2 FILLER_170_927 ();
 FILLCELL_X2 FILLER_170_943 ();
 FILLCELL_X1 FILLER_170_945 ();
 FILLCELL_X4 FILLER_170_993 ();
 FILLCELL_X2 FILLER_170_997 ();
 FILLCELL_X1 FILLER_170_999 ();
 FILLCELL_X1 FILLER_170_1020 ();
 FILLCELL_X2 FILLER_170_1041 ();
 FILLCELL_X8 FILLER_170_1050 ();
 FILLCELL_X1 FILLER_170_1058 ();
 FILLCELL_X2 FILLER_170_1066 ();
 FILLCELL_X1 FILLER_170_1068 ();
 FILLCELL_X32 FILLER_170_1099 ();
 FILLCELL_X32 FILLER_170_1131 ();
 FILLCELL_X32 FILLER_170_1163 ();
 FILLCELL_X32 FILLER_170_1195 ();
 FILLCELL_X32 FILLER_170_1227 ();
 FILLCELL_X32 FILLER_170_1259 ();
 FILLCELL_X32 FILLER_170_1291 ();
 FILLCELL_X32 FILLER_170_1323 ();
 FILLCELL_X32 FILLER_170_1355 ();
 FILLCELL_X32 FILLER_170_1387 ();
 FILLCELL_X32 FILLER_170_1419 ();
 FILLCELL_X32 FILLER_170_1451 ();
 FILLCELL_X32 FILLER_170_1483 ();
 FILLCELL_X32 FILLER_170_1515 ();
 FILLCELL_X32 FILLER_170_1547 ();
 FILLCELL_X32 FILLER_170_1579 ();
 FILLCELL_X32 FILLER_170_1611 ();
 FILLCELL_X8 FILLER_170_1643 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X16 FILLER_171_33 ();
 FILLCELL_X2 FILLER_171_49 ();
 FILLCELL_X2 FILLER_171_78 ();
 FILLCELL_X1 FILLER_171_80 ();
 FILLCELL_X2 FILLER_171_88 ();
 FILLCELL_X1 FILLER_171_90 ();
 FILLCELL_X4 FILLER_171_118 ();
 FILLCELL_X1 FILLER_171_122 ();
 FILLCELL_X4 FILLER_171_128 ();
 FILLCELL_X2 FILLER_171_132 ();
 FILLCELL_X1 FILLER_171_134 ();
 FILLCELL_X4 FILLER_171_142 ();
 FILLCELL_X32 FILLER_171_173 ();
 FILLCELL_X16 FILLER_171_205 ();
 FILLCELL_X8 FILLER_171_241 ();
 FILLCELL_X8 FILLER_171_293 ();
 FILLCELL_X4 FILLER_171_301 ();
 FILLCELL_X2 FILLER_171_305 ();
 FILLCELL_X8 FILLER_171_311 ();
 FILLCELL_X4 FILLER_171_319 ();
 FILLCELL_X2 FILLER_171_347 ();
 FILLCELL_X4 FILLER_171_372 ();
 FILLCELL_X1 FILLER_171_388 ();
 FILLCELL_X16 FILLER_171_422 ();
 FILLCELL_X1 FILLER_171_438 ();
 FILLCELL_X4 FILLER_171_446 ();
 FILLCELL_X1 FILLER_171_472 ();
 FILLCELL_X2 FILLER_171_493 ();
 FILLCELL_X2 FILLER_171_498 ();
 FILLCELL_X2 FILLER_171_509 ();
 FILLCELL_X1 FILLER_171_511 ();
 FILLCELL_X2 FILLER_171_535 ();
 FILLCELL_X1 FILLER_171_537 ();
 FILLCELL_X2 FILLER_171_542 ();
 FILLCELL_X1 FILLER_171_544 ();
 FILLCELL_X8 FILLER_171_548 ();
 FILLCELL_X1 FILLER_171_580 ();
 FILLCELL_X8 FILLER_171_584 ();
 FILLCELL_X4 FILLER_171_592 ();
 FILLCELL_X2 FILLER_171_596 ();
 FILLCELL_X1 FILLER_171_602 ();
 FILLCELL_X8 FILLER_171_626 ();
 FILLCELL_X2 FILLER_171_638 ();
 FILLCELL_X4 FILLER_171_663 ();
 FILLCELL_X2 FILLER_171_667 ();
 FILLCELL_X1 FILLER_171_669 ();
 FILLCELL_X2 FILLER_171_698 ();
 FILLCELL_X2 FILLER_171_727 ();
 FILLCELL_X1 FILLER_171_729 ();
 FILLCELL_X8 FILLER_171_749 ();
 FILLCELL_X2 FILLER_171_757 ();
 FILLCELL_X1 FILLER_171_779 ();
 FILLCELL_X4 FILLER_171_808 ();
 FILLCELL_X1 FILLER_171_832 ();
 FILLCELL_X2 FILLER_171_853 ();
 FILLCELL_X16 FILLER_171_864 ();
 FILLCELL_X4 FILLER_171_880 ();
 FILLCELL_X1 FILLER_171_884 ();
 FILLCELL_X1 FILLER_171_894 ();
 FILLCELL_X2 FILLER_171_900 ();
 FILLCELL_X1 FILLER_171_902 ();
 FILLCELL_X2 FILLER_171_908 ();
 FILLCELL_X1 FILLER_171_910 ();
 FILLCELL_X1 FILLER_171_920 ();
 FILLCELL_X2 FILLER_171_934 ();
 FILLCELL_X1 FILLER_171_936 ();
 FILLCELL_X2 FILLER_171_944 ();
 FILLCELL_X2 FILLER_171_953 ();
 FILLCELL_X1 FILLER_171_969 ();
 FILLCELL_X1 FILLER_171_1000 ();
 FILLCELL_X4 FILLER_171_1012 ();
 FILLCELL_X1 FILLER_171_1016 ();
 FILLCELL_X8 FILLER_171_1024 ();
 FILLCELL_X1 FILLER_171_1032 ();
 FILLCELL_X1 FILLER_171_1046 ();
 FILLCELL_X32 FILLER_171_1067 ();
 FILLCELL_X32 FILLER_171_1099 ();
 FILLCELL_X32 FILLER_171_1131 ();
 FILLCELL_X32 FILLER_171_1163 ();
 FILLCELL_X32 FILLER_171_1195 ();
 FILLCELL_X32 FILLER_171_1227 ();
 FILLCELL_X4 FILLER_171_1259 ();
 FILLCELL_X32 FILLER_171_1264 ();
 FILLCELL_X32 FILLER_171_1296 ();
 FILLCELL_X32 FILLER_171_1328 ();
 FILLCELL_X32 FILLER_171_1360 ();
 FILLCELL_X32 FILLER_171_1392 ();
 FILLCELL_X32 FILLER_171_1424 ();
 FILLCELL_X32 FILLER_171_1456 ();
 FILLCELL_X32 FILLER_171_1488 ();
 FILLCELL_X32 FILLER_171_1520 ();
 FILLCELL_X32 FILLER_171_1552 ();
 FILLCELL_X32 FILLER_171_1584 ();
 FILLCELL_X32 FILLER_171_1616 ();
 FILLCELL_X2 FILLER_171_1648 ();
 FILLCELL_X1 FILLER_171_1650 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X16 FILLER_172_33 ();
 FILLCELL_X8 FILLER_172_49 ();
 FILLCELL_X4 FILLER_172_57 ();
 FILLCELL_X1 FILLER_172_61 ();
 FILLCELL_X2 FILLER_172_69 ();
 FILLCELL_X1 FILLER_172_71 ();
 FILLCELL_X1 FILLER_172_97 ();
 FILLCELL_X8 FILLER_172_109 ();
 FILLCELL_X4 FILLER_172_117 ();
 FILLCELL_X4 FILLER_172_141 ();
 FILLCELL_X4 FILLER_172_175 ();
 FILLCELL_X4 FILLER_172_188 ();
 FILLCELL_X1 FILLER_172_219 ();
 FILLCELL_X4 FILLER_172_253 ();
 FILLCELL_X2 FILLER_172_257 ();
 FILLCELL_X1 FILLER_172_259 ();
 FILLCELL_X8 FILLER_172_267 ();
 FILLCELL_X2 FILLER_172_275 ();
 FILLCELL_X1 FILLER_172_277 ();
 FILLCELL_X1 FILLER_172_282 ();
 FILLCELL_X2 FILLER_172_286 ();
 FILLCELL_X1 FILLER_172_288 ();
 FILLCELL_X2 FILLER_172_314 ();
 FILLCELL_X1 FILLER_172_336 ();
 FILLCELL_X1 FILLER_172_349 ();
 FILLCELL_X8 FILLER_172_354 ();
 FILLCELL_X4 FILLER_172_362 ();
 FILLCELL_X2 FILLER_172_366 ();
 FILLCELL_X8 FILLER_172_394 ();
 FILLCELL_X1 FILLER_172_402 ();
 FILLCELL_X1 FILLER_172_407 ();
 FILLCELL_X8 FILLER_172_439 ();
 FILLCELL_X2 FILLER_172_447 ();
 FILLCELL_X4 FILLER_172_473 ();
 FILLCELL_X2 FILLER_172_477 ();
 FILLCELL_X16 FILLER_172_510 ();
 FILLCELL_X8 FILLER_172_526 ();
 FILLCELL_X1 FILLER_172_534 ();
 FILLCELL_X8 FILLER_172_539 ();
 FILLCELL_X2 FILLER_172_547 ();
 FILLCELL_X1 FILLER_172_549 ();
 FILLCELL_X1 FILLER_172_565 ();
 FILLCELL_X4 FILLER_172_569 ();
 FILLCELL_X2 FILLER_172_573 ();
 FILLCELL_X8 FILLER_172_582 ();
 FILLCELL_X1 FILLER_172_590 ();
 FILLCELL_X1 FILLER_172_618 ();
 FILLCELL_X1 FILLER_172_630 ();
 FILLCELL_X2 FILLER_172_632 ();
 FILLCELL_X1 FILLER_172_634 ();
 FILLCELL_X1 FILLER_172_642 ();
 FILLCELL_X2 FILLER_172_688 ();
 FILLCELL_X1 FILLER_172_690 ();
 FILLCELL_X16 FILLER_172_707 ();
 FILLCELL_X8 FILLER_172_723 ();
 FILLCELL_X1 FILLER_172_731 ();
 FILLCELL_X1 FILLER_172_761 ();
 FILLCELL_X1 FILLER_172_767 ();
 FILLCELL_X1 FILLER_172_774 ();
 FILLCELL_X4 FILLER_172_782 ();
 FILLCELL_X1 FILLER_172_786 ();
 FILLCELL_X16 FILLER_172_794 ();
 FILLCELL_X8 FILLER_172_810 ();
 FILLCELL_X2 FILLER_172_821 ();
 FILLCELL_X2 FILLER_172_832 ();
 FILLCELL_X2 FILLER_172_841 ();
 FILLCELL_X1 FILLER_172_877 ();
 FILLCELL_X2 FILLER_172_882 ();
 FILLCELL_X2 FILLER_172_891 ();
 FILLCELL_X1 FILLER_172_893 ();
 FILLCELL_X1 FILLER_172_896 ();
 FILLCELL_X2 FILLER_172_901 ();
 FILLCELL_X1 FILLER_172_903 ();
 FILLCELL_X4 FILLER_172_918 ();
 FILLCELL_X2 FILLER_172_922 ();
 FILLCELL_X8 FILLER_172_931 ();
 FILLCELL_X1 FILLER_172_939 ();
 FILLCELL_X1 FILLER_172_953 ();
 FILLCELL_X2 FILLER_172_961 ();
 FILLCELL_X1 FILLER_172_968 ();
 FILLCELL_X16 FILLER_172_992 ();
 FILLCELL_X1 FILLER_172_1008 ();
 FILLCELL_X4 FILLER_172_1057 ();
 FILLCELL_X2 FILLER_172_1061 ();
 FILLCELL_X1 FILLER_172_1063 ();
 FILLCELL_X32 FILLER_172_1091 ();
 FILLCELL_X32 FILLER_172_1123 ();
 FILLCELL_X32 FILLER_172_1155 ();
 FILLCELL_X32 FILLER_172_1187 ();
 FILLCELL_X32 FILLER_172_1219 ();
 FILLCELL_X32 FILLER_172_1251 ();
 FILLCELL_X32 FILLER_172_1283 ();
 FILLCELL_X32 FILLER_172_1315 ();
 FILLCELL_X32 FILLER_172_1347 ();
 FILLCELL_X32 FILLER_172_1379 ();
 FILLCELL_X32 FILLER_172_1411 ();
 FILLCELL_X32 FILLER_172_1443 ();
 FILLCELL_X32 FILLER_172_1475 ();
 FILLCELL_X32 FILLER_172_1507 ();
 FILLCELL_X32 FILLER_172_1539 ();
 FILLCELL_X32 FILLER_172_1571 ();
 FILLCELL_X32 FILLER_172_1603 ();
 FILLCELL_X16 FILLER_172_1635 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X16 FILLER_173_33 ();
 FILLCELL_X8 FILLER_173_49 ();
 FILLCELL_X2 FILLER_173_57 ();
 FILLCELL_X1 FILLER_173_59 ();
 FILLCELL_X8 FILLER_173_80 ();
 FILLCELL_X2 FILLER_173_88 ();
 FILLCELL_X1 FILLER_173_116 ();
 FILLCELL_X1 FILLER_173_144 ();
 FILLCELL_X1 FILLER_173_150 ();
 FILLCELL_X1 FILLER_173_164 ();
 FILLCELL_X4 FILLER_173_192 ();
 FILLCELL_X1 FILLER_173_196 ();
 FILLCELL_X1 FILLER_173_233 ();
 FILLCELL_X8 FILLER_173_253 ();
 FILLCELL_X4 FILLER_173_261 ();
 FILLCELL_X2 FILLER_173_269 ();
 FILLCELL_X2 FILLER_173_274 ();
 FILLCELL_X4 FILLER_173_281 ();
 FILLCELL_X2 FILLER_173_285 ();
 FILLCELL_X1 FILLER_173_287 ();
 FILLCELL_X1 FILLER_173_292 ();
 FILLCELL_X1 FILLER_173_296 ();
 FILLCELL_X1 FILLER_173_302 ();
 FILLCELL_X2 FILLER_173_307 ();
 FILLCELL_X2 FILLER_173_312 ();
 FILLCELL_X1 FILLER_173_314 ();
 FILLCELL_X2 FILLER_173_322 ();
 FILLCELL_X2 FILLER_173_331 ();
 FILLCELL_X2 FILLER_173_337 ();
 FILLCELL_X1 FILLER_173_339 ();
 FILLCELL_X2 FILLER_173_346 ();
 FILLCELL_X1 FILLER_173_348 ();
 FILLCELL_X1 FILLER_173_369 ();
 FILLCELL_X2 FILLER_173_390 ();
 FILLCELL_X2 FILLER_173_435 ();
 FILLCELL_X1 FILLER_173_437 ();
 FILLCELL_X1 FILLER_173_449 ();
 FILLCELL_X2 FILLER_173_470 ();
 FILLCELL_X16 FILLER_173_475 ();
 FILLCELL_X2 FILLER_173_491 ();
 FILLCELL_X1 FILLER_173_493 ();
 FILLCELL_X1 FILLER_173_531 ();
 FILLCELL_X1 FILLER_173_552 ();
 FILLCELL_X1 FILLER_173_573 ();
 FILLCELL_X1 FILLER_173_594 ();
 FILLCELL_X1 FILLER_173_632 ();
 FILLCELL_X8 FILLER_173_653 ();
 FILLCELL_X4 FILLER_173_661 ();
 FILLCELL_X2 FILLER_173_665 ();
 FILLCELL_X1 FILLER_173_667 ();
 FILLCELL_X8 FILLER_173_716 ();
 FILLCELL_X4 FILLER_173_724 ();
 FILLCELL_X1 FILLER_173_728 ();
 FILLCELL_X1 FILLER_173_770 ();
 FILLCELL_X2 FILLER_173_796 ();
 FILLCELL_X1 FILLER_173_798 ();
 FILLCELL_X8 FILLER_173_803 ();
 FILLCELL_X16 FILLER_173_834 ();
 FILLCELL_X1 FILLER_173_884 ();
 FILLCELL_X2 FILLER_173_903 ();
 FILLCELL_X4 FILLER_173_918 ();
 FILLCELL_X8 FILLER_173_939 ();
 FILLCELL_X4 FILLER_173_947 ();
 FILLCELL_X1 FILLER_173_951 ();
 FILLCELL_X2 FILLER_173_1005 ();
 FILLCELL_X1 FILLER_173_1007 ();
 FILLCELL_X2 FILLER_173_1028 ();
 FILLCELL_X1 FILLER_173_1030 ();
 FILLCELL_X2 FILLER_173_1058 ();
 FILLCELL_X1 FILLER_173_1060 ();
 FILLCELL_X32 FILLER_173_1088 ();
 FILLCELL_X32 FILLER_173_1120 ();
 FILLCELL_X32 FILLER_173_1152 ();
 FILLCELL_X32 FILLER_173_1184 ();
 FILLCELL_X32 FILLER_173_1216 ();
 FILLCELL_X8 FILLER_173_1248 ();
 FILLCELL_X4 FILLER_173_1256 ();
 FILLCELL_X2 FILLER_173_1260 ();
 FILLCELL_X1 FILLER_173_1262 ();
 FILLCELL_X32 FILLER_173_1264 ();
 FILLCELL_X32 FILLER_173_1296 ();
 FILLCELL_X32 FILLER_173_1328 ();
 FILLCELL_X32 FILLER_173_1360 ();
 FILLCELL_X32 FILLER_173_1392 ();
 FILLCELL_X32 FILLER_173_1424 ();
 FILLCELL_X32 FILLER_173_1456 ();
 FILLCELL_X32 FILLER_173_1488 ();
 FILLCELL_X32 FILLER_173_1520 ();
 FILLCELL_X32 FILLER_173_1552 ();
 FILLCELL_X32 FILLER_173_1584 ();
 FILLCELL_X32 FILLER_173_1616 ();
 FILLCELL_X2 FILLER_173_1648 ();
 FILLCELL_X1 FILLER_173_1650 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X8 FILLER_174_33 ();
 FILLCELL_X2 FILLER_174_41 ();
 FILLCELL_X8 FILLER_174_92 ();
 FILLCELL_X1 FILLER_174_100 ();
 FILLCELL_X8 FILLER_174_156 ();
 FILLCELL_X4 FILLER_174_164 ();
 FILLCELL_X1 FILLER_174_168 ();
 FILLCELL_X4 FILLER_174_203 ();
 FILLCELL_X2 FILLER_174_207 ();
 FILLCELL_X1 FILLER_174_218 ();
 FILLCELL_X4 FILLER_174_228 ();
 FILLCELL_X4 FILLER_174_239 ();
 FILLCELL_X2 FILLER_174_243 ();
 FILLCELL_X4 FILLER_174_252 ();
 FILLCELL_X1 FILLER_174_256 ();
 FILLCELL_X1 FILLER_174_277 ();
 FILLCELL_X1 FILLER_174_318 ();
 FILLCELL_X2 FILLER_174_324 ();
 FILLCELL_X4 FILLER_174_346 ();
 FILLCELL_X2 FILLER_174_350 ();
 FILLCELL_X1 FILLER_174_352 ();
 FILLCELL_X2 FILLER_174_360 ();
 FILLCELL_X4 FILLER_174_369 ();
 FILLCELL_X2 FILLER_174_373 ();
 FILLCELL_X4 FILLER_174_382 ();
 FILLCELL_X2 FILLER_174_386 ();
 FILLCELL_X1 FILLER_174_388 ();
 FILLCELL_X4 FILLER_174_402 ();
 FILLCELL_X1 FILLER_174_406 ();
 FILLCELL_X4 FILLER_174_420 ();
 FILLCELL_X2 FILLER_174_424 ();
 FILLCELL_X1 FILLER_174_426 ();
 FILLCELL_X16 FILLER_174_431 ();
 FILLCELL_X2 FILLER_174_515 ();
 FILLCELL_X1 FILLER_174_517 ();
 FILLCELL_X4 FILLER_174_538 ();
 FILLCELL_X1 FILLER_174_542 ();
 FILLCELL_X4 FILLER_174_546 ();
 FILLCELL_X2 FILLER_174_550 ();
 FILLCELL_X1 FILLER_174_561 ();
 FILLCELL_X4 FILLER_174_566 ();
 FILLCELL_X2 FILLER_174_573 ();
 FILLCELL_X4 FILLER_174_589 ();
 FILLCELL_X4 FILLER_174_620 ();
 FILLCELL_X4 FILLER_174_660 ();
 FILLCELL_X2 FILLER_174_664 ();
 FILLCELL_X1 FILLER_174_666 ();
 FILLCELL_X8 FILLER_174_680 ();
 FILLCELL_X4 FILLER_174_688 ();
 FILLCELL_X1 FILLER_174_692 ();
 FILLCELL_X1 FILLER_174_700 ();
 FILLCELL_X8 FILLER_174_728 ();
 FILLCELL_X2 FILLER_174_736 ();
 FILLCELL_X1 FILLER_174_738 ();
 FILLCELL_X1 FILLER_174_746 ();
 FILLCELL_X4 FILLER_174_761 ();
 FILLCELL_X4 FILLER_174_792 ();
 FILLCELL_X2 FILLER_174_796 ();
 FILLCELL_X4 FILLER_174_818 ();
 FILLCELL_X2 FILLER_174_822 ();
 FILLCELL_X2 FILLER_174_844 ();
 FILLCELL_X8 FILLER_174_868 ();
 FILLCELL_X4 FILLER_174_876 ();
 FILLCELL_X4 FILLER_174_887 ();
 FILLCELL_X2 FILLER_174_891 ();
 FILLCELL_X2 FILLER_174_898 ();
 FILLCELL_X1 FILLER_174_916 ();
 FILLCELL_X1 FILLER_174_922 ();
 FILLCELL_X4 FILLER_174_936 ();
 FILLCELL_X1 FILLER_174_940 ();
 FILLCELL_X2 FILLER_174_948 ();
 FILLCELL_X8 FILLER_174_957 ();
 FILLCELL_X4 FILLER_174_965 ();
 FILLCELL_X4 FILLER_174_996 ();
 FILLCELL_X2 FILLER_174_1000 ();
 FILLCELL_X1 FILLER_174_1002 ();
 FILLCELL_X8 FILLER_174_1016 ();
 FILLCELL_X4 FILLER_174_1024 ();
 FILLCELL_X2 FILLER_174_1028 ();
 FILLCELL_X1 FILLER_174_1030 ();
 FILLCELL_X2 FILLER_174_1038 ();
 FILLCELL_X1 FILLER_174_1040 ();
 FILLCELL_X8 FILLER_174_1055 ();
 FILLCELL_X1 FILLER_174_1063 ();
 FILLCELL_X32 FILLER_174_1091 ();
 FILLCELL_X32 FILLER_174_1123 ();
 FILLCELL_X32 FILLER_174_1155 ();
 FILLCELL_X32 FILLER_174_1187 ();
 FILLCELL_X32 FILLER_174_1219 ();
 FILLCELL_X32 FILLER_174_1251 ();
 FILLCELL_X32 FILLER_174_1283 ();
 FILLCELL_X32 FILLER_174_1315 ();
 FILLCELL_X32 FILLER_174_1347 ();
 FILLCELL_X32 FILLER_174_1379 ();
 FILLCELL_X32 FILLER_174_1411 ();
 FILLCELL_X32 FILLER_174_1443 ();
 FILLCELL_X32 FILLER_174_1475 ();
 FILLCELL_X32 FILLER_174_1507 ();
 FILLCELL_X32 FILLER_174_1539 ();
 FILLCELL_X32 FILLER_174_1571 ();
 FILLCELL_X32 FILLER_174_1603 ();
 FILLCELL_X16 FILLER_174_1635 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X16 FILLER_175_33 ();
 FILLCELL_X8 FILLER_175_49 ();
 FILLCELL_X2 FILLER_175_57 ();
 FILLCELL_X8 FILLER_175_67 ();
 FILLCELL_X1 FILLER_175_129 ();
 FILLCELL_X16 FILLER_175_164 ();
 FILLCELL_X4 FILLER_175_180 ();
 FILLCELL_X1 FILLER_175_184 ();
 FILLCELL_X4 FILLER_175_192 ();
 FILLCELL_X2 FILLER_175_196 ();
 FILLCELL_X8 FILLER_175_207 ();
 FILLCELL_X1 FILLER_175_215 ();
 FILLCELL_X4 FILLER_175_252 ();
 FILLCELL_X1 FILLER_175_276 ();
 FILLCELL_X4 FILLER_175_297 ();
 FILLCELL_X2 FILLER_175_301 ();
 FILLCELL_X2 FILLER_175_323 ();
 FILLCELL_X1 FILLER_175_325 ();
 FILLCELL_X2 FILLER_175_346 ();
 FILLCELL_X4 FILLER_175_368 ();
 FILLCELL_X16 FILLER_175_379 ();
 FILLCELL_X4 FILLER_175_395 ();
 FILLCELL_X2 FILLER_175_419 ();
 FILLCELL_X2 FILLER_175_428 ();
 FILLCELL_X1 FILLER_175_443 ();
 FILLCELL_X1 FILLER_175_464 ();
 FILLCELL_X1 FILLER_175_485 ();
 FILLCELL_X2 FILLER_175_489 ();
 FILLCELL_X1 FILLER_175_519 ();
 FILLCELL_X2 FILLER_175_526 ();
 FILLCELL_X1 FILLER_175_548 ();
 FILLCELL_X2 FILLER_175_552 ();
 FILLCELL_X2 FILLER_175_559 ();
 FILLCELL_X1 FILLER_175_581 ();
 FILLCELL_X1 FILLER_175_594 ();
 FILLCELL_X4 FILLER_175_604 ();
 FILLCELL_X2 FILLER_175_608 ();
 FILLCELL_X16 FILLER_175_630 ();
 FILLCELL_X4 FILLER_175_646 ();
 FILLCELL_X2 FILLER_175_650 ();
 FILLCELL_X16 FILLER_175_659 ();
 FILLCELL_X2 FILLER_175_675 ();
 FILLCELL_X1 FILLER_175_677 ();
 FILLCELL_X4 FILLER_175_704 ();
 FILLCELL_X16 FILLER_175_717 ();
 FILLCELL_X4 FILLER_175_733 ();
 FILLCELL_X4 FILLER_175_744 ();
 FILLCELL_X2 FILLER_175_748 ();
 FILLCELL_X1 FILLER_175_750 ();
 FILLCELL_X16 FILLER_175_765 ();
 FILLCELL_X2 FILLER_175_781 ();
 FILLCELL_X8 FILLER_175_812 ();
 FILLCELL_X1 FILLER_175_820 ();
 FILLCELL_X2 FILLER_175_828 ();
 FILLCELL_X4 FILLER_175_837 ();
 FILLCELL_X1 FILLER_175_841 ();
 FILLCELL_X8 FILLER_175_854 ();
 FILLCELL_X4 FILLER_175_862 ();
 FILLCELL_X1 FILLER_175_866 ();
 FILLCELL_X2 FILLER_175_874 ();
 FILLCELL_X2 FILLER_175_912 ();
 FILLCELL_X1 FILLER_175_914 ();
 FILLCELL_X4 FILLER_175_924 ();
 FILLCELL_X2 FILLER_175_928 ();
 FILLCELL_X2 FILLER_175_950 ();
 FILLCELL_X4 FILLER_175_972 ();
 FILLCELL_X2 FILLER_175_983 ();
 FILLCELL_X1 FILLER_175_985 ();
 FILLCELL_X4 FILLER_175_1013 ();
 FILLCELL_X1 FILLER_175_1017 ();
 FILLCELL_X32 FILLER_175_1051 ();
 FILLCELL_X32 FILLER_175_1083 ();
 FILLCELL_X32 FILLER_175_1115 ();
 FILLCELL_X32 FILLER_175_1147 ();
 FILLCELL_X32 FILLER_175_1179 ();
 FILLCELL_X32 FILLER_175_1211 ();
 FILLCELL_X16 FILLER_175_1243 ();
 FILLCELL_X4 FILLER_175_1259 ();
 FILLCELL_X32 FILLER_175_1264 ();
 FILLCELL_X32 FILLER_175_1296 ();
 FILLCELL_X32 FILLER_175_1328 ();
 FILLCELL_X32 FILLER_175_1360 ();
 FILLCELL_X32 FILLER_175_1392 ();
 FILLCELL_X32 FILLER_175_1424 ();
 FILLCELL_X32 FILLER_175_1456 ();
 FILLCELL_X32 FILLER_175_1488 ();
 FILLCELL_X32 FILLER_175_1520 ();
 FILLCELL_X32 FILLER_175_1552 ();
 FILLCELL_X32 FILLER_175_1584 ();
 FILLCELL_X32 FILLER_175_1616 ();
 FILLCELL_X2 FILLER_175_1648 ();
 FILLCELL_X1 FILLER_175_1650 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X16 FILLER_176_33 ();
 FILLCELL_X2 FILLER_176_49 ();
 FILLCELL_X1 FILLER_176_51 ();
 FILLCELL_X4 FILLER_176_86 ();
 FILLCELL_X16 FILLER_176_95 ();
 FILLCELL_X2 FILLER_176_111 ();
 FILLCELL_X1 FILLER_176_113 ();
 FILLCELL_X16 FILLER_176_141 ();
 FILLCELL_X2 FILLER_176_157 ();
 FILLCELL_X1 FILLER_176_159 ();
 FILLCELL_X4 FILLER_176_174 ();
 FILLCELL_X1 FILLER_176_178 ();
 FILLCELL_X2 FILLER_176_199 ();
 FILLCELL_X1 FILLER_176_201 ();
 FILLCELL_X2 FILLER_176_231 ();
 FILLCELL_X1 FILLER_176_233 ();
 FILLCELL_X8 FILLER_176_254 ();
 FILLCELL_X1 FILLER_176_262 ();
 FILLCELL_X2 FILLER_176_267 ();
 FILLCELL_X1 FILLER_176_272 ();
 FILLCELL_X2 FILLER_176_280 ();
 FILLCELL_X4 FILLER_176_286 ();
 FILLCELL_X4 FILLER_176_300 ();
 FILLCELL_X1 FILLER_176_304 ();
 FILLCELL_X1 FILLER_176_327 ();
 FILLCELL_X1 FILLER_176_348 ();
 FILLCELL_X1 FILLER_176_369 ();
 FILLCELL_X1 FILLER_176_384 ();
 FILLCELL_X2 FILLER_176_389 ();
 FILLCELL_X2 FILLER_176_394 ();
 FILLCELL_X2 FILLER_176_401 ();
 FILLCELL_X1 FILLER_176_403 ();
 FILLCELL_X1 FILLER_176_445 ();
 FILLCELL_X4 FILLER_176_450 ();
 FILLCELL_X1 FILLER_176_454 ();
 FILLCELL_X8 FILLER_176_458 ();
 FILLCELL_X1 FILLER_176_466 ();
 FILLCELL_X2 FILLER_176_495 ();
 FILLCELL_X4 FILLER_176_501 ();
 FILLCELL_X1 FILLER_176_505 ();
 FILLCELL_X4 FILLER_176_509 ();
 FILLCELL_X1 FILLER_176_513 ();
 FILLCELL_X8 FILLER_176_519 ();
 FILLCELL_X2 FILLER_176_527 ();
 FILLCELL_X4 FILLER_176_560 ();
 FILLCELL_X1 FILLER_176_564 ();
 FILLCELL_X2 FILLER_176_569 ();
 FILLCELL_X4 FILLER_176_627 ();
 FILLCELL_X1 FILLER_176_655 ();
 FILLCELL_X1 FILLER_176_676 ();
 FILLCELL_X1 FILLER_176_694 ();
 FILLCELL_X16 FILLER_176_711 ();
 FILLCELL_X8 FILLER_176_727 ();
 FILLCELL_X4 FILLER_176_735 ();
 FILLCELL_X1 FILLER_176_739 ();
 FILLCELL_X2 FILLER_176_771 ();
 FILLCELL_X1 FILLER_176_773 ();
 FILLCELL_X4 FILLER_176_795 ();
 FILLCELL_X2 FILLER_176_806 ();
 FILLCELL_X2 FILLER_176_812 ();
 FILLCELL_X4 FILLER_176_834 ();
 FILLCELL_X1 FILLER_176_838 ();
 FILLCELL_X2 FILLER_176_866 ();
 FILLCELL_X1 FILLER_176_868 ();
 FILLCELL_X16 FILLER_176_889 ();
 FILLCELL_X2 FILLER_176_905 ();
 FILLCELL_X1 FILLER_176_907 ();
 FILLCELL_X2 FILLER_176_921 ();
 FILLCELL_X16 FILLER_176_936 ();
 FILLCELL_X8 FILLER_176_960 ();
 FILLCELL_X4 FILLER_176_968 ();
 FILLCELL_X2 FILLER_176_972 ();
 FILLCELL_X1 FILLER_176_974 ();
 FILLCELL_X16 FILLER_176_1008 ();
 FILLCELL_X8 FILLER_176_1024 ();
 FILLCELL_X32 FILLER_176_1045 ();
 FILLCELL_X32 FILLER_176_1077 ();
 FILLCELL_X32 FILLER_176_1109 ();
 FILLCELL_X32 FILLER_176_1141 ();
 FILLCELL_X32 FILLER_176_1173 ();
 FILLCELL_X32 FILLER_176_1205 ();
 FILLCELL_X32 FILLER_176_1237 ();
 FILLCELL_X32 FILLER_176_1269 ();
 FILLCELL_X32 FILLER_176_1301 ();
 FILLCELL_X32 FILLER_176_1333 ();
 FILLCELL_X32 FILLER_176_1365 ();
 FILLCELL_X32 FILLER_176_1397 ();
 FILLCELL_X32 FILLER_176_1429 ();
 FILLCELL_X32 FILLER_176_1461 ();
 FILLCELL_X32 FILLER_176_1493 ();
 FILLCELL_X32 FILLER_176_1525 ();
 FILLCELL_X32 FILLER_176_1557 ();
 FILLCELL_X32 FILLER_176_1589 ();
 FILLCELL_X16 FILLER_176_1621 ();
 FILLCELL_X8 FILLER_176_1637 ();
 FILLCELL_X4 FILLER_176_1645 ();
 FILLCELL_X2 FILLER_176_1649 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X8 FILLER_177_65 ();
 FILLCELL_X4 FILLER_177_73 ();
 FILLCELL_X1 FILLER_177_77 ();
 FILLCELL_X1 FILLER_177_127 ();
 FILLCELL_X2 FILLER_177_133 ();
 FILLCELL_X1 FILLER_177_135 ();
 FILLCELL_X2 FILLER_177_150 ();
 FILLCELL_X1 FILLER_177_152 ();
 FILLCELL_X8 FILLER_177_180 ();
 FILLCELL_X2 FILLER_177_188 ();
 FILLCELL_X4 FILLER_177_197 ();
 FILLCELL_X2 FILLER_177_201 ();
 FILLCELL_X8 FILLER_177_257 ();
 FILLCELL_X2 FILLER_177_265 ();
 FILLCELL_X1 FILLER_177_267 ();
 FILLCELL_X2 FILLER_177_288 ();
 FILLCELL_X8 FILLER_177_317 ();
 FILLCELL_X2 FILLER_177_325 ();
 FILLCELL_X1 FILLER_177_327 ();
 FILLCELL_X4 FILLER_177_333 ();
 FILLCELL_X1 FILLER_177_337 ();
 FILLCELL_X2 FILLER_177_349 ();
 FILLCELL_X1 FILLER_177_351 ();
 FILLCELL_X2 FILLER_177_356 ();
 FILLCELL_X2 FILLER_177_361 ();
 FILLCELL_X1 FILLER_177_363 ();
 FILLCELL_X2 FILLER_177_369 ();
 FILLCELL_X1 FILLER_177_371 ();
 FILLCELL_X2 FILLER_177_378 ();
 FILLCELL_X4 FILLER_177_406 ();
 FILLCELL_X1 FILLER_177_410 ();
 FILLCELL_X8 FILLER_177_418 ();
 FILLCELL_X2 FILLER_177_426 ();
 FILLCELL_X8 FILLER_177_432 ();
 FILLCELL_X2 FILLER_177_440 ();
 FILLCELL_X4 FILLER_177_465 ();
 FILLCELL_X2 FILLER_177_469 ();
 FILLCELL_X2 FILLER_177_478 ();
 FILLCELL_X8 FILLER_177_488 ();
 FILLCELL_X1 FILLER_177_496 ();
 FILLCELL_X2 FILLER_177_517 ();
 FILLCELL_X2 FILLER_177_539 ();
 FILLCELL_X1 FILLER_177_590 ();
 FILLCELL_X2 FILLER_177_605 ();
 FILLCELL_X2 FILLER_177_627 ();
 FILLCELL_X1 FILLER_177_629 ();
 FILLCELL_X2 FILLER_177_644 ();
 FILLCELL_X8 FILLER_177_666 ();
 FILLCELL_X4 FILLER_177_674 ();
 FILLCELL_X2 FILLER_177_678 ();
 FILLCELL_X2 FILLER_177_726 ();
 FILLCELL_X16 FILLER_177_774 ();
 FILLCELL_X8 FILLER_177_790 ();
 FILLCELL_X2 FILLER_177_798 ();
 FILLCELL_X2 FILLER_177_813 ();
 FILLCELL_X4 FILLER_177_824 ();
 FILLCELL_X2 FILLER_177_828 ();
 FILLCELL_X1 FILLER_177_834 ();
 FILLCELL_X4 FILLER_177_844 ();
 FILLCELL_X1 FILLER_177_848 ();
 FILLCELL_X4 FILLER_177_858 ();
 FILLCELL_X8 FILLER_177_882 ();
 FILLCELL_X4 FILLER_177_890 ();
 FILLCELL_X2 FILLER_177_894 ();
 FILLCELL_X4 FILLER_177_918 ();
 FILLCELL_X4 FILLER_177_926 ();
 FILLCELL_X2 FILLER_177_934 ();
 FILLCELL_X4 FILLER_177_938 ();
 FILLCELL_X2 FILLER_177_950 ();
 FILLCELL_X2 FILLER_177_956 ();
 FILLCELL_X2 FILLER_177_985 ();
 FILLCELL_X8 FILLER_177_1021 ();
 FILLCELL_X4 FILLER_177_1042 ();
 FILLCELL_X1 FILLER_177_1046 ();
 FILLCELL_X2 FILLER_177_1060 ();
 FILLCELL_X1 FILLER_177_1062 ();
 FILLCELL_X32 FILLER_177_1076 ();
 FILLCELL_X32 FILLER_177_1108 ();
 FILLCELL_X32 FILLER_177_1140 ();
 FILLCELL_X32 FILLER_177_1172 ();
 FILLCELL_X32 FILLER_177_1204 ();
 FILLCELL_X16 FILLER_177_1236 ();
 FILLCELL_X8 FILLER_177_1252 ();
 FILLCELL_X2 FILLER_177_1260 ();
 FILLCELL_X1 FILLER_177_1262 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X32 FILLER_177_1296 ();
 FILLCELL_X32 FILLER_177_1328 ();
 FILLCELL_X32 FILLER_177_1360 ();
 FILLCELL_X32 FILLER_177_1392 ();
 FILLCELL_X32 FILLER_177_1424 ();
 FILLCELL_X32 FILLER_177_1456 ();
 FILLCELL_X32 FILLER_177_1488 ();
 FILLCELL_X32 FILLER_177_1520 ();
 FILLCELL_X32 FILLER_177_1552 ();
 FILLCELL_X32 FILLER_177_1584 ();
 FILLCELL_X32 FILLER_177_1616 ();
 FILLCELL_X2 FILLER_177_1648 ();
 FILLCELL_X1 FILLER_177_1650 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X16 FILLER_178_97 ();
 FILLCELL_X8 FILLER_178_113 ();
 FILLCELL_X4 FILLER_178_141 ();
 FILLCELL_X4 FILLER_178_165 ();
 FILLCELL_X8 FILLER_178_178 ();
 FILLCELL_X8 FILLER_178_206 ();
 FILLCELL_X2 FILLER_178_214 ();
 FILLCELL_X1 FILLER_178_216 ();
 FILLCELL_X1 FILLER_178_224 ();
 FILLCELL_X4 FILLER_178_232 ();
 FILLCELL_X2 FILLER_178_236 ();
 FILLCELL_X1 FILLER_178_238 ();
 FILLCELL_X4 FILLER_178_251 ();
 FILLCELL_X2 FILLER_178_255 ();
 FILLCELL_X1 FILLER_178_257 ();
 FILLCELL_X2 FILLER_178_307 ();
 FILLCELL_X16 FILLER_178_329 ();
 FILLCELL_X8 FILLER_178_345 ();
 FILLCELL_X1 FILLER_178_353 ();
 FILLCELL_X4 FILLER_178_358 ();
 FILLCELL_X4 FILLER_178_365 ();
 FILLCELL_X2 FILLER_178_374 ();
 FILLCELL_X1 FILLER_178_376 ();
 FILLCELL_X4 FILLER_178_417 ();
 FILLCELL_X1 FILLER_178_446 ();
 FILLCELL_X1 FILLER_178_471 ();
 FILLCELL_X4 FILLER_178_492 ();
 FILLCELL_X1 FILLER_178_496 ();
 FILLCELL_X2 FILLER_178_542 ();
 FILLCELL_X4 FILLER_178_557 ();
 FILLCELL_X1 FILLER_178_561 ();
 FILLCELL_X2 FILLER_178_585 ();
 FILLCELL_X2 FILLER_178_592 ();
 FILLCELL_X4 FILLER_178_603 ();
 FILLCELL_X8 FILLER_178_614 ();
 FILLCELL_X2 FILLER_178_622 ();
 FILLCELL_X2 FILLER_178_646 ();
 FILLCELL_X8 FILLER_178_666 ();
 FILLCELL_X2 FILLER_178_674 ();
 FILLCELL_X8 FILLER_178_685 ();
 FILLCELL_X2 FILLER_178_693 ();
 FILLCELL_X1 FILLER_178_695 ();
 FILLCELL_X2 FILLER_178_723 ();
 FILLCELL_X2 FILLER_178_738 ();
 FILLCELL_X1 FILLER_178_740 ();
 FILLCELL_X2 FILLER_178_744 ();
 FILLCELL_X16 FILLER_178_780 ();
 FILLCELL_X4 FILLER_178_796 ();
 FILLCELL_X2 FILLER_178_800 ();
 FILLCELL_X1 FILLER_178_802 ();
 FILLCELL_X2 FILLER_178_810 ();
 FILLCELL_X1 FILLER_178_812 ();
 FILLCELL_X1 FILLER_178_839 ();
 FILLCELL_X2 FILLER_178_858 ();
 FILLCELL_X4 FILLER_178_868 ();
 FILLCELL_X1 FILLER_178_872 ();
 FILLCELL_X4 FILLER_178_876 ();
 FILLCELL_X4 FILLER_178_887 ();
 FILLCELL_X2 FILLER_178_891 ();
 FILLCELL_X1 FILLER_178_893 ();
 FILLCELL_X4 FILLER_178_929 ();
 FILLCELL_X2 FILLER_178_933 ();
 FILLCELL_X1 FILLER_178_935 ();
 FILLCELL_X8 FILLER_178_984 ();
 FILLCELL_X4 FILLER_178_992 ();
 FILLCELL_X2 FILLER_178_996 ();
 FILLCELL_X4 FILLER_178_1005 ();
 FILLCELL_X1 FILLER_178_1009 ();
 FILLCELL_X32 FILLER_178_1051 ();
 FILLCELL_X32 FILLER_178_1083 ();
 FILLCELL_X32 FILLER_178_1115 ();
 FILLCELL_X32 FILLER_178_1147 ();
 FILLCELL_X32 FILLER_178_1179 ();
 FILLCELL_X32 FILLER_178_1211 ();
 FILLCELL_X32 FILLER_178_1243 ();
 FILLCELL_X32 FILLER_178_1275 ();
 FILLCELL_X32 FILLER_178_1307 ();
 FILLCELL_X32 FILLER_178_1339 ();
 FILLCELL_X32 FILLER_178_1371 ();
 FILLCELL_X32 FILLER_178_1403 ();
 FILLCELL_X32 FILLER_178_1435 ();
 FILLCELL_X32 FILLER_178_1467 ();
 FILLCELL_X32 FILLER_178_1499 ();
 FILLCELL_X32 FILLER_178_1531 ();
 FILLCELL_X32 FILLER_178_1563 ();
 FILLCELL_X32 FILLER_178_1595 ();
 FILLCELL_X16 FILLER_178_1627 ();
 FILLCELL_X8 FILLER_178_1643 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X16 FILLER_179_129 ();
 FILLCELL_X4 FILLER_179_152 ();
 FILLCELL_X2 FILLER_179_156 ();
 FILLCELL_X1 FILLER_179_158 ();
 FILLCELL_X8 FILLER_179_188 ();
 FILLCELL_X2 FILLER_179_196 ();
 FILLCELL_X1 FILLER_179_198 ();
 FILLCELL_X1 FILLER_179_213 ();
 FILLCELL_X1 FILLER_179_234 ();
 FILLCELL_X4 FILLER_179_240 ();
 FILLCELL_X1 FILLER_179_269 ();
 FILLCELL_X1 FILLER_179_297 ();
 FILLCELL_X1 FILLER_179_318 ();
 FILLCELL_X1 FILLER_179_346 ();
 FILLCELL_X1 FILLER_179_367 ();
 FILLCELL_X2 FILLER_179_388 ();
 FILLCELL_X1 FILLER_179_398 ();
 FILLCELL_X8 FILLER_179_403 ();
 FILLCELL_X1 FILLER_179_421 ();
 FILLCELL_X1 FILLER_179_440 ();
 FILLCELL_X4 FILLER_179_465 ();
 FILLCELL_X2 FILLER_179_469 ();
 FILLCELL_X1 FILLER_179_471 ();
 FILLCELL_X1 FILLER_179_479 ();
 FILLCELL_X1 FILLER_179_507 ();
 FILLCELL_X4 FILLER_179_515 ();
 FILLCELL_X1 FILLER_179_519 ();
 FILLCELL_X4 FILLER_179_534 ();
 FILLCELL_X2 FILLER_179_538 ();
 FILLCELL_X1 FILLER_179_540 ();
 FILLCELL_X2 FILLER_179_563 ();
 FILLCELL_X1 FILLER_179_565 ();
 FILLCELL_X4 FILLER_179_569 ();
 FILLCELL_X2 FILLER_179_573 ();
 FILLCELL_X1 FILLER_179_579 ();
 FILLCELL_X4 FILLER_179_584 ();
 FILLCELL_X2 FILLER_179_606 ();
 FILLCELL_X4 FILLER_179_668 ();
 FILLCELL_X1 FILLER_179_672 ();
 FILLCELL_X16 FILLER_179_736 ();
 FILLCELL_X8 FILLER_179_752 ();
 FILLCELL_X2 FILLER_179_760 ();
 FILLCELL_X4 FILLER_179_791 ();
 FILLCELL_X2 FILLER_179_795 ();
 FILLCELL_X1 FILLER_179_808 ();
 FILLCELL_X8 FILLER_179_816 ();
 FILLCELL_X4 FILLER_179_824 ();
 FILLCELL_X4 FILLER_179_846 ();
 FILLCELL_X1 FILLER_179_850 ();
 FILLCELL_X2 FILLER_179_864 ();
 FILLCELL_X1 FILLER_179_871 ();
 FILLCELL_X8 FILLER_179_897 ();
 FILLCELL_X1 FILLER_179_905 ();
 FILLCELL_X16 FILLER_179_959 ();
 FILLCELL_X4 FILLER_179_985 ();
 FILLCELL_X1 FILLER_179_989 ();
 FILLCELL_X4 FILLER_179_995 ();
 FILLCELL_X1 FILLER_179_1031 ();
 FILLCELL_X32 FILLER_179_1059 ();
 FILLCELL_X32 FILLER_179_1091 ();
 FILLCELL_X32 FILLER_179_1123 ();
 FILLCELL_X32 FILLER_179_1155 ();
 FILLCELL_X32 FILLER_179_1187 ();
 FILLCELL_X32 FILLER_179_1219 ();
 FILLCELL_X8 FILLER_179_1251 ();
 FILLCELL_X4 FILLER_179_1259 ();
 FILLCELL_X32 FILLER_179_1264 ();
 FILLCELL_X32 FILLER_179_1296 ();
 FILLCELL_X32 FILLER_179_1328 ();
 FILLCELL_X32 FILLER_179_1360 ();
 FILLCELL_X32 FILLER_179_1392 ();
 FILLCELL_X32 FILLER_179_1424 ();
 FILLCELL_X32 FILLER_179_1456 ();
 FILLCELL_X32 FILLER_179_1488 ();
 FILLCELL_X32 FILLER_179_1520 ();
 FILLCELL_X32 FILLER_179_1552 ();
 FILLCELL_X32 FILLER_179_1584 ();
 FILLCELL_X32 FILLER_179_1616 ();
 FILLCELL_X2 FILLER_179_1648 ();
 FILLCELL_X1 FILLER_179_1650 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X4 FILLER_180_129 ();
 FILLCELL_X2 FILLER_180_133 ();
 FILLCELL_X1 FILLER_180_135 ();
 FILLCELL_X4 FILLER_180_175 ();
 FILLCELL_X2 FILLER_180_192 ();
 FILLCELL_X4 FILLER_180_203 ();
 FILLCELL_X4 FILLER_180_227 ();
 FILLCELL_X2 FILLER_180_236 ();
 FILLCELL_X1 FILLER_180_238 ();
 FILLCELL_X16 FILLER_180_246 ();
 FILLCELL_X2 FILLER_180_262 ();
 FILLCELL_X4 FILLER_180_267 ();
 FILLCELL_X2 FILLER_180_271 ();
 FILLCELL_X1 FILLER_180_273 ();
 FILLCELL_X2 FILLER_180_301 ();
 FILLCELL_X2 FILLER_180_330 ();
 FILLCELL_X2 FILLER_180_337 ();
 FILLCELL_X2 FILLER_180_344 ();
 FILLCELL_X8 FILLER_180_379 ();
 FILLCELL_X2 FILLER_180_387 ();
 FILLCELL_X4 FILLER_180_409 ();
 FILLCELL_X2 FILLER_180_433 ();
 FILLCELL_X16 FILLER_180_491 ();
 FILLCELL_X8 FILLER_180_507 ();
 FILLCELL_X2 FILLER_180_515 ();
 FILLCELL_X1 FILLER_180_517 ();
 FILLCELL_X16 FILLER_180_526 ();
 FILLCELL_X8 FILLER_180_542 ();
 FILLCELL_X1 FILLER_180_568 ();
 FILLCELL_X1 FILLER_180_578 ();
 FILLCELL_X8 FILLER_180_599 ();
 FILLCELL_X16 FILLER_180_611 ();
 FILLCELL_X4 FILLER_180_627 ();
 FILLCELL_X8 FILLER_180_636 ();
 FILLCELL_X2 FILLER_180_644 ();
 FILLCELL_X8 FILLER_180_679 ();
 FILLCELL_X16 FILLER_180_725 ();
 FILLCELL_X2 FILLER_180_741 ();
 FILLCELL_X1 FILLER_180_743 ();
 FILLCELL_X4 FILLER_180_751 ();
 FILLCELL_X2 FILLER_180_755 ();
 FILLCELL_X2 FILLER_180_768 ();
 FILLCELL_X2 FILLER_180_774 ();
 FILLCELL_X1 FILLER_180_776 ();
 FILLCELL_X8 FILLER_180_784 ();
 FILLCELL_X4 FILLER_180_792 ();
 FILLCELL_X4 FILLER_180_823 ();
 FILLCELL_X1 FILLER_180_827 ();
 FILLCELL_X4 FILLER_180_846 ();
 FILLCELL_X4 FILLER_180_857 ();
 FILLCELL_X4 FILLER_180_881 ();
 FILLCELL_X2 FILLER_180_885 ();
 FILLCELL_X4 FILLER_180_891 ();
 FILLCELL_X4 FILLER_180_912 ();
 FILLCELL_X2 FILLER_180_916 ();
 FILLCELL_X2 FILLER_180_935 ();
 FILLCELL_X1 FILLER_180_937 ();
 FILLCELL_X1 FILLER_180_971 ();
 FILLCELL_X2 FILLER_180_979 ();
 FILLCELL_X1 FILLER_180_988 ();
 FILLCELL_X2 FILLER_180_994 ();
 FILLCELL_X4 FILLER_180_1016 ();
 FILLCELL_X1 FILLER_180_1020 ();
 FILLCELL_X2 FILLER_180_1025 ();
 FILLCELL_X2 FILLER_180_1047 ();
 FILLCELL_X1 FILLER_180_1049 ();
 FILLCELL_X32 FILLER_180_1063 ();
 FILLCELL_X32 FILLER_180_1095 ();
 FILLCELL_X32 FILLER_180_1127 ();
 FILLCELL_X32 FILLER_180_1159 ();
 FILLCELL_X32 FILLER_180_1191 ();
 FILLCELL_X32 FILLER_180_1223 ();
 FILLCELL_X32 FILLER_180_1255 ();
 FILLCELL_X32 FILLER_180_1287 ();
 FILLCELL_X32 FILLER_180_1319 ();
 FILLCELL_X32 FILLER_180_1351 ();
 FILLCELL_X32 FILLER_180_1383 ();
 FILLCELL_X32 FILLER_180_1415 ();
 FILLCELL_X32 FILLER_180_1447 ();
 FILLCELL_X32 FILLER_180_1479 ();
 FILLCELL_X32 FILLER_180_1511 ();
 FILLCELL_X32 FILLER_180_1543 ();
 FILLCELL_X32 FILLER_180_1575 ();
 FILLCELL_X32 FILLER_180_1607 ();
 FILLCELL_X8 FILLER_180_1639 ();
 FILLCELL_X4 FILLER_180_1647 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X16 FILLER_181_97 ();
 FILLCELL_X8 FILLER_181_113 ();
 FILLCELL_X4 FILLER_181_121 ();
 FILLCELL_X2 FILLER_181_145 ();
 FILLCELL_X1 FILLER_181_147 ();
 FILLCELL_X16 FILLER_181_186 ();
 FILLCELL_X1 FILLER_181_202 ();
 FILLCELL_X4 FILLER_181_223 ();
 FILLCELL_X8 FILLER_181_261 ();
 FILLCELL_X1 FILLER_181_269 ();
 FILLCELL_X8 FILLER_181_307 ();
 FILLCELL_X2 FILLER_181_315 ();
 FILLCELL_X8 FILLER_181_321 ();
 FILLCELL_X4 FILLER_181_364 ();
 FILLCELL_X2 FILLER_181_368 ();
 FILLCELL_X4 FILLER_181_383 ();
 FILLCELL_X2 FILLER_181_387 ();
 FILLCELL_X4 FILLER_181_396 ();
 FILLCELL_X2 FILLER_181_400 ();
 FILLCELL_X16 FILLER_181_416 ();
 FILLCELL_X1 FILLER_181_475 ();
 FILLCELL_X1 FILLER_181_509 ();
 FILLCELL_X2 FILLER_181_512 ();
 FILLCELL_X1 FILLER_181_514 ();
 FILLCELL_X4 FILLER_181_532 ();
 FILLCELL_X2 FILLER_181_536 ();
 FILLCELL_X1 FILLER_181_542 ();
 FILLCELL_X4 FILLER_181_602 ();
 FILLCELL_X2 FILLER_181_606 ();
 FILLCELL_X4 FILLER_181_617 ();
 FILLCELL_X1 FILLER_181_621 ();
 FILLCELL_X1 FILLER_181_631 ();
 FILLCELL_X8 FILLER_181_634 ();
 FILLCELL_X2 FILLER_181_649 ();
 FILLCELL_X1 FILLER_181_651 ();
 FILLCELL_X8 FILLER_181_666 ();
 FILLCELL_X2 FILLER_181_674 ();
 FILLCELL_X16 FILLER_181_709 ();
 FILLCELL_X2 FILLER_181_725 ();
 FILLCELL_X1 FILLER_181_727 ();
 FILLCELL_X1 FILLER_181_771 ();
 FILLCELL_X2 FILLER_181_781 ();
 FILLCELL_X1 FILLER_181_783 ();
 FILLCELL_X1 FILLER_181_849 ();
 FILLCELL_X8 FILLER_181_903 ();
 FILLCELL_X2 FILLER_181_911 ();
 FILLCELL_X1 FILLER_181_913 ();
 FILLCELL_X16 FILLER_181_941 ();
 FILLCELL_X8 FILLER_181_957 ();
 FILLCELL_X1 FILLER_181_965 ();
 FILLCELL_X8 FILLER_181_970 ();
 FILLCELL_X1 FILLER_181_978 ();
 FILLCELL_X2 FILLER_181_1013 ();
 FILLCELL_X8 FILLER_181_1022 ();
 FILLCELL_X32 FILLER_181_1039 ();
 FILLCELL_X32 FILLER_181_1071 ();
 FILLCELL_X32 FILLER_181_1103 ();
 FILLCELL_X32 FILLER_181_1135 ();
 FILLCELL_X32 FILLER_181_1167 ();
 FILLCELL_X32 FILLER_181_1199 ();
 FILLCELL_X32 FILLER_181_1231 ();
 FILLCELL_X32 FILLER_181_1264 ();
 FILLCELL_X32 FILLER_181_1296 ();
 FILLCELL_X32 FILLER_181_1328 ();
 FILLCELL_X32 FILLER_181_1360 ();
 FILLCELL_X32 FILLER_181_1392 ();
 FILLCELL_X32 FILLER_181_1424 ();
 FILLCELL_X32 FILLER_181_1456 ();
 FILLCELL_X32 FILLER_181_1488 ();
 FILLCELL_X32 FILLER_181_1520 ();
 FILLCELL_X32 FILLER_181_1552 ();
 FILLCELL_X32 FILLER_181_1584 ();
 FILLCELL_X32 FILLER_181_1616 ();
 FILLCELL_X2 FILLER_181_1648 ();
 FILLCELL_X1 FILLER_181_1650 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X16 FILLER_182_97 ();
 FILLCELL_X8 FILLER_182_113 ();
 FILLCELL_X4 FILLER_182_121 ();
 FILLCELL_X16 FILLER_182_152 ();
 FILLCELL_X4 FILLER_182_168 ();
 FILLCELL_X4 FILLER_182_199 ();
 FILLCELL_X2 FILLER_182_203 ();
 FILLCELL_X1 FILLER_182_205 ();
 FILLCELL_X2 FILLER_182_213 ();
 FILLCELL_X1 FILLER_182_240 ();
 FILLCELL_X1 FILLER_182_279 ();
 FILLCELL_X8 FILLER_182_288 ();
 FILLCELL_X4 FILLER_182_296 ();
 FILLCELL_X1 FILLER_182_300 ();
 FILLCELL_X4 FILLER_182_308 ();
 FILLCELL_X2 FILLER_182_312 ();
 FILLCELL_X2 FILLER_182_341 ();
 FILLCELL_X8 FILLER_182_355 ();
 FILLCELL_X2 FILLER_182_363 ();
 FILLCELL_X1 FILLER_182_365 ();
 FILLCELL_X8 FILLER_182_378 ();
 FILLCELL_X4 FILLER_182_386 ();
 FILLCELL_X2 FILLER_182_390 ();
 FILLCELL_X2 FILLER_182_419 ();
 FILLCELL_X4 FILLER_182_428 ();
 FILLCELL_X1 FILLER_182_432 ();
 FILLCELL_X4 FILLER_182_440 ();
 FILLCELL_X1 FILLER_182_444 ();
 FILLCELL_X1 FILLER_182_456 ();
 FILLCELL_X2 FILLER_182_479 ();
 FILLCELL_X8 FILLER_182_526 ();
 FILLCELL_X4 FILLER_182_552 ();
 FILLCELL_X2 FILLER_182_567 ();
 FILLCELL_X4 FILLER_182_578 ();
 FILLCELL_X1 FILLER_182_606 ();
 FILLCELL_X2 FILLER_182_628 ();
 FILLCELL_X1 FILLER_182_630 ();
 FILLCELL_X1 FILLER_182_632 ();
 FILLCELL_X16 FILLER_182_657 ();
 FILLCELL_X4 FILLER_182_680 ();
 FILLCELL_X1 FILLER_182_684 ();
 FILLCELL_X8 FILLER_182_719 ();
 FILLCELL_X1 FILLER_182_734 ();
 FILLCELL_X2 FILLER_182_744 ();
 FILLCELL_X1 FILLER_182_773 ();
 FILLCELL_X1 FILLER_182_794 ();
 FILLCELL_X1 FILLER_182_802 ();
 FILLCELL_X2 FILLER_182_820 ();
 FILLCELL_X8 FILLER_182_825 ();
 FILLCELL_X2 FILLER_182_833 ();
 FILLCELL_X1 FILLER_182_835 ();
 FILLCELL_X4 FILLER_182_863 ();
 FILLCELL_X1 FILLER_182_895 ();
 FILLCELL_X4 FILLER_182_923 ();
 FILLCELL_X16 FILLER_182_947 ();
 FILLCELL_X8 FILLER_182_968 ();
 FILLCELL_X4 FILLER_182_976 ();
 FILLCELL_X2 FILLER_182_987 ();
 FILLCELL_X4 FILLER_182_994 ();
 FILLCELL_X16 FILLER_182_1003 ();
 FILLCELL_X32 FILLER_182_1039 ();
 FILLCELL_X32 FILLER_182_1071 ();
 FILLCELL_X32 FILLER_182_1103 ();
 FILLCELL_X32 FILLER_182_1135 ();
 FILLCELL_X32 FILLER_182_1167 ();
 FILLCELL_X32 FILLER_182_1199 ();
 FILLCELL_X32 FILLER_182_1231 ();
 FILLCELL_X32 FILLER_182_1263 ();
 FILLCELL_X32 FILLER_182_1295 ();
 FILLCELL_X32 FILLER_182_1327 ();
 FILLCELL_X32 FILLER_182_1359 ();
 FILLCELL_X32 FILLER_182_1391 ();
 FILLCELL_X32 FILLER_182_1423 ();
 FILLCELL_X32 FILLER_182_1455 ();
 FILLCELL_X32 FILLER_182_1487 ();
 FILLCELL_X32 FILLER_182_1519 ();
 FILLCELL_X32 FILLER_182_1551 ();
 FILLCELL_X32 FILLER_182_1583 ();
 FILLCELL_X32 FILLER_182_1615 ();
 FILLCELL_X4 FILLER_182_1647 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X8 FILLER_183_129 ();
 FILLCELL_X4 FILLER_183_137 ();
 FILLCELL_X2 FILLER_183_141 ();
 FILLCELL_X1 FILLER_183_143 ();
 FILLCELL_X8 FILLER_183_151 ();
 FILLCELL_X4 FILLER_183_159 ();
 FILLCELL_X1 FILLER_183_163 ();
 FILLCELL_X2 FILLER_183_191 ();
 FILLCELL_X4 FILLER_183_220 ();
 FILLCELL_X2 FILLER_183_224 ();
 FILLCELL_X1 FILLER_183_311 ();
 FILLCELL_X8 FILLER_183_344 ();
 FILLCELL_X2 FILLER_183_404 ();
 FILLCELL_X2 FILLER_183_434 ();
 FILLCELL_X4 FILLER_183_456 ();
 FILLCELL_X2 FILLER_183_460 ();
 FILLCELL_X1 FILLER_183_475 ();
 FILLCELL_X4 FILLER_183_478 ();
 FILLCELL_X2 FILLER_183_482 ();
 FILLCELL_X4 FILLER_183_489 ();
 FILLCELL_X1 FILLER_183_493 ();
 FILLCELL_X16 FILLER_183_503 ();
 FILLCELL_X4 FILLER_183_519 ();
 FILLCELL_X2 FILLER_183_523 ();
 FILLCELL_X2 FILLER_183_534 ();
 FILLCELL_X1 FILLER_183_536 ();
 FILLCELL_X4 FILLER_183_546 ();
 FILLCELL_X4 FILLER_183_559 ();
 FILLCELL_X2 FILLER_183_563 ();
 FILLCELL_X1 FILLER_183_565 ();
 FILLCELL_X8 FILLER_183_589 ();
 FILLCELL_X2 FILLER_183_597 ();
 FILLCELL_X2 FILLER_183_617 ();
 FILLCELL_X1 FILLER_183_619 ();
 FILLCELL_X4 FILLER_183_628 ();
 FILLCELL_X8 FILLER_183_650 ();
 FILLCELL_X4 FILLER_183_677 ();
 FILLCELL_X2 FILLER_183_681 ();
 FILLCELL_X1 FILLER_183_683 ();
 FILLCELL_X16 FILLER_183_691 ();
 FILLCELL_X4 FILLER_183_707 ();
 FILLCELL_X1 FILLER_183_711 ();
 FILLCELL_X1 FILLER_183_735 ();
 FILLCELL_X8 FILLER_183_752 ();
 FILLCELL_X4 FILLER_183_760 ();
 FILLCELL_X1 FILLER_183_771 ();
 FILLCELL_X2 FILLER_183_802 ();
 FILLCELL_X8 FILLER_183_859 ();
 FILLCELL_X1 FILLER_183_867 ();
 FILLCELL_X2 FILLER_183_896 ();
 FILLCELL_X4 FILLER_183_909 ();
 FILLCELL_X2 FILLER_183_913 ();
 FILLCELL_X2 FILLER_183_922 ();
 FILLCELL_X1 FILLER_183_931 ();
 FILLCELL_X2 FILLER_183_968 ();
 FILLCELL_X1 FILLER_183_990 ();
 FILLCELL_X2 FILLER_183_1018 ();
 FILLCELL_X1 FILLER_183_1020 ();
 FILLCELL_X32 FILLER_183_1048 ();
 FILLCELL_X32 FILLER_183_1080 ();
 FILLCELL_X32 FILLER_183_1112 ();
 FILLCELL_X32 FILLER_183_1144 ();
 FILLCELL_X32 FILLER_183_1176 ();
 FILLCELL_X32 FILLER_183_1208 ();
 FILLCELL_X16 FILLER_183_1240 ();
 FILLCELL_X4 FILLER_183_1256 ();
 FILLCELL_X2 FILLER_183_1260 ();
 FILLCELL_X1 FILLER_183_1262 ();
 FILLCELL_X32 FILLER_183_1264 ();
 FILLCELL_X32 FILLER_183_1296 ();
 FILLCELL_X32 FILLER_183_1328 ();
 FILLCELL_X32 FILLER_183_1360 ();
 FILLCELL_X32 FILLER_183_1392 ();
 FILLCELL_X32 FILLER_183_1424 ();
 FILLCELL_X32 FILLER_183_1456 ();
 FILLCELL_X32 FILLER_183_1488 ();
 FILLCELL_X32 FILLER_183_1520 ();
 FILLCELL_X32 FILLER_183_1552 ();
 FILLCELL_X32 FILLER_183_1584 ();
 FILLCELL_X32 FILLER_183_1616 ();
 FILLCELL_X2 FILLER_183_1648 ();
 FILLCELL_X1 FILLER_183_1650 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X8 FILLER_184_129 ();
 FILLCELL_X4 FILLER_184_137 ();
 FILLCELL_X1 FILLER_184_141 ();
 FILLCELL_X4 FILLER_184_192 ();
 FILLCELL_X4 FILLER_184_223 ();
 FILLCELL_X1 FILLER_184_227 ();
 FILLCELL_X8 FILLER_184_256 ();
 FILLCELL_X1 FILLER_184_264 ();
 FILLCELL_X2 FILLER_184_290 ();
 FILLCELL_X1 FILLER_184_292 ();
 FILLCELL_X4 FILLER_184_323 ();
 FILLCELL_X2 FILLER_184_327 ();
 FILLCELL_X2 FILLER_184_334 ();
 FILLCELL_X16 FILLER_184_352 ();
 FILLCELL_X1 FILLER_184_368 ();
 FILLCELL_X2 FILLER_184_437 ();
 FILLCELL_X4 FILLER_184_448 ();
 FILLCELL_X2 FILLER_184_452 ();
 FILLCELL_X1 FILLER_184_454 ();
 FILLCELL_X1 FILLER_184_462 ();
 FILLCELL_X8 FILLER_184_485 ();
 FILLCELL_X1 FILLER_184_496 ();
 FILLCELL_X1 FILLER_184_501 ();
 FILLCELL_X2 FILLER_184_509 ();
 FILLCELL_X8 FILLER_184_515 ();
 FILLCELL_X2 FILLER_184_523 ();
 FILLCELL_X8 FILLER_184_545 ();
 FILLCELL_X1 FILLER_184_562 ();
 FILLCELL_X1 FILLER_184_566 ();
 FILLCELL_X1 FILLER_184_571 ();
 FILLCELL_X1 FILLER_184_575 ();
 FILLCELL_X4 FILLER_184_600 ();
 FILLCELL_X2 FILLER_184_621 ();
 FILLCELL_X2 FILLER_184_625 ();
 FILLCELL_X1 FILLER_184_630 ();
 FILLCELL_X4 FILLER_184_657 ();
 FILLCELL_X1 FILLER_184_661 ();
 FILLCELL_X16 FILLER_184_674 ();
 FILLCELL_X4 FILLER_184_690 ();
 FILLCELL_X4 FILLER_184_701 ();
 FILLCELL_X2 FILLER_184_705 ();
 FILLCELL_X1 FILLER_184_707 ();
 FILLCELL_X2 FILLER_184_721 ();
 FILLCELL_X1 FILLER_184_723 ();
 FILLCELL_X4 FILLER_184_744 ();
 FILLCELL_X8 FILLER_184_768 ();
 FILLCELL_X4 FILLER_184_776 ();
 FILLCELL_X2 FILLER_184_780 ();
 FILLCELL_X2 FILLER_184_787 ();
 FILLCELL_X4 FILLER_184_816 ();
 FILLCELL_X2 FILLER_184_820 ();
 FILLCELL_X8 FILLER_184_862 ();
 FILLCELL_X8 FILLER_184_896 ();
 FILLCELL_X2 FILLER_184_904 ();
 FILLCELL_X4 FILLER_184_926 ();
 FILLCELL_X1 FILLER_184_930 ();
 FILLCELL_X2 FILLER_184_938 ();
 FILLCELL_X4 FILLER_184_967 ();
 FILLCELL_X8 FILLER_184_1001 ();
 FILLCELL_X2 FILLER_184_1009 ();
 FILLCELL_X2 FILLER_184_1023 ();
 FILLCELL_X1 FILLER_184_1025 ();
 FILLCELL_X4 FILLER_184_1037 ();
 FILLCELL_X32 FILLER_184_1054 ();
 FILLCELL_X32 FILLER_184_1086 ();
 FILLCELL_X32 FILLER_184_1118 ();
 FILLCELL_X32 FILLER_184_1150 ();
 FILLCELL_X32 FILLER_184_1182 ();
 FILLCELL_X32 FILLER_184_1214 ();
 FILLCELL_X32 FILLER_184_1246 ();
 FILLCELL_X32 FILLER_184_1278 ();
 FILLCELL_X32 FILLER_184_1310 ();
 FILLCELL_X32 FILLER_184_1342 ();
 FILLCELL_X32 FILLER_184_1374 ();
 FILLCELL_X32 FILLER_184_1406 ();
 FILLCELL_X32 FILLER_184_1438 ();
 FILLCELL_X32 FILLER_184_1470 ();
 FILLCELL_X32 FILLER_184_1502 ();
 FILLCELL_X32 FILLER_184_1534 ();
 FILLCELL_X32 FILLER_184_1566 ();
 FILLCELL_X32 FILLER_184_1598 ();
 FILLCELL_X16 FILLER_184_1630 ();
 FILLCELL_X4 FILLER_184_1646 ();
 FILLCELL_X1 FILLER_184_1650 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X16 FILLER_185_129 ();
 FILLCELL_X2 FILLER_185_145 ();
 FILLCELL_X1 FILLER_185_147 ();
 FILLCELL_X8 FILLER_185_153 ();
 FILLCELL_X4 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_185 ();
 FILLCELL_X4 FILLER_185_217 ();
 FILLCELL_X2 FILLER_185_221 ();
 FILLCELL_X1 FILLER_185_243 ();
 FILLCELL_X8 FILLER_185_269 ();
 FILLCELL_X4 FILLER_185_277 ();
 FILLCELL_X8 FILLER_185_290 ();
 FILLCELL_X1 FILLER_185_305 ();
 FILLCELL_X1 FILLER_185_326 ();
 FILLCELL_X1 FILLER_185_347 ();
 FILLCELL_X1 FILLER_185_355 ();
 FILLCELL_X4 FILLER_185_368 ();
 FILLCELL_X2 FILLER_185_386 ();
 FILLCELL_X4 FILLER_185_440 ();
 FILLCELL_X2 FILLER_185_448 ();
 FILLCELL_X1 FILLER_185_450 ();
 FILLCELL_X2 FILLER_185_471 ();
 FILLCELL_X4 FILLER_185_483 ();
 FILLCELL_X1 FILLER_185_487 ();
 FILLCELL_X8 FILLER_185_516 ();
 FILLCELL_X1 FILLER_185_524 ();
 FILLCELL_X1 FILLER_185_529 ();
 FILLCELL_X8 FILLER_185_542 ();
 FILLCELL_X4 FILLER_185_550 ();
 FILLCELL_X8 FILLER_185_602 ();
 FILLCELL_X8 FILLER_185_623 ();
 FILLCELL_X4 FILLER_185_631 ();
 FILLCELL_X2 FILLER_185_635 ();
 FILLCELL_X4 FILLER_185_665 ();
 FILLCELL_X2 FILLER_185_669 ();
 FILLCELL_X2 FILLER_185_685 ();
 FILLCELL_X1 FILLER_185_687 ();
 FILLCELL_X2 FILLER_185_695 ();
 FILLCELL_X1 FILLER_185_697 ();
 FILLCELL_X4 FILLER_185_742 ();
 FILLCELL_X1 FILLER_185_764 ();
 FILLCELL_X8 FILLER_185_785 ();
 FILLCELL_X1 FILLER_185_800 ();
 FILLCELL_X8 FILLER_185_819 ();
 FILLCELL_X4 FILLER_185_827 ();
 FILLCELL_X2 FILLER_185_871 ();
 FILLCELL_X4 FILLER_185_886 ();
 FILLCELL_X32 FILLER_185_924 ();
 FILLCELL_X8 FILLER_185_956 ();
 FILLCELL_X4 FILLER_185_964 ();
 FILLCELL_X2 FILLER_185_968 ();
 FILLCELL_X8 FILLER_185_988 ();
 FILLCELL_X4 FILLER_185_996 ();
 FILLCELL_X1 FILLER_185_1000 ();
 FILLCELL_X4 FILLER_185_1008 ();
 FILLCELL_X1 FILLER_185_1012 ();
 FILLCELL_X8 FILLER_185_1033 ();
 FILLCELL_X4 FILLER_185_1041 ();
 FILLCELL_X1 FILLER_185_1045 ();
 FILLCELL_X32 FILLER_185_1059 ();
 FILLCELL_X32 FILLER_185_1091 ();
 FILLCELL_X32 FILLER_185_1123 ();
 FILLCELL_X32 FILLER_185_1155 ();
 FILLCELL_X32 FILLER_185_1187 ();
 FILLCELL_X32 FILLER_185_1219 ();
 FILLCELL_X8 FILLER_185_1251 ();
 FILLCELL_X4 FILLER_185_1259 ();
 FILLCELL_X32 FILLER_185_1264 ();
 FILLCELL_X32 FILLER_185_1296 ();
 FILLCELL_X32 FILLER_185_1328 ();
 FILLCELL_X32 FILLER_185_1360 ();
 FILLCELL_X32 FILLER_185_1392 ();
 FILLCELL_X32 FILLER_185_1424 ();
 FILLCELL_X32 FILLER_185_1456 ();
 FILLCELL_X32 FILLER_185_1488 ();
 FILLCELL_X32 FILLER_185_1520 ();
 FILLCELL_X32 FILLER_185_1552 ();
 FILLCELL_X32 FILLER_185_1584 ();
 FILLCELL_X32 FILLER_185_1616 ();
 FILLCELL_X2 FILLER_185_1648 ();
 FILLCELL_X1 FILLER_185_1650 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X4 FILLER_186_161 ();
 FILLCELL_X2 FILLER_186_165 ();
 FILLCELL_X16 FILLER_186_190 ();
 FILLCELL_X2 FILLER_186_206 ();
 FILLCELL_X1 FILLER_186_208 ();
 FILLCELL_X8 FILLER_186_265 ();
 FILLCELL_X4 FILLER_186_293 ();
 FILLCELL_X2 FILLER_186_322 ();
 FILLCELL_X1 FILLER_186_324 ();
 FILLCELL_X1 FILLER_186_372 ();
 FILLCELL_X4 FILLER_186_384 ();
 FILLCELL_X1 FILLER_186_388 ();
 FILLCELL_X2 FILLER_186_391 ();
 FILLCELL_X1 FILLER_186_393 ();
 FILLCELL_X1 FILLER_186_405 ();
 FILLCELL_X4 FILLER_186_410 ();
 FILLCELL_X1 FILLER_186_414 ();
 FILLCELL_X16 FILLER_186_419 ();
 FILLCELL_X2 FILLER_186_435 ();
 FILLCELL_X1 FILLER_186_437 ();
 FILLCELL_X8 FILLER_186_447 ();
 FILLCELL_X2 FILLER_186_455 ();
 FILLCELL_X2 FILLER_186_461 ();
 FILLCELL_X2 FILLER_186_466 ();
 FILLCELL_X1 FILLER_186_475 ();
 FILLCELL_X8 FILLER_186_553 ();
 FILLCELL_X1 FILLER_186_565 ();
 FILLCELL_X4 FILLER_186_569 ();
 FILLCELL_X8 FILLER_186_593 ();
 FILLCELL_X8 FILLER_186_632 ();
 FILLCELL_X2 FILLER_186_640 ();
 FILLCELL_X1 FILLER_186_642 ();
 FILLCELL_X16 FILLER_186_659 ();
 FILLCELL_X2 FILLER_186_675 ();
 FILLCELL_X2 FILLER_186_686 ();
 FILLCELL_X4 FILLER_186_716 ();
 FILLCELL_X4 FILLER_186_745 ();
 FILLCELL_X2 FILLER_186_749 ();
 FILLCELL_X1 FILLER_186_751 ();
 FILLCELL_X4 FILLER_186_779 ();
 FILLCELL_X2 FILLER_186_783 ();
 FILLCELL_X1 FILLER_186_805 ();
 FILLCELL_X4 FILLER_186_813 ();
 FILLCELL_X1 FILLER_186_817 ();
 FILLCELL_X16 FILLER_186_845 ();
 FILLCELL_X8 FILLER_186_861 ();
 FILLCELL_X2 FILLER_186_869 ();
 FILLCELL_X1 FILLER_186_871 ();
 FILLCELL_X2 FILLER_186_908 ();
 FILLCELL_X4 FILLER_186_937 ();
 FILLCELL_X2 FILLER_186_941 ();
 FILLCELL_X1 FILLER_186_943 ();
 FILLCELL_X16 FILLER_186_949 ();
 FILLCELL_X4 FILLER_186_965 ();
 FILLCELL_X2 FILLER_186_969 ();
 FILLCELL_X4 FILLER_186_991 ();
 FILLCELL_X2 FILLER_186_995 ();
 FILLCELL_X32 FILLER_186_1037 ();
 FILLCELL_X32 FILLER_186_1069 ();
 FILLCELL_X32 FILLER_186_1101 ();
 FILLCELL_X32 FILLER_186_1133 ();
 FILLCELL_X32 FILLER_186_1165 ();
 FILLCELL_X32 FILLER_186_1197 ();
 FILLCELL_X32 FILLER_186_1229 ();
 FILLCELL_X32 FILLER_186_1261 ();
 FILLCELL_X32 FILLER_186_1293 ();
 FILLCELL_X32 FILLER_186_1325 ();
 FILLCELL_X32 FILLER_186_1357 ();
 FILLCELL_X32 FILLER_186_1389 ();
 FILLCELL_X32 FILLER_186_1421 ();
 FILLCELL_X32 FILLER_186_1453 ();
 FILLCELL_X32 FILLER_186_1485 ();
 FILLCELL_X32 FILLER_186_1517 ();
 FILLCELL_X32 FILLER_186_1549 ();
 FILLCELL_X32 FILLER_186_1581 ();
 FILLCELL_X32 FILLER_186_1613 ();
 FILLCELL_X4 FILLER_186_1645 ();
 FILLCELL_X2 FILLER_186_1649 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X8 FILLER_187_161 ();
 FILLCELL_X2 FILLER_187_169 ();
 FILLCELL_X16 FILLER_187_231 ();
 FILLCELL_X16 FILLER_187_254 ();
 FILLCELL_X2 FILLER_187_270 ();
 FILLCELL_X1 FILLER_187_272 ();
 FILLCELL_X1 FILLER_187_287 ();
 FILLCELL_X8 FILLER_187_300 ();
 FILLCELL_X4 FILLER_187_308 ();
 FILLCELL_X2 FILLER_187_312 ();
 FILLCELL_X1 FILLER_187_314 ();
 FILLCELL_X8 FILLER_187_322 ();
 FILLCELL_X4 FILLER_187_334 ();
 FILLCELL_X2 FILLER_187_345 ();
 FILLCELL_X2 FILLER_187_367 ();
 FILLCELL_X1 FILLER_187_369 ();
 FILLCELL_X4 FILLER_187_390 ();
 FILLCELL_X1 FILLER_187_394 ();
 FILLCELL_X8 FILLER_187_422 ();
 FILLCELL_X1 FILLER_187_450 ();
 FILLCELL_X16 FILLER_187_474 ();
 FILLCELL_X2 FILLER_187_490 ();
 FILLCELL_X1 FILLER_187_516 ();
 FILLCELL_X1 FILLER_187_529 ();
 FILLCELL_X1 FILLER_187_555 ();
 FILLCELL_X4 FILLER_187_576 ();
 FILLCELL_X2 FILLER_187_580 ();
 FILLCELL_X1 FILLER_187_582 ();
 FILLCELL_X8 FILLER_187_590 ();
 FILLCELL_X4 FILLER_187_598 ();
 FILLCELL_X2 FILLER_187_602 ();
 FILLCELL_X8 FILLER_187_609 ();
 FILLCELL_X8 FILLER_187_630 ();
 FILLCELL_X2 FILLER_187_638 ();
 FILLCELL_X1 FILLER_187_640 ();
 FILLCELL_X8 FILLER_187_657 ();
 FILLCELL_X1 FILLER_187_665 ();
 FILLCELL_X2 FILLER_187_700 ();
 FILLCELL_X8 FILLER_187_709 ();
 FILLCELL_X2 FILLER_187_717 ();
 FILLCELL_X2 FILLER_187_739 ();
 FILLCELL_X1 FILLER_187_741 ();
 FILLCELL_X1 FILLER_187_769 ();
 FILLCELL_X4 FILLER_187_790 ();
 FILLCELL_X4 FILLER_187_801 ();
 FILLCELL_X2 FILLER_187_805 ();
 FILLCELL_X1 FILLER_187_807 ();
 FILLCELL_X2 FILLER_187_828 ();
 FILLCELL_X1 FILLER_187_830 ();
 FILLCELL_X4 FILLER_187_838 ();
 FILLCELL_X2 FILLER_187_842 ();
 FILLCELL_X1 FILLER_187_844 ();
 FILLCELL_X2 FILLER_187_853 ();
 FILLCELL_X1 FILLER_187_855 ();
 FILLCELL_X8 FILLER_187_865 ();
 FILLCELL_X4 FILLER_187_873 ();
 FILLCELL_X1 FILLER_187_877 ();
 FILLCELL_X4 FILLER_187_905 ();
 FILLCELL_X1 FILLER_187_909 ();
 FILLCELL_X8 FILLER_187_917 ();
 FILLCELL_X2 FILLER_187_925 ();
 FILLCELL_X4 FILLER_187_957 ();
 FILLCELL_X4 FILLER_187_1002 ();
 FILLCELL_X2 FILLER_187_1006 ();
 FILLCELL_X1 FILLER_187_1015 ();
 FILLCELL_X32 FILLER_187_1028 ();
 FILLCELL_X32 FILLER_187_1060 ();
 FILLCELL_X32 FILLER_187_1092 ();
 FILLCELL_X32 FILLER_187_1124 ();
 FILLCELL_X32 FILLER_187_1156 ();
 FILLCELL_X32 FILLER_187_1188 ();
 FILLCELL_X32 FILLER_187_1220 ();
 FILLCELL_X8 FILLER_187_1252 ();
 FILLCELL_X2 FILLER_187_1260 ();
 FILLCELL_X1 FILLER_187_1262 ();
 FILLCELL_X32 FILLER_187_1264 ();
 FILLCELL_X32 FILLER_187_1296 ();
 FILLCELL_X32 FILLER_187_1328 ();
 FILLCELL_X32 FILLER_187_1360 ();
 FILLCELL_X32 FILLER_187_1392 ();
 FILLCELL_X32 FILLER_187_1424 ();
 FILLCELL_X32 FILLER_187_1456 ();
 FILLCELL_X32 FILLER_187_1488 ();
 FILLCELL_X32 FILLER_187_1520 ();
 FILLCELL_X32 FILLER_187_1552 ();
 FILLCELL_X32 FILLER_187_1584 ();
 FILLCELL_X32 FILLER_187_1616 ();
 FILLCELL_X2 FILLER_187_1648 ();
 FILLCELL_X1 FILLER_187_1650 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X16 FILLER_188_193 ();
 FILLCELL_X4 FILLER_188_209 ();
 FILLCELL_X1 FILLER_188_213 ();
 FILLCELL_X16 FILLER_188_256 ();
 FILLCELL_X4 FILLER_188_292 ();
 FILLCELL_X16 FILLER_188_302 ();
 FILLCELL_X8 FILLER_188_338 ();
 FILLCELL_X2 FILLER_188_346 ();
 FILLCELL_X8 FILLER_188_352 ();
 FILLCELL_X4 FILLER_188_360 ();
 FILLCELL_X1 FILLER_188_364 ();
 FILLCELL_X8 FILLER_188_403 ();
 FILLCELL_X8 FILLER_188_431 ();
 FILLCELL_X1 FILLER_188_439 ();
 FILLCELL_X2 FILLER_188_449 ();
 FILLCELL_X4 FILLER_188_462 ();
 FILLCELL_X2 FILLER_188_466 ();
 FILLCELL_X4 FILLER_188_492 ();
 FILLCELL_X2 FILLER_188_496 ();
 FILLCELL_X4 FILLER_188_505 ();
 FILLCELL_X2 FILLER_188_509 ();
 FILLCELL_X1 FILLER_188_511 ();
 FILLCELL_X16 FILLER_188_523 ();
 FILLCELL_X1 FILLER_188_542 ();
 FILLCELL_X2 FILLER_188_575 ();
 FILLCELL_X1 FILLER_188_577 ();
 FILLCELL_X2 FILLER_188_598 ();
 FILLCELL_X16 FILLER_188_608 ();
 FILLCELL_X4 FILLER_188_624 ();
 FILLCELL_X2 FILLER_188_628 ();
 FILLCELL_X1 FILLER_188_630 ();
 FILLCELL_X4 FILLER_188_650 ();
 FILLCELL_X2 FILLER_188_659 ();
 FILLCELL_X1 FILLER_188_661 ();
 FILLCELL_X8 FILLER_188_739 ();
 FILLCELL_X4 FILLER_188_774 ();
 FILLCELL_X4 FILLER_188_798 ();
 FILLCELL_X2 FILLER_188_802 ();
 FILLCELL_X1 FILLER_188_804 ();
 FILLCELL_X16 FILLER_188_810 ();
 FILLCELL_X4 FILLER_188_826 ();
 FILLCELL_X1 FILLER_188_830 ();
 FILLCELL_X4 FILLER_188_838 ();
 FILLCELL_X1 FILLER_188_842 ();
 FILLCELL_X1 FILLER_188_876 ();
 FILLCELL_X4 FILLER_188_891 ();
 FILLCELL_X2 FILLER_188_895 ();
 FILLCELL_X1 FILLER_188_897 ();
 FILLCELL_X1 FILLER_188_918 ();
 FILLCELL_X2 FILLER_188_944 ();
 FILLCELL_X2 FILLER_188_966 ();
 FILLCELL_X1 FILLER_188_968 ();
 FILLCELL_X8 FILLER_188_989 ();
 FILLCELL_X4 FILLER_188_997 ();
 FILLCELL_X2 FILLER_188_1001 ();
 FILLCELL_X32 FILLER_188_1023 ();
 FILLCELL_X32 FILLER_188_1055 ();
 FILLCELL_X32 FILLER_188_1087 ();
 FILLCELL_X32 FILLER_188_1119 ();
 FILLCELL_X32 FILLER_188_1151 ();
 FILLCELL_X32 FILLER_188_1183 ();
 FILLCELL_X32 FILLER_188_1215 ();
 FILLCELL_X32 FILLER_188_1247 ();
 FILLCELL_X32 FILLER_188_1279 ();
 FILLCELL_X32 FILLER_188_1311 ();
 FILLCELL_X32 FILLER_188_1343 ();
 FILLCELL_X32 FILLER_188_1375 ();
 FILLCELL_X32 FILLER_188_1407 ();
 FILLCELL_X32 FILLER_188_1439 ();
 FILLCELL_X32 FILLER_188_1471 ();
 FILLCELL_X32 FILLER_188_1503 ();
 FILLCELL_X32 FILLER_188_1535 ();
 FILLCELL_X32 FILLER_188_1567 ();
 FILLCELL_X32 FILLER_188_1599 ();
 FILLCELL_X16 FILLER_188_1631 ();
 FILLCELL_X4 FILLER_188_1647 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X8 FILLER_189_193 ();
 FILLCELL_X4 FILLER_189_201 ();
 FILLCELL_X2 FILLER_189_225 ();
 FILLCELL_X1 FILLER_189_227 ();
 FILLCELL_X4 FILLER_189_231 ();
 FILLCELL_X2 FILLER_189_235 ();
 FILLCELL_X8 FILLER_189_264 ();
 FILLCELL_X1 FILLER_189_297 ();
 FILLCELL_X4 FILLER_189_318 ();
 FILLCELL_X2 FILLER_189_322 ();
 FILLCELL_X16 FILLER_189_331 ();
 FILLCELL_X1 FILLER_189_354 ();
 FILLCELL_X1 FILLER_189_362 ();
 FILLCELL_X8 FILLER_189_374 ();
 FILLCELL_X2 FILLER_189_382 ();
 FILLCELL_X16 FILLER_189_397 ();
 FILLCELL_X1 FILLER_189_417 ();
 FILLCELL_X8 FILLER_189_422 ();
 FILLCELL_X1 FILLER_189_430 ();
 FILLCELL_X1 FILLER_189_505 ();
 FILLCELL_X2 FILLER_189_510 ();
 FILLCELL_X1 FILLER_189_515 ();
 FILLCELL_X1 FILLER_189_525 ();
 FILLCELL_X4 FILLER_189_530 ();
 FILLCELL_X1 FILLER_189_534 ();
 FILLCELL_X8 FILLER_189_545 ();
 FILLCELL_X1 FILLER_189_590 ();
 FILLCELL_X2 FILLER_189_613 ();
 FILLCELL_X1 FILLER_189_644 ();
 FILLCELL_X1 FILLER_189_677 ();
 FILLCELL_X16 FILLER_189_706 ();
 FILLCELL_X4 FILLER_189_722 ();
 FILLCELL_X1 FILLER_189_726 ();
 FILLCELL_X4 FILLER_189_729 ();
 FILLCELL_X1 FILLER_189_733 ();
 FILLCELL_X16 FILLER_189_737 ();
 FILLCELL_X2 FILLER_189_753 ();
 FILLCELL_X1 FILLER_189_755 ();
 FILLCELL_X16 FILLER_189_781 ();
 FILLCELL_X2 FILLER_189_797 ();
 FILLCELL_X1 FILLER_189_799 ();
 FILLCELL_X16 FILLER_189_818 ();
 FILLCELL_X2 FILLER_189_842 ();
 FILLCELL_X4 FILLER_189_848 ();
 FILLCELL_X8 FILLER_189_876 ();
 FILLCELL_X16 FILLER_189_904 ();
 FILLCELL_X2 FILLER_189_920 ();
 FILLCELL_X4 FILLER_189_924 ();
 FILLCELL_X32 FILLER_189_939 ();
 FILLCELL_X32 FILLER_189_971 ();
 FILLCELL_X32 FILLER_189_1003 ();
 FILLCELL_X32 FILLER_189_1035 ();
 FILLCELL_X32 FILLER_189_1067 ();
 FILLCELL_X32 FILLER_189_1099 ();
 FILLCELL_X32 FILLER_189_1131 ();
 FILLCELL_X32 FILLER_189_1163 ();
 FILLCELL_X32 FILLER_189_1195 ();
 FILLCELL_X32 FILLER_189_1227 ();
 FILLCELL_X4 FILLER_189_1259 ();
 FILLCELL_X32 FILLER_189_1264 ();
 FILLCELL_X32 FILLER_189_1296 ();
 FILLCELL_X32 FILLER_189_1328 ();
 FILLCELL_X32 FILLER_189_1360 ();
 FILLCELL_X32 FILLER_189_1392 ();
 FILLCELL_X32 FILLER_189_1424 ();
 FILLCELL_X32 FILLER_189_1456 ();
 FILLCELL_X32 FILLER_189_1488 ();
 FILLCELL_X32 FILLER_189_1520 ();
 FILLCELL_X32 FILLER_189_1552 ();
 FILLCELL_X32 FILLER_189_1584 ();
 FILLCELL_X32 FILLER_189_1616 ();
 FILLCELL_X2 FILLER_189_1648 ();
 FILLCELL_X1 FILLER_189_1650 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X16 FILLER_190_193 ();
 FILLCELL_X1 FILLER_190_209 ();
 FILLCELL_X8 FILLER_190_237 ();
 FILLCELL_X4 FILLER_190_245 ();
 FILLCELL_X1 FILLER_190_269 ();
 FILLCELL_X4 FILLER_190_279 ();
 FILLCELL_X8 FILLER_190_310 ();
 FILLCELL_X2 FILLER_190_318 ();
 FILLCELL_X1 FILLER_190_320 ();
 FILLCELL_X4 FILLER_190_341 ();
 FILLCELL_X1 FILLER_190_349 ();
 FILLCELL_X8 FILLER_190_370 ();
 FILLCELL_X1 FILLER_190_378 ();
 FILLCELL_X1 FILLER_190_387 ();
 FILLCELL_X4 FILLER_190_426 ();
 FILLCELL_X2 FILLER_190_430 ();
 FILLCELL_X1 FILLER_190_432 ();
 FILLCELL_X8 FILLER_190_449 ();
 FILLCELL_X4 FILLER_190_457 ();
 FILLCELL_X1 FILLER_190_461 ();
 FILLCELL_X4 FILLER_190_465 ();
 FILLCELL_X4 FILLER_190_473 ();
 FILLCELL_X2 FILLER_190_477 ();
 FILLCELL_X1 FILLER_190_479 ();
 FILLCELL_X1 FILLER_190_499 ();
 FILLCELL_X2 FILLER_190_520 ();
 FILLCELL_X1 FILLER_190_522 ();
 FILLCELL_X4 FILLER_190_546 ();
 FILLCELL_X2 FILLER_190_555 ();
 FILLCELL_X1 FILLER_190_597 ();
 FILLCELL_X1 FILLER_190_603 ();
 FILLCELL_X8 FILLER_190_639 ();
 FILLCELL_X4 FILLER_190_647 ();
 FILLCELL_X2 FILLER_190_651 ();
 FILLCELL_X1 FILLER_190_653 ();
 FILLCELL_X4 FILLER_190_694 ();
 FILLCELL_X2 FILLER_190_698 ();
 FILLCELL_X2 FILLER_190_757 ();
 FILLCELL_X1 FILLER_190_759 ();
 FILLCELL_X1 FILLER_190_772 ();
 FILLCELL_X4 FILLER_190_804 ();
 FILLCELL_X2 FILLER_190_808 ();
 FILLCELL_X2 FILLER_190_856 ();
 FILLCELL_X4 FILLER_190_865 ();
 FILLCELL_X1 FILLER_190_869 ();
 FILLCELL_X4 FILLER_190_894 ();
 FILLCELL_X1 FILLER_190_905 ();
 FILLCELL_X2 FILLER_190_926 ();
 FILLCELL_X32 FILLER_190_955 ();
 FILLCELL_X32 FILLER_190_987 ();
 FILLCELL_X32 FILLER_190_1019 ();
 FILLCELL_X32 FILLER_190_1051 ();
 FILLCELL_X32 FILLER_190_1083 ();
 FILLCELL_X32 FILLER_190_1115 ();
 FILLCELL_X32 FILLER_190_1147 ();
 FILLCELL_X32 FILLER_190_1179 ();
 FILLCELL_X32 FILLER_190_1211 ();
 FILLCELL_X32 FILLER_190_1243 ();
 FILLCELL_X32 FILLER_190_1275 ();
 FILLCELL_X32 FILLER_190_1307 ();
 FILLCELL_X32 FILLER_190_1339 ();
 FILLCELL_X32 FILLER_190_1371 ();
 FILLCELL_X32 FILLER_190_1403 ();
 FILLCELL_X32 FILLER_190_1435 ();
 FILLCELL_X32 FILLER_190_1467 ();
 FILLCELL_X32 FILLER_190_1499 ();
 FILLCELL_X32 FILLER_190_1531 ();
 FILLCELL_X32 FILLER_190_1563 ();
 FILLCELL_X32 FILLER_190_1595 ();
 FILLCELL_X16 FILLER_190_1627 ();
 FILLCELL_X8 FILLER_190_1643 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X16 FILLER_191_193 ();
 FILLCELL_X8 FILLER_191_209 ();
 FILLCELL_X16 FILLER_191_229 ();
 FILLCELL_X8 FILLER_191_245 ();
 FILLCELL_X4 FILLER_191_267 ();
 FILLCELL_X2 FILLER_191_271 ();
 FILLCELL_X8 FILLER_191_353 ();
 FILLCELL_X4 FILLER_191_361 ();
 FILLCELL_X2 FILLER_191_365 ();
 FILLCELL_X2 FILLER_191_421 ();
 FILLCELL_X1 FILLER_191_423 ();
 FILLCELL_X2 FILLER_191_458 ();
 FILLCELL_X1 FILLER_191_471 ();
 FILLCELL_X8 FILLER_191_479 ();
 FILLCELL_X4 FILLER_191_487 ();
 FILLCELL_X1 FILLER_191_491 ();
 FILLCELL_X2 FILLER_191_496 ();
 FILLCELL_X1 FILLER_191_498 ();
 FILLCELL_X16 FILLER_191_502 ();
 FILLCELL_X8 FILLER_191_518 ();
 FILLCELL_X2 FILLER_191_526 ();
 FILLCELL_X1 FILLER_191_528 ();
 FILLCELL_X2 FILLER_191_538 ();
 FILLCELL_X2 FILLER_191_571 ();
 FILLCELL_X1 FILLER_191_573 ();
 FILLCELL_X1 FILLER_191_577 ();
 FILLCELL_X8 FILLER_191_585 ();
 FILLCELL_X2 FILLER_191_593 ();
 FILLCELL_X1 FILLER_191_595 ();
 FILLCELL_X4 FILLER_191_614 ();
 FILLCELL_X2 FILLER_191_618 ();
 FILLCELL_X1 FILLER_191_620 ();
 FILLCELL_X2 FILLER_191_643 ();
 FILLCELL_X4 FILLER_191_651 ();
 FILLCELL_X2 FILLER_191_655 ();
 FILLCELL_X1 FILLER_191_657 ();
 FILLCELL_X4 FILLER_191_665 ();
 FILLCELL_X2 FILLER_191_669 ();
 FILLCELL_X1 FILLER_191_671 ();
 FILLCELL_X2 FILLER_191_690 ();
 FILLCELL_X1 FILLER_191_692 ();
 FILLCELL_X8 FILLER_191_700 ();
 FILLCELL_X4 FILLER_191_708 ();
 FILLCELL_X2 FILLER_191_719 ();
 FILLCELL_X1 FILLER_191_775 ();
 FILLCELL_X16 FILLER_191_783 ();
 FILLCELL_X1 FILLER_191_806 ();
 FILLCELL_X8 FILLER_191_818 ();
 FILLCELL_X2 FILLER_191_826 ();
 FILLCELL_X8 FILLER_191_864 ();
 FILLCELL_X1 FILLER_191_872 ();
 FILLCELL_X4 FILLER_191_885 ();
 FILLCELL_X1 FILLER_191_889 ();
 FILLCELL_X2 FILLER_191_917 ();
 FILLCELL_X4 FILLER_191_926 ();
 FILLCELL_X1 FILLER_191_930 ();
 FILLCELL_X32 FILLER_191_960 ();
 FILLCELL_X32 FILLER_191_992 ();
 FILLCELL_X32 FILLER_191_1024 ();
 FILLCELL_X32 FILLER_191_1056 ();
 FILLCELL_X32 FILLER_191_1088 ();
 FILLCELL_X32 FILLER_191_1120 ();
 FILLCELL_X32 FILLER_191_1152 ();
 FILLCELL_X32 FILLER_191_1184 ();
 FILLCELL_X32 FILLER_191_1216 ();
 FILLCELL_X8 FILLER_191_1248 ();
 FILLCELL_X4 FILLER_191_1256 ();
 FILLCELL_X2 FILLER_191_1260 ();
 FILLCELL_X1 FILLER_191_1262 ();
 FILLCELL_X32 FILLER_191_1264 ();
 FILLCELL_X32 FILLER_191_1296 ();
 FILLCELL_X32 FILLER_191_1328 ();
 FILLCELL_X32 FILLER_191_1360 ();
 FILLCELL_X32 FILLER_191_1392 ();
 FILLCELL_X32 FILLER_191_1424 ();
 FILLCELL_X32 FILLER_191_1456 ();
 FILLCELL_X32 FILLER_191_1488 ();
 FILLCELL_X32 FILLER_191_1520 ();
 FILLCELL_X32 FILLER_191_1552 ();
 FILLCELL_X32 FILLER_191_1584 ();
 FILLCELL_X32 FILLER_191_1616 ();
 FILLCELL_X2 FILLER_191_1648 ();
 FILLCELL_X1 FILLER_191_1650 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X16 FILLER_192_225 ();
 FILLCELL_X8 FILLER_192_241 ();
 FILLCELL_X4 FILLER_192_249 ();
 FILLCELL_X2 FILLER_192_253 ();
 FILLCELL_X1 FILLER_192_305 ();
 FILLCELL_X2 FILLER_192_313 ();
 FILLCELL_X1 FILLER_192_315 ();
 FILLCELL_X2 FILLER_192_323 ();
 FILLCELL_X1 FILLER_192_325 ();
 FILLCELL_X2 FILLER_192_365 ();
 FILLCELL_X1 FILLER_192_367 ();
 FILLCELL_X4 FILLER_192_403 ();
 FILLCELL_X2 FILLER_192_407 ();
 FILLCELL_X1 FILLER_192_409 ();
 FILLCELL_X16 FILLER_192_414 ();
 FILLCELL_X2 FILLER_192_430 ();
 FILLCELL_X1 FILLER_192_432 ();
 FILLCELL_X2 FILLER_192_442 ();
 FILLCELL_X2 FILLER_192_487 ();
 FILLCELL_X1 FILLER_192_489 ();
 FILLCELL_X2 FILLER_192_510 ();
 FILLCELL_X1 FILLER_192_528 ();
 FILLCELL_X2 FILLER_192_549 ();
 FILLCELL_X1 FILLER_192_555 ();
 FILLCELL_X2 FILLER_192_559 ();
 FILLCELL_X16 FILLER_192_568 ();
 FILLCELL_X1 FILLER_192_632 ();
 FILLCELL_X1 FILLER_192_642 ();
 FILLCELL_X1 FILLER_192_650 ();
 FILLCELL_X1 FILLER_192_671 ();
 FILLCELL_X16 FILLER_192_697 ();
 FILLCELL_X8 FILLER_192_713 ();
 FILLCELL_X4 FILLER_192_748 ();
 FILLCELL_X2 FILLER_192_752 ();
 FILLCELL_X1 FILLER_192_754 ();
 FILLCELL_X2 FILLER_192_759 ();
 FILLCELL_X8 FILLER_192_768 ();
 FILLCELL_X1 FILLER_192_776 ();
 FILLCELL_X32 FILLER_192_817 ();
 FILLCELL_X2 FILLER_192_849 ();
 FILLCELL_X4 FILLER_192_864 ();
 FILLCELL_X2 FILLER_192_868 ();
 FILLCELL_X1 FILLER_192_870 ();
 FILLCELL_X4 FILLER_192_880 ();
 FILLCELL_X2 FILLER_192_884 ();
 FILLCELL_X1 FILLER_192_886 ();
 FILLCELL_X2 FILLER_192_894 ();
 FILLCELL_X1 FILLER_192_896 ();
 FILLCELL_X8 FILLER_192_922 ();
 FILLCELL_X32 FILLER_192_957 ();
 FILLCELL_X32 FILLER_192_989 ();
 FILLCELL_X32 FILLER_192_1021 ();
 FILLCELL_X32 FILLER_192_1053 ();
 FILLCELL_X32 FILLER_192_1085 ();
 FILLCELL_X32 FILLER_192_1117 ();
 FILLCELL_X32 FILLER_192_1149 ();
 FILLCELL_X32 FILLER_192_1181 ();
 FILLCELL_X32 FILLER_192_1213 ();
 FILLCELL_X32 FILLER_192_1245 ();
 FILLCELL_X32 FILLER_192_1277 ();
 FILLCELL_X32 FILLER_192_1309 ();
 FILLCELL_X32 FILLER_192_1341 ();
 FILLCELL_X32 FILLER_192_1373 ();
 FILLCELL_X32 FILLER_192_1405 ();
 FILLCELL_X32 FILLER_192_1437 ();
 FILLCELL_X32 FILLER_192_1469 ();
 FILLCELL_X32 FILLER_192_1501 ();
 FILLCELL_X32 FILLER_192_1533 ();
 FILLCELL_X32 FILLER_192_1565 ();
 FILLCELL_X32 FILLER_192_1597 ();
 FILLCELL_X16 FILLER_192_1629 ();
 FILLCELL_X4 FILLER_192_1645 ();
 FILLCELL_X2 FILLER_192_1649 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X8 FILLER_193_257 ();
 FILLCELL_X4 FILLER_193_265 ();
 FILLCELL_X2 FILLER_193_269 ();
 FILLCELL_X1 FILLER_193_271 ();
 FILLCELL_X4 FILLER_193_279 ();
 FILLCELL_X1 FILLER_193_283 ();
 FILLCELL_X16 FILLER_193_324 ();
 FILLCELL_X8 FILLER_193_340 ();
 FILLCELL_X4 FILLER_193_348 ();
 FILLCELL_X4 FILLER_193_359 ();
 FILLCELL_X2 FILLER_193_363 ();
 FILLCELL_X16 FILLER_193_372 ();
 FILLCELL_X4 FILLER_193_388 ();
 FILLCELL_X2 FILLER_193_392 ();
 FILLCELL_X1 FILLER_193_394 ();
 FILLCELL_X2 FILLER_193_413 ();
 FILLCELL_X1 FILLER_193_415 ();
 FILLCELL_X4 FILLER_193_420 ();
 FILLCELL_X1 FILLER_193_424 ();
 FILLCELL_X1 FILLER_193_447 ();
 FILLCELL_X2 FILLER_193_455 ();
 FILLCELL_X4 FILLER_193_477 ();
 FILLCELL_X2 FILLER_193_481 ();
 FILLCELL_X2 FILLER_193_503 ();
 FILLCELL_X4 FILLER_193_525 ();
 FILLCELL_X2 FILLER_193_529 ();
 FILLCELL_X4 FILLER_193_541 ();
 FILLCELL_X2 FILLER_193_545 ();
 FILLCELL_X4 FILLER_193_576 ();
 FILLCELL_X2 FILLER_193_580 ();
 FILLCELL_X8 FILLER_193_612 ();
 FILLCELL_X4 FILLER_193_620 ();
 FILLCELL_X2 FILLER_193_661 ();
 FILLCELL_X4 FILLER_193_670 ();
 FILLCELL_X2 FILLER_193_674 ();
 FILLCELL_X1 FILLER_193_676 ();
 FILLCELL_X1 FILLER_193_679 ();
 FILLCELL_X1 FILLER_193_687 ();
 FILLCELL_X2 FILLER_193_711 ();
 FILLCELL_X8 FILLER_193_724 ();
 FILLCELL_X4 FILLER_193_732 ();
 FILLCELL_X2 FILLER_193_736 ();
 FILLCELL_X4 FILLER_193_749 ();
 FILLCELL_X2 FILLER_193_753 ();
 FILLCELL_X1 FILLER_193_755 ();
 FILLCELL_X2 FILLER_193_776 ();
 FILLCELL_X1 FILLER_193_778 ();
 FILLCELL_X8 FILLER_193_786 ();
 FILLCELL_X2 FILLER_193_794 ();
 FILLCELL_X1 FILLER_193_796 ();
 FILLCELL_X8 FILLER_193_826 ();
 FILLCELL_X2 FILLER_193_834 ();
 FILLCELL_X4 FILLER_193_845 ();
 FILLCELL_X2 FILLER_193_849 ();
 FILLCELL_X1 FILLER_193_851 ();
 FILLCELL_X2 FILLER_193_891 ();
 FILLCELL_X1 FILLER_193_893 ();
 FILLCELL_X4 FILLER_193_901 ();
 FILLCELL_X1 FILLER_193_905 ();
 FILLCELL_X32 FILLER_193_933 ();
 FILLCELL_X32 FILLER_193_965 ();
 FILLCELL_X32 FILLER_193_997 ();
 FILLCELL_X32 FILLER_193_1029 ();
 FILLCELL_X32 FILLER_193_1061 ();
 FILLCELL_X32 FILLER_193_1093 ();
 FILLCELL_X32 FILLER_193_1125 ();
 FILLCELL_X32 FILLER_193_1157 ();
 FILLCELL_X32 FILLER_193_1189 ();
 FILLCELL_X32 FILLER_193_1221 ();
 FILLCELL_X8 FILLER_193_1253 ();
 FILLCELL_X2 FILLER_193_1261 ();
 FILLCELL_X32 FILLER_193_1264 ();
 FILLCELL_X32 FILLER_193_1296 ();
 FILLCELL_X32 FILLER_193_1328 ();
 FILLCELL_X32 FILLER_193_1360 ();
 FILLCELL_X32 FILLER_193_1392 ();
 FILLCELL_X32 FILLER_193_1424 ();
 FILLCELL_X32 FILLER_193_1456 ();
 FILLCELL_X32 FILLER_193_1488 ();
 FILLCELL_X32 FILLER_193_1520 ();
 FILLCELL_X32 FILLER_193_1552 ();
 FILLCELL_X32 FILLER_193_1584 ();
 FILLCELL_X32 FILLER_193_1616 ();
 FILLCELL_X2 FILLER_193_1648 ();
 FILLCELL_X1 FILLER_193_1650 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X16 FILLER_194_257 ();
 FILLCELL_X8 FILLER_194_273 ();
 FILLCELL_X8 FILLER_194_301 ();
 FILLCELL_X4 FILLER_194_309 ();
 FILLCELL_X2 FILLER_194_313 ();
 FILLCELL_X8 FILLER_194_331 ();
 FILLCELL_X4 FILLER_194_339 ();
 FILLCELL_X1 FILLER_194_354 ();
 FILLCELL_X1 FILLER_194_362 ();
 FILLCELL_X2 FILLER_194_370 ();
 FILLCELL_X4 FILLER_194_392 ();
 FILLCELL_X2 FILLER_194_416 ();
 FILLCELL_X8 FILLER_194_425 ();
 FILLCELL_X4 FILLER_194_433 ();
 FILLCELL_X1 FILLER_194_437 ();
 FILLCELL_X16 FILLER_194_469 ();
 FILLCELL_X4 FILLER_194_485 ();
 FILLCELL_X1 FILLER_194_489 ();
 FILLCELL_X1 FILLER_194_494 ();
 FILLCELL_X1 FILLER_194_498 ();
 FILLCELL_X1 FILLER_194_503 ();
 FILLCELL_X1 FILLER_194_507 ();
 FILLCELL_X2 FILLER_194_528 ();
 FILLCELL_X2 FILLER_194_550 ();
 FILLCELL_X2 FILLER_194_556 ();
 FILLCELL_X1 FILLER_194_558 ();
 FILLCELL_X1 FILLER_194_577 ();
 FILLCELL_X2 FILLER_194_596 ();
 FILLCELL_X1 FILLER_194_611 ();
 FILLCELL_X8 FILLER_194_616 ();
 FILLCELL_X4 FILLER_194_624 ();
 FILLCELL_X2 FILLER_194_628 ();
 FILLCELL_X1 FILLER_194_630 ();
 FILLCELL_X1 FILLER_194_699 ();
 FILLCELL_X8 FILLER_194_720 ();
 FILLCELL_X4 FILLER_194_728 ();
 FILLCELL_X1 FILLER_194_732 ();
 FILLCELL_X1 FILLER_194_751 ();
 FILLCELL_X1 FILLER_194_765 ();
 FILLCELL_X1 FILLER_194_775 ();
 FILLCELL_X4 FILLER_194_796 ();
 FILLCELL_X2 FILLER_194_807 ();
 FILLCELL_X1 FILLER_194_809 ();
 FILLCELL_X2 FILLER_194_846 ();
 FILLCELL_X1 FILLER_194_848 ();
 FILLCELL_X2 FILLER_194_867 ();
 FILLCELL_X1 FILLER_194_876 ();
 FILLCELL_X2 FILLER_194_884 ();
 FILLCELL_X1 FILLER_194_893 ();
 FILLCELL_X2 FILLER_194_914 ();
 FILLCELL_X32 FILLER_194_943 ();
 FILLCELL_X32 FILLER_194_975 ();
 FILLCELL_X32 FILLER_194_1007 ();
 FILLCELL_X32 FILLER_194_1039 ();
 FILLCELL_X32 FILLER_194_1071 ();
 FILLCELL_X32 FILLER_194_1103 ();
 FILLCELL_X32 FILLER_194_1135 ();
 FILLCELL_X32 FILLER_194_1167 ();
 FILLCELL_X32 FILLER_194_1199 ();
 FILLCELL_X32 FILLER_194_1231 ();
 FILLCELL_X32 FILLER_194_1263 ();
 FILLCELL_X32 FILLER_194_1295 ();
 FILLCELL_X32 FILLER_194_1327 ();
 FILLCELL_X32 FILLER_194_1359 ();
 FILLCELL_X32 FILLER_194_1391 ();
 FILLCELL_X32 FILLER_194_1423 ();
 FILLCELL_X32 FILLER_194_1455 ();
 FILLCELL_X32 FILLER_194_1487 ();
 FILLCELL_X32 FILLER_194_1519 ();
 FILLCELL_X32 FILLER_194_1551 ();
 FILLCELL_X32 FILLER_194_1583 ();
 FILLCELL_X32 FILLER_194_1615 ();
 FILLCELL_X4 FILLER_194_1647 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X16 FILLER_195_289 ();
 FILLCELL_X2 FILLER_195_325 ();
 FILLCELL_X1 FILLER_195_327 ();
 FILLCELL_X2 FILLER_195_355 ();
 FILLCELL_X2 FILLER_195_360 ();
 FILLCELL_X2 FILLER_195_366 ();
 FILLCELL_X1 FILLER_195_402 ();
 FILLCELL_X1 FILLER_195_407 ();
 FILLCELL_X1 FILLER_195_415 ();
 FILLCELL_X8 FILLER_195_420 ();
 FILLCELL_X4 FILLER_195_428 ();
 FILLCELL_X1 FILLER_195_432 ();
 FILLCELL_X8 FILLER_195_460 ();
 FILLCELL_X2 FILLER_195_468 ();
 FILLCELL_X1 FILLER_195_470 ();
 FILLCELL_X4 FILLER_195_475 ();
 FILLCELL_X1 FILLER_195_514 ();
 FILLCELL_X1 FILLER_195_519 ();
 FILLCELL_X8 FILLER_195_523 ();
 FILLCELL_X1 FILLER_195_531 ();
 FILLCELL_X2 FILLER_195_536 ();
 FILLCELL_X1 FILLER_195_546 ();
 FILLCELL_X16 FILLER_195_576 ();
 FILLCELL_X2 FILLER_195_592 ();
 FILLCELL_X1 FILLER_195_614 ();
 FILLCELL_X1 FILLER_195_624 ();
 FILLCELL_X1 FILLER_195_634 ();
 FILLCELL_X1 FILLER_195_655 ();
 FILLCELL_X4 FILLER_195_663 ();
 FILLCELL_X16 FILLER_195_671 ();
 FILLCELL_X4 FILLER_195_687 ();
 FILLCELL_X8 FILLER_195_698 ();
 FILLCELL_X1 FILLER_195_711 ();
 FILLCELL_X8 FILLER_195_716 ();
 FILLCELL_X2 FILLER_195_724 ();
 FILLCELL_X4 FILLER_195_733 ();
 FILLCELL_X2 FILLER_195_737 ();
 FILLCELL_X2 FILLER_195_757 ();
 FILLCELL_X4 FILLER_195_777 ();
 FILLCELL_X2 FILLER_195_781 ();
 FILLCELL_X1 FILLER_195_783 ();
 FILLCELL_X4 FILLER_195_815 ();
 FILLCELL_X2 FILLER_195_819 ();
 FILLCELL_X1 FILLER_195_821 ();
 FILLCELL_X1 FILLER_195_829 ();
 FILLCELL_X1 FILLER_195_864 ();
 FILLCELL_X8 FILLER_195_890 ();
 FILLCELL_X2 FILLER_195_898 ();
 FILLCELL_X8 FILLER_195_907 ();
 FILLCELL_X2 FILLER_195_915 ();
 FILLCELL_X1 FILLER_195_917 ();
 FILLCELL_X32 FILLER_195_953 ();
 FILLCELL_X32 FILLER_195_985 ();
 FILLCELL_X32 FILLER_195_1017 ();
 FILLCELL_X32 FILLER_195_1049 ();
 FILLCELL_X32 FILLER_195_1081 ();
 FILLCELL_X32 FILLER_195_1113 ();
 FILLCELL_X32 FILLER_195_1145 ();
 FILLCELL_X32 FILLER_195_1177 ();
 FILLCELL_X32 FILLER_195_1209 ();
 FILLCELL_X16 FILLER_195_1241 ();
 FILLCELL_X4 FILLER_195_1257 ();
 FILLCELL_X2 FILLER_195_1261 ();
 FILLCELL_X32 FILLER_195_1264 ();
 FILLCELL_X32 FILLER_195_1296 ();
 FILLCELL_X32 FILLER_195_1328 ();
 FILLCELL_X32 FILLER_195_1360 ();
 FILLCELL_X32 FILLER_195_1392 ();
 FILLCELL_X32 FILLER_195_1424 ();
 FILLCELL_X32 FILLER_195_1456 ();
 FILLCELL_X32 FILLER_195_1488 ();
 FILLCELL_X32 FILLER_195_1520 ();
 FILLCELL_X32 FILLER_195_1552 ();
 FILLCELL_X32 FILLER_195_1584 ();
 FILLCELL_X32 FILLER_195_1616 ();
 FILLCELL_X2 FILLER_195_1648 ();
 FILLCELL_X1 FILLER_195_1650 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X16 FILLER_196_289 ();
 FILLCELL_X4 FILLER_196_332 ();
 FILLCELL_X8 FILLER_196_343 ();
 FILLCELL_X4 FILLER_196_351 ();
 FILLCELL_X1 FILLER_196_355 ();
 FILLCELL_X1 FILLER_196_363 ();
 FILLCELL_X8 FILLER_196_384 ();
 FILLCELL_X1 FILLER_196_392 ();
 FILLCELL_X16 FILLER_196_424 ();
 FILLCELL_X4 FILLER_196_440 ();
 FILLCELL_X4 FILLER_196_446 ();
 FILLCELL_X1 FILLER_196_450 ();
 FILLCELL_X8 FILLER_196_471 ();
 FILLCELL_X4 FILLER_196_479 ();
 FILLCELL_X2 FILLER_196_485 ();
 FILLCELL_X1 FILLER_196_494 ();
 FILLCELL_X1 FILLER_196_514 ();
 FILLCELL_X4 FILLER_196_519 ();
 FILLCELL_X2 FILLER_196_526 ();
 FILLCELL_X1 FILLER_196_528 ();
 FILLCELL_X2 FILLER_196_549 ();
 FILLCELL_X2 FILLER_196_555 ();
 FILLCELL_X1 FILLER_196_557 ();
 FILLCELL_X2 FILLER_196_567 ();
 FILLCELL_X1 FILLER_196_569 ();
 FILLCELL_X2 FILLER_196_579 ();
 FILLCELL_X1 FILLER_196_581 ();
 FILLCELL_X2 FILLER_196_589 ();
 FILLCELL_X4 FILLER_196_618 ();
 FILLCELL_X2 FILLER_196_622 ();
 FILLCELL_X4 FILLER_196_652 ();
 FILLCELL_X2 FILLER_196_656 ();
 FILLCELL_X1 FILLER_196_658 ();
 FILLCELL_X1 FILLER_196_664 ();
 FILLCELL_X8 FILLER_196_672 ();
 FILLCELL_X2 FILLER_196_680 ();
 FILLCELL_X1 FILLER_196_682 ();
 FILLCELL_X8 FILLER_196_690 ();
 FILLCELL_X2 FILLER_196_698 ();
 FILLCELL_X2 FILLER_196_716 ();
 FILLCELL_X4 FILLER_196_742 ();
 FILLCELL_X1 FILLER_196_746 ();
 FILLCELL_X4 FILLER_196_775 ();
 FILLCELL_X16 FILLER_196_786 ();
 FILLCELL_X4 FILLER_196_802 ();
 FILLCELL_X2 FILLER_196_806 ();
 FILLCELL_X8 FILLER_196_828 ();
 FILLCELL_X4 FILLER_196_836 ();
 FILLCELL_X1 FILLER_196_840 ();
 FILLCELL_X4 FILLER_196_850 ();
 FILLCELL_X1 FILLER_196_854 ();
 FILLCELL_X8 FILLER_196_868 ();
 FILLCELL_X2 FILLER_196_876 ();
 FILLCELL_X8 FILLER_196_882 ();
 FILLCELL_X2 FILLER_196_890 ();
 FILLCELL_X1 FILLER_196_892 ();
 FILLCELL_X4 FILLER_196_900 ();
 FILLCELL_X1 FILLER_196_904 ();
 FILLCELL_X1 FILLER_196_932 ();
 FILLCELL_X32 FILLER_196_940 ();
 FILLCELL_X32 FILLER_196_972 ();
 FILLCELL_X32 FILLER_196_1004 ();
 FILLCELL_X32 FILLER_196_1036 ();
 FILLCELL_X32 FILLER_196_1068 ();
 FILLCELL_X32 FILLER_196_1100 ();
 FILLCELL_X32 FILLER_196_1132 ();
 FILLCELL_X32 FILLER_196_1164 ();
 FILLCELL_X32 FILLER_196_1196 ();
 FILLCELL_X32 FILLER_196_1228 ();
 FILLCELL_X32 FILLER_196_1260 ();
 FILLCELL_X32 FILLER_196_1292 ();
 FILLCELL_X32 FILLER_196_1324 ();
 FILLCELL_X32 FILLER_196_1356 ();
 FILLCELL_X32 FILLER_196_1388 ();
 FILLCELL_X32 FILLER_196_1420 ();
 FILLCELL_X32 FILLER_196_1452 ();
 FILLCELL_X32 FILLER_196_1484 ();
 FILLCELL_X32 FILLER_196_1516 ();
 FILLCELL_X32 FILLER_196_1548 ();
 FILLCELL_X32 FILLER_196_1580 ();
 FILLCELL_X32 FILLER_196_1612 ();
 FILLCELL_X4 FILLER_196_1644 ();
 FILLCELL_X2 FILLER_196_1648 ();
 FILLCELL_X1 FILLER_196_1650 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X8 FILLER_197_321 ();
 FILLCELL_X4 FILLER_197_329 ();
 FILLCELL_X1 FILLER_197_333 ();
 FILLCELL_X8 FILLER_197_354 ();
 FILLCELL_X2 FILLER_197_362 ();
 FILLCELL_X4 FILLER_197_404 ();
 FILLCELL_X2 FILLER_197_408 ();
 FILLCELL_X16 FILLER_197_430 ();
 FILLCELL_X1 FILLER_197_446 ();
 FILLCELL_X2 FILLER_197_467 ();
 FILLCELL_X4 FILLER_197_476 ();
 FILLCELL_X2 FILLER_197_480 ();
 FILLCELL_X1 FILLER_197_482 ();
 FILLCELL_X2 FILLER_197_532 ();
 FILLCELL_X1 FILLER_197_534 ();
 FILLCELL_X4 FILLER_197_546 ();
 FILLCELL_X2 FILLER_197_550 ();
 FILLCELL_X1 FILLER_197_552 ();
 FILLCELL_X1 FILLER_197_597 ();
 FILLCELL_X2 FILLER_197_607 ();
 FILLCELL_X2 FILLER_197_618 ();
 FILLCELL_X8 FILLER_197_636 ();
 FILLCELL_X2 FILLER_197_644 ();
 FILLCELL_X1 FILLER_197_646 ();
 FILLCELL_X8 FILLER_197_674 ();
 FILLCELL_X2 FILLER_197_682 ();
 FILLCELL_X4 FILLER_197_693 ();
 FILLCELL_X2 FILLER_197_697 ();
 FILLCELL_X2 FILLER_197_719 ();
 FILLCELL_X1 FILLER_197_721 ();
 FILLCELL_X2 FILLER_197_749 ();
 FILLCELL_X4 FILLER_197_755 ();
 FILLCELL_X2 FILLER_197_759 ();
 FILLCELL_X4 FILLER_197_774 ();
 FILLCELL_X16 FILLER_197_798 ();
 FILLCELL_X2 FILLER_197_814 ();
 FILLCELL_X1 FILLER_197_836 ();
 FILLCELL_X2 FILLER_197_848 ();
 FILLCELL_X1 FILLER_197_863 ();
 FILLCELL_X4 FILLER_197_882 ();
 FILLCELL_X1 FILLER_197_886 ();
 FILLCELL_X4 FILLER_197_914 ();
 FILLCELL_X32 FILLER_197_945 ();
 FILLCELL_X32 FILLER_197_977 ();
 FILLCELL_X32 FILLER_197_1009 ();
 FILLCELL_X32 FILLER_197_1041 ();
 FILLCELL_X32 FILLER_197_1073 ();
 FILLCELL_X32 FILLER_197_1105 ();
 FILLCELL_X32 FILLER_197_1137 ();
 FILLCELL_X32 FILLER_197_1169 ();
 FILLCELL_X32 FILLER_197_1201 ();
 FILLCELL_X16 FILLER_197_1233 ();
 FILLCELL_X8 FILLER_197_1249 ();
 FILLCELL_X4 FILLER_197_1257 ();
 FILLCELL_X2 FILLER_197_1261 ();
 FILLCELL_X32 FILLER_197_1264 ();
 FILLCELL_X32 FILLER_197_1296 ();
 FILLCELL_X32 FILLER_197_1328 ();
 FILLCELL_X32 FILLER_197_1360 ();
 FILLCELL_X32 FILLER_197_1392 ();
 FILLCELL_X32 FILLER_197_1424 ();
 FILLCELL_X32 FILLER_197_1456 ();
 FILLCELL_X32 FILLER_197_1488 ();
 FILLCELL_X32 FILLER_197_1520 ();
 FILLCELL_X32 FILLER_197_1552 ();
 FILLCELL_X32 FILLER_197_1584 ();
 FILLCELL_X32 FILLER_197_1616 ();
 FILLCELL_X2 FILLER_197_1648 ();
 FILLCELL_X1 FILLER_197_1650 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X16 FILLER_198_289 ();
 FILLCELL_X8 FILLER_198_305 ();
 FILLCELL_X2 FILLER_198_313 ();
 FILLCELL_X1 FILLER_198_315 ();
 FILLCELL_X4 FILLER_198_343 ();
 FILLCELL_X2 FILLER_198_347 ();
 FILLCELL_X8 FILLER_198_363 ();
 FILLCELL_X4 FILLER_198_371 ();
 FILLCELL_X2 FILLER_198_375 ();
 FILLCELL_X4 FILLER_198_391 ();
 FILLCELL_X2 FILLER_198_402 ();
 FILLCELL_X1 FILLER_198_404 ();
 FILLCELL_X4 FILLER_198_445 ();
 FILLCELL_X2 FILLER_198_449 ();
 FILLCELL_X1 FILLER_198_458 ();
 FILLCELL_X4 FILLER_198_499 ();
 FILLCELL_X2 FILLER_198_503 ();
 FILLCELL_X2 FILLER_198_525 ();
 FILLCELL_X2 FILLER_198_558 ();
 FILLCELL_X8 FILLER_198_570 ();
 FILLCELL_X1 FILLER_198_578 ();
 FILLCELL_X2 FILLER_198_611 ();
 FILLCELL_X4 FILLER_198_620 ();
 FILLCELL_X4 FILLER_198_632 ();
 FILLCELL_X4 FILLER_198_654 ();
 FILLCELL_X1 FILLER_198_658 ();
 FILLCELL_X2 FILLER_198_661 ();
 FILLCELL_X1 FILLER_198_663 ();
 FILLCELL_X4 FILLER_198_695 ();
 FILLCELL_X1 FILLER_198_699 ();
 FILLCELL_X4 FILLER_198_709 ();
 FILLCELL_X2 FILLER_198_713 ();
 FILLCELL_X1 FILLER_198_715 ();
 FILLCELL_X2 FILLER_198_736 ();
 FILLCELL_X1 FILLER_198_738 ();
 FILLCELL_X1 FILLER_198_771 ();
 FILLCELL_X1 FILLER_198_781 ();
 FILLCELL_X1 FILLER_198_800 ();
 FILLCELL_X1 FILLER_198_886 ();
 FILLCELL_X32 FILLER_198_935 ();
 FILLCELL_X32 FILLER_198_967 ();
 FILLCELL_X32 FILLER_198_999 ();
 FILLCELL_X32 FILLER_198_1031 ();
 FILLCELL_X32 FILLER_198_1063 ();
 FILLCELL_X32 FILLER_198_1095 ();
 FILLCELL_X32 FILLER_198_1127 ();
 FILLCELL_X32 FILLER_198_1159 ();
 FILLCELL_X32 FILLER_198_1191 ();
 FILLCELL_X32 FILLER_198_1223 ();
 FILLCELL_X32 FILLER_198_1255 ();
 FILLCELL_X32 FILLER_198_1287 ();
 FILLCELL_X32 FILLER_198_1319 ();
 FILLCELL_X32 FILLER_198_1351 ();
 FILLCELL_X32 FILLER_198_1383 ();
 FILLCELL_X32 FILLER_198_1415 ();
 FILLCELL_X32 FILLER_198_1447 ();
 FILLCELL_X32 FILLER_198_1479 ();
 FILLCELL_X32 FILLER_198_1511 ();
 FILLCELL_X32 FILLER_198_1543 ();
 FILLCELL_X32 FILLER_198_1575 ();
 FILLCELL_X32 FILLER_198_1607 ();
 FILLCELL_X8 FILLER_198_1639 ();
 FILLCELL_X4 FILLER_198_1647 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X4 FILLER_199_321 ();
 FILLCELL_X1 FILLER_199_334 ();
 FILLCELL_X2 FILLER_199_355 ();
 FILLCELL_X2 FILLER_199_377 ();
 FILLCELL_X16 FILLER_199_404 ();
 FILLCELL_X1 FILLER_199_420 ();
 FILLCELL_X8 FILLER_199_457 ();
 FILLCELL_X8 FILLER_199_474 ();
 FILLCELL_X1 FILLER_199_482 ();
 FILLCELL_X2 FILLER_199_510 ();
 FILLCELL_X1 FILLER_199_516 ();
 FILLCELL_X4 FILLER_199_520 ();
 FILLCELL_X2 FILLER_199_524 ();
 FILLCELL_X2 FILLER_199_530 ();
 FILLCELL_X1 FILLER_199_532 ();
 FILLCELL_X8 FILLER_199_537 ();
 FILLCELL_X4 FILLER_199_545 ();
 FILLCELL_X1 FILLER_199_549 ();
 FILLCELL_X4 FILLER_199_570 ();
 FILLCELL_X4 FILLER_199_677 ();
 FILLCELL_X2 FILLER_199_699 ();
 FILLCELL_X8 FILLER_199_710 ();
 FILLCELL_X2 FILLER_199_718 ();
 FILLCELL_X1 FILLER_199_720 ();
 FILLCELL_X1 FILLER_199_728 ();
 FILLCELL_X16 FILLER_199_773 ();
 FILLCELL_X8 FILLER_199_827 ();
 FILLCELL_X2 FILLER_199_835 ();
 FILLCELL_X4 FILLER_199_850 ();
 FILLCELL_X4 FILLER_199_861 ();
 FILLCELL_X1 FILLER_199_878 ();
 FILLCELL_X32 FILLER_199_908 ();
 FILLCELL_X32 FILLER_199_940 ();
 FILLCELL_X32 FILLER_199_972 ();
 FILLCELL_X32 FILLER_199_1004 ();
 FILLCELL_X32 FILLER_199_1036 ();
 FILLCELL_X32 FILLER_199_1068 ();
 FILLCELL_X32 FILLER_199_1100 ();
 FILLCELL_X32 FILLER_199_1132 ();
 FILLCELL_X32 FILLER_199_1164 ();
 FILLCELL_X32 FILLER_199_1196 ();
 FILLCELL_X32 FILLER_199_1228 ();
 FILLCELL_X2 FILLER_199_1260 ();
 FILLCELL_X1 FILLER_199_1262 ();
 FILLCELL_X32 FILLER_199_1264 ();
 FILLCELL_X32 FILLER_199_1296 ();
 FILLCELL_X32 FILLER_199_1328 ();
 FILLCELL_X32 FILLER_199_1360 ();
 FILLCELL_X32 FILLER_199_1392 ();
 FILLCELL_X32 FILLER_199_1424 ();
 FILLCELL_X32 FILLER_199_1456 ();
 FILLCELL_X32 FILLER_199_1488 ();
 FILLCELL_X32 FILLER_199_1520 ();
 FILLCELL_X32 FILLER_199_1552 ();
 FILLCELL_X32 FILLER_199_1584 ();
 FILLCELL_X32 FILLER_199_1616 ();
 FILLCELL_X2 FILLER_199_1648 ();
 FILLCELL_X1 FILLER_199_1650 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X8 FILLER_200_321 ();
 FILLCELL_X2 FILLER_200_329 ();
 FILLCELL_X8 FILLER_200_336 ();
 FILLCELL_X4 FILLER_200_344 ();
 FILLCELL_X2 FILLER_200_348 ();
 FILLCELL_X1 FILLER_200_350 ();
 FILLCELL_X8 FILLER_200_358 ();
 FILLCELL_X4 FILLER_200_366 ();
 FILLCELL_X2 FILLER_200_370 ();
 FILLCELL_X2 FILLER_200_399 ();
 FILLCELL_X16 FILLER_200_408 ();
 FILLCELL_X1 FILLER_200_433 ();
 FILLCELL_X4 FILLER_200_452 ();
 FILLCELL_X1 FILLER_200_456 ();
 FILLCELL_X2 FILLER_200_464 ();
 FILLCELL_X1 FILLER_200_466 ();
 FILLCELL_X4 FILLER_200_480 ();
 FILLCELL_X2 FILLER_200_484 ();
 FILLCELL_X1 FILLER_200_486 ();
 FILLCELL_X4 FILLER_200_505 ();
 FILLCELL_X1 FILLER_200_509 ();
 FILLCELL_X2 FILLER_200_528 ();
 FILLCELL_X1 FILLER_200_530 ();
 FILLCELL_X32 FILLER_200_555 ();
 FILLCELL_X16 FILLER_200_587 ();
 FILLCELL_X8 FILLER_200_603 ();
 FILLCELL_X1 FILLER_200_611 ();
 FILLCELL_X1 FILLER_200_630 ();
 FILLCELL_X16 FILLER_200_632 ();
 FILLCELL_X2 FILLER_200_648 ();
 FILLCELL_X1 FILLER_200_650 ();
 FILLCELL_X1 FILLER_200_671 ();
 FILLCELL_X1 FILLER_200_676 ();
 FILLCELL_X1 FILLER_200_684 ();
 FILLCELL_X2 FILLER_200_690 ();
 FILLCELL_X2 FILLER_200_696 ();
 FILLCELL_X16 FILLER_200_702 ();
 FILLCELL_X4 FILLER_200_718 ();
 FILLCELL_X8 FILLER_200_742 ();
 FILLCELL_X2 FILLER_200_750 ();
 FILLCELL_X1 FILLER_200_752 ();
 FILLCELL_X4 FILLER_200_778 ();
 FILLCELL_X2 FILLER_200_782 ();
 FILLCELL_X1 FILLER_200_784 ();
 FILLCELL_X1 FILLER_200_787 ();
 FILLCELL_X4 FILLER_200_793 ();
 FILLCELL_X2 FILLER_200_797 ();
 FILLCELL_X1 FILLER_200_799 ();
 FILLCELL_X1 FILLER_200_822 ();
 FILLCELL_X4 FILLER_200_850 ();
 FILLCELL_X1 FILLER_200_854 ();
 FILLCELL_X1 FILLER_200_875 ();
 FILLCELL_X1 FILLER_200_881 ();
 FILLCELL_X1 FILLER_200_884 ();
 FILLCELL_X32 FILLER_200_892 ();
 FILLCELL_X32 FILLER_200_924 ();
 FILLCELL_X32 FILLER_200_956 ();
 FILLCELL_X32 FILLER_200_988 ();
 FILLCELL_X32 FILLER_200_1020 ();
 FILLCELL_X32 FILLER_200_1052 ();
 FILLCELL_X32 FILLER_200_1084 ();
 FILLCELL_X32 FILLER_200_1116 ();
 FILLCELL_X32 FILLER_200_1148 ();
 FILLCELL_X32 FILLER_200_1180 ();
 FILLCELL_X32 FILLER_200_1212 ();
 FILLCELL_X32 FILLER_200_1244 ();
 FILLCELL_X32 FILLER_200_1276 ();
 FILLCELL_X32 FILLER_200_1308 ();
 FILLCELL_X32 FILLER_200_1340 ();
 FILLCELL_X32 FILLER_200_1372 ();
 FILLCELL_X32 FILLER_200_1404 ();
 FILLCELL_X32 FILLER_200_1436 ();
 FILLCELL_X32 FILLER_200_1468 ();
 FILLCELL_X32 FILLER_200_1500 ();
 FILLCELL_X32 FILLER_200_1532 ();
 FILLCELL_X32 FILLER_200_1564 ();
 FILLCELL_X32 FILLER_200_1596 ();
 FILLCELL_X16 FILLER_200_1628 ();
 FILLCELL_X4 FILLER_200_1644 ();
 FILLCELL_X2 FILLER_200_1648 ();
 FILLCELL_X1 FILLER_200_1650 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X16 FILLER_201_321 ();
 FILLCELL_X4 FILLER_201_337 ();
 FILLCELL_X2 FILLER_201_341 ();
 FILLCELL_X4 FILLER_201_370 ();
 FILLCELL_X1 FILLER_201_374 ();
 FILLCELL_X1 FILLER_201_382 ();
 FILLCELL_X2 FILLER_201_395 ();
 FILLCELL_X1 FILLER_201_417 ();
 FILLCELL_X2 FILLER_201_422 ();
 FILLCELL_X1 FILLER_201_433 ();
 FILLCELL_X1 FILLER_201_443 ();
 FILLCELL_X2 FILLER_201_464 ();
 FILLCELL_X2 FILLER_201_469 ();
 FILLCELL_X2 FILLER_201_480 ();
 FILLCELL_X1 FILLER_201_482 ();
 FILLCELL_X4 FILLER_201_503 ();
 FILLCELL_X1 FILLER_201_527 ();
 FILLCELL_X1 FILLER_201_532 ();
 FILLCELL_X1 FILLER_201_536 ();
 FILLCELL_X1 FILLER_201_569 ();
 FILLCELL_X8 FILLER_201_573 ();
 FILLCELL_X1 FILLER_201_581 ();
 FILLCELL_X4 FILLER_201_591 ();
 FILLCELL_X1 FILLER_201_595 ();
 FILLCELL_X8 FILLER_201_605 ();
 FILLCELL_X4 FILLER_201_613 ();
 FILLCELL_X1 FILLER_201_617 ();
 FILLCELL_X16 FILLER_201_631 ();
 FILLCELL_X8 FILLER_201_647 ();
 FILLCELL_X1 FILLER_201_655 ();
 FILLCELL_X2 FILLER_201_663 ();
 FILLCELL_X1 FILLER_201_665 ();
 FILLCELL_X2 FILLER_201_674 ();
 FILLCELL_X2 FILLER_201_700 ();
 FILLCELL_X1 FILLER_201_702 ();
 FILLCELL_X2 FILLER_201_707 ();
 FILLCELL_X1 FILLER_201_709 ();
 FILLCELL_X8 FILLER_201_714 ();
 FILLCELL_X4 FILLER_201_722 ();
 FILLCELL_X8 FILLER_201_733 ();
 FILLCELL_X2 FILLER_201_761 ();
 FILLCELL_X4 FILLER_201_770 ();
 FILLCELL_X2 FILLER_201_774 ();
 FILLCELL_X2 FILLER_201_803 ();
 FILLCELL_X2 FILLER_201_812 ();
 FILLCELL_X8 FILLER_201_821 ();
 FILLCELL_X2 FILLER_201_829 ();
 FILLCELL_X1 FILLER_201_831 ();
 FILLCELL_X2 FILLER_201_859 ();
 FILLCELL_X2 FILLER_201_863 ();
 FILLCELL_X32 FILLER_201_885 ();
 FILLCELL_X32 FILLER_201_917 ();
 FILLCELL_X32 FILLER_201_949 ();
 FILLCELL_X32 FILLER_201_981 ();
 FILLCELL_X32 FILLER_201_1013 ();
 FILLCELL_X32 FILLER_201_1045 ();
 FILLCELL_X32 FILLER_201_1077 ();
 FILLCELL_X32 FILLER_201_1109 ();
 FILLCELL_X32 FILLER_201_1141 ();
 FILLCELL_X32 FILLER_201_1173 ();
 FILLCELL_X32 FILLER_201_1205 ();
 FILLCELL_X16 FILLER_201_1237 ();
 FILLCELL_X8 FILLER_201_1253 ();
 FILLCELL_X2 FILLER_201_1261 ();
 FILLCELL_X32 FILLER_201_1264 ();
 FILLCELL_X32 FILLER_201_1296 ();
 FILLCELL_X32 FILLER_201_1328 ();
 FILLCELL_X32 FILLER_201_1360 ();
 FILLCELL_X32 FILLER_201_1392 ();
 FILLCELL_X32 FILLER_201_1424 ();
 FILLCELL_X32 FILLER_201_1456 ();
 FILLCELL_X32 FILLER_201_1488 ();
 FILLCELL_X32 FILLER_201_1520 ();
 FILLCELL_X32 FILLER_201_1552 ();
 FILLCELL_X32 FILLER_201_1584 ();
 FILLCELL_X32 FILLER_201_1616 ();
 FILLCELL_X2 FILLER_201_1648 ();
 FILLCELL_X1 FILLER_201_1650 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X2 FILLER_202_393 ();
 FILLCELL_X8 FILLER_202_415 ();
 FILLCELL_X1 FILLER_202_423 ();
 FILLCELL_X4 FILLER_202_442 ();
 FILLCELL_X1 FILLER_202_490 ();
 FILLCELL_X2 FILLER_202_495 ();
 FILLCELL_X1 FILLER_202_497 ();
 FILLCELL_X4 FILLER_202_506 ();
 FILLCELL_X1 FILLER_202_513 ();
 FILLCELL_X4 FILLER_202_537 ();
 FILLCELL_X1 FILLER_202_541 ();
 FILLCELL_X2 FILLER_202_585 ();
 FILLCELL_X4 FILLER_202_607 ();
 FILLCELL_X2 FILLER_202_611 ();
 FILLCELL_X2 FILLER_202_632 ();
 FILLCELL_X1 FILLER_202_634 ();
 FILLCELL_X1 FILLER_202_639 ();
 FILLCELL_X16 FILLER_202_660 ();
 FILLCELL_X1 FILLER_202_676 ();
 FILLCELL_X1 FILLER_202_700 ();
 FILLCELL_X2 FILLER_202_708 ();
 FILLCELL_X8 FILLER_202_730 ();
 FILLCELL_X4 FILLER_202_738 ();
 FILLCELL_X1 FILLER_202_742 ();
 FILLCELL_X8 FILLER_202_750 ();
 FILLCELL_X2 FILLER_202_758 ();
 FILLCELL_X1 FILLER_202_760 ();
 FILLCELL_X1 FILLER_202_781 ();
 FILLCELL_X4 FILLER_202_802 ();
 FILLCELL_X1 FILLER_202_806 ();
 FILLCELL_X16 FILLER_202_834 ();
 FILLCELL_X1 FILLER_202_868 ();
 FILLCELL_X32 FILLER_202_896 ();
 FILLCELL_X32 FILLER_202_928 ();
 FILLCELL_X32 FILLER_202_960 ();
 FILLCELL_X32 FILLER_202_992 ();
 FILLCELL_X32 FILLER_202_1024 ();
 FILLCELL_X32 FILLER_202_1056 ();
 FILLCELL_X32 FILLER_202_1088 ();
 FILLCELL_X32 FILLER_202_1120 ();
 FILLCELL_X32 FILLER_202_1152 ();
 FILLCELL_X32 FILLER_202_1184 ();
 FILLCELL_X32 FILLER_202_1216 ();
 FILLCELL_X32 FILLER_202_1248 ();
 FILLCELL_X32 FILLER_202_1280 ();
 FILLCELL_X32 FILLER_202_1312 ();
 FILLCELL_X32 FILLER_202_1344 ();
 FILLCELL_X32 FILLER_202_1376 ();
 FILLCELL_X32 FILLER_202_1408 ();
 FILLCELL_X32 FILLER_202_1440 ();
 FILLCELL_X32 FILLER_202_1472 ();
 FILLCELL_X32 FILLER_202_1504 ();
 FILLCELL_X32 FILLER_202_1536 ();
 FILLCELL_X32 FILLER_202_1568 ();
 FILLCELL_X32 FILLER_202_1600 ();
 FILLCELL_X16 FILLER_202_1632 ();
 FILLCELL_X2 FILLER_202_1648 ();
 FILLCELL_X1 FILLER_202_1650 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X16 FILLER_203_353 ();
 FILLCELL_X2 FILLER_203_369 ();
 FILLCELL_X1 FILLER_203_371 ();
 FILLCELL_X1 FILLER_203_399 ();
 FILLCELL_X8 FILLER_203_444 ();
 FILLCELL_X4 FILLER_203_452 ();
 FILLCELL_X1 FILLER_203_456 ();
 FILLCELL_X4 FILLER_203_521 ();
 FILLCELL_X1 FILLER_203_525 ();
 FILLCELL_X8 FILLER_203_533 ();
 FILLCELL_X8 FILLER_203_566 ();
 FILLCELL_X2 FILLER_203_594 ();
 FILLCELL_X1 FILLER_203_641 ();
 FILLCELL_X2 FILLER_203_671 ();
 FILLCELL_X2 FILLER_203_677 ();
 FILLCELL_X8 FILLER_203_695 ();
 FILLCELL_X2 FILLER_203_703 ();
 FILLCELL_X1 FILLER_203_705 ();
 FILLCELL_X2 FILLER_203_729 ();
 FILLCELL_X1 FILLER_203_751 ();
 FILLCELL_X4 FILLER_203_759 ();
 FILLCELL_X2 FILLER_203_763 ();
 FILLCELL_X1 FILLER_203_765 ();
 FILLCELL_X2 FILLER_203_768 ();
 FILLCELL_X1 FILLER_203_770 ();
 FILLCELL_X4 FILLER_203_773 ();
 FILLCELL_X1 FILLER_203_777 ();
 FILLCELL_X8 FILLER_203_798 ();
 FILLCELL_X2 FILLER_203_823 ();
 FILLCELL_X1 FILLER_203_845 ();
 FILLCELL_X16 FILLER_203_853 ();
 FILLCELL_X32 FILLER_203_896 ();
 FILLCELL_X32 FILLER_203_928 ();
 FILLCELL_X32 FILLER_203_960 ();
 FILLCELL_X32 FILLER_203_992 ();
 FILLCELL_X32 FILLER_203_1024 ();
 FILLCELL_X32 FILLER_203_1056 ();
 FILLCELL_X32 FILLER_203_1088 ();
 FILLCELL_X32 FILLER_203_1120 ();
 FILLCELL_X32 FILLER_203_1152 ();
 FILLCELL_X32 FILLER_203_1184 ();
 FILLCELL_X32 FILLER_203_1216 ();
 FILLCELL_X8 FILLER_203_1248 ();
 FILLCELL_X4 FILLER_203_1256 ();
 FILLCELL_X2 FILLER_203_1260 ();
 FILLCELL_X1 FILLER_203_1262 ();
 FILLCELL_X32 FILLER_203_1264 ();
 FILLCELL_X32 FILLER_203_1296 ();
 FILLCELL_X32 FILLER_203_1328 ();
 FILLCELL_X32 FILLER_203_1360 ();
 FILLCELL_X32 FILLER_203_1392 ();
 FILLCELL_X32 FILLER_203_1424 ();
 FILLCELL_X32 FILLER_203_1456 ();
 FILLCELL_X32 FILLER_203_1488 ();
 FILLCELL_X32 FILLER_203_1520 ();
 FILLCELL_X32 FILLER_203_1552 ();
 FILLCELL_X32 FILLER_203_1584 ();
 FILLCELL_X32 FILLER_203_1616 ();
 FILLCELL_X2 FILLER_203_1648 ();
 FILLCELL_X1 FILLER_203_1650 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X32 FILLER_204_353 ();
 FILLCELL_X8 FILLER_204_385 ();
 FILLCELL_X16 FILLER_204_400 ();
 FILLCELL_X8 FILLER_204_416 ();
 FILLCELL_X1 FILLER_204_424 ();
 FILLCELL_X16 FILLER_204_434 ();
 FILLCELL_X4 FILLER_204_450 ();
 FILLCELL_X1 FILLER_204_474 ();
 FILLCELL_X1 FILLER_204_495 ();
 FILLCELL_X2 FILLER_204_519 ();
 FILLCELL_X1 FILLER_204_521 ();
 FILLCELL_X4 FILLER_204_542 ();
 FILLCELL_X2 FILLER_204_546 ();
 FILLCELL_X1 FILLER_204_552 ();
 FILLCELL_X8 FILLER_204_556 ();
 FILLCELL_X2 FILLER_204_564 ();
 FILLCELL_X1 FILLER_204_586 ();
 FILLCELL_X4 FILLER_204_594 ();
 FILLCELL_X1 FILLER_204_598 ();
 FILLCELL_X4 FILLER_204_610 ();
 FILLCELL_X4 FILLER_204_641 ();
 FILLCELL_X4 FILLER_204_649 ();
 FILLCELL_X2 FILLER_204_653 ();
 FILLCELL_X8 FILLER_204_669 ();
 FILLCELL_X4 FILLER_204_677 ();
 FILLCELL_X1 FILLER_204_681 ();
 FILLCELL_X4 FILLER_204_702 ();
 FILLCELL_X4 FILLER_204_747 ();
 FILLCELL_X2 FILLER_204_751 ();
 FILLCELL_X2 FILLER_204_780 ();
 FILLCELL_X4 FILLER_204_794 ();
 FILLCELL_X2 FILLER_204_798 ();
 FILLCELL_X4 FILLER_204_834 ();
 FILLCELL_X2 FILLER_204_838 ();
 FILLCELL_X32 FILLER_204_867 ();
 FILLCELL_X32 FILLER_204_899 ();
 FILLCELL_X32 FILLER_204_931 ();
 FILLCELL_X32 FILLER_204_963 ();
 FILLCELL_X32 FILLER_204_995 ();
 FILLCELL_X32 FILLER_204_1027 ();
 FILLCELL_X32 FILLER_204_1059 ();
 FILLCELL_X32 FILLER_204_1091 ();
 FILLCELL_X32 FILLER_204_1123 ();
 FILLCELL_X32 FILLER_204_1155 ();
 FILLCELL_X32 FILLER_204_1187 ();
 FILLCELL_X32 FILLER_204_1219 ();
 FILLCELL_X32 FILLER_204_1251 ();
 FILLCELL_X32 FILLER_204_1283 ();
 FILLCELL_X32 FILLER_204_1315 ();
 FILLCELL_X32 FILLER_204_1347 ();
 FILLCELL_X32 FILLER_204_1379 ();
 FILLCELL_X32 FILLER_204_1411 ();
 FILLCELL_X32 FILLER_204_1443 ();
 FILLCELL_X32 FILLER_204_1475 ();
 FILLCELL_X32 FILLER_204_1507 ();
 FILLCELL_X32 FILLER_204_1539 ();
 FILLCELL_X32 FILLER_204_1571 ();
 FILLCELL_X32 FILLER_204_1603 ();
 FILLCELL_X16 FILLER_204_1635 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X32 FILLER_205_353 ();
 FILLCELL_X32 FILLER_205_385 ();
 FILLCELL_X32 FILLER_205_417 ();
 FILLCELL_X16 FILLER_205_449 ();
 FILLCELL_X4 FILLER_205_465 ();
 FILLCELL_X1 FILLER_205_469 ();
 FILLCELL_X4 FILLER_205_472 ();
 FILLCELL_X2 FILLER_205_476 ();
 FILLCELL_X1 FILLER_205_478 ();
 FILLCELL_X8 FILLER_205_483 ();
 FILLCELL_X32 FILLER_205_494 ();
 FILLCELL_X16 FILLER_205_526 ();
 FILLCELL_X2 FILLER_205_542 ();
 FILLCELL_X1 FILLER_205_544 ();
 FILLCELL_X8 FILLER_205_565 ();
 FILLCELL_X2 FILLER_205_573 ();
 FILLCELL_X1 FILLER_205_575 ();
 FILLCELL_X2 FILLER_205_603 ();
 FILLCELL_X2 FILLER_205_632 ();
 FILLCELL_X1 FILLER_205_634 ();
 FILLCELL_X8 FILLER_205_644 ();
 FILLCELL_X4 FILLER_205_652 ();
 FILLCELL_X1 FILLER_205_681 ();
 FILLCELL_X8 FILLER_205_702 ();
 FILLCELL_X1 FILLER_205_710 ();
 FILLCELL_X1 FILLER_205_731 ();
 FILLCELL_X1 FILLER_205_752 ();
 FILLCELL_X1 FILLER_205_760 ();
 FILLCELL_X4 FILLER_205_841 ();
 FILLCELL_X2 FILLER_205_845 ();
 FILLCELL_X1 FILLER_205_847 ();
 FILLCELL_X32 FILLER_205_868 ();
 FILLCELL_X32 FILLER_205_900 ();
 FILLCELL_X32 FILLER_205_932 ();
 FILLCELL_X32 FILLER_205_964 ();
 FILLCELL_X32 FILLER_205_996 ();
 FILLCELL_X32 FILLER_205_1028 ();
 FILLCELL_X32 FILLER_205_1060 ();
 FILLCELL_X32 FILLER_205_1092 ();
 FILLCELL_X32 FILLER_205_1124 ();
 FILLCELL_X32 FILLER_205_1156 ();
 FILLCELL_X32 FILLER_205_1188 ();
 FILLCELL_X32 FILLER_205_1220 ();
 FILLCELL_X8 FILLER_205_1252 ();
 FILLCELL_X2 FILLER_205_1260 ();
 FILLCELL_X1 FILLER_205_1262 ();
 FILLCELL_X32 FILLER_205_1264 ();
 FILLCELL_X32 FILLER_205_1296 ();
 FILLCELL_X32 FILLER_205_1328 ();
 FILLCELL_X32 FILLER_205_1360 ();
 FILLCELL_X32 FILLER_205_1392 ();
 FILLCELL_X32 FILLER_205_1424 ();
 FILLCELL_X32 FILLER_205_1456 ();
 FILLCELL_X32 FILLER_205_1488 ();
 FILLCELL_X32 FILLER_205_1520 ();
 FILLCELL_X32 FILLER_205_1552 ();
 FILLCELL_X32 FILLER_205_1584 ();
 FILLCELL_X32 FILLER_205_1616 ();
 FILLCELL_X2 FILLER_205_1648 ();
 FILLCELL_X1 FILLER_205_1650 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X32 FILLER_206_353 ();
 FILLCELL_X32 FILLER_206_385 ();
 FILLCELL_X32 FILLER_206_417 ();
 FILLCELL_X32 FILLER_206_449 ();
 FILLCELL_X32 FILLER_206_481 ();
 FILLCELL_X32 FILLER_206_513 ();
 FILLCELL_X16 FILLER_206_545 ();
 FILLCELL_X8 FILLER_206_561 ();
 FILLCELL_X2 FILLER_206_589 ();
 FILLCELL_X8 FILLER_206_618 ();
 FILLCELL_X4 FILLER_206_626 ();
 FILLCELL_X1 FILLER_206_630 ();
 FILLCELL_X1 FILLER_206_632 ();
 FILLCELL_X1 FILLER_206_716 ();
 FILLCELL_X8 FILLER_206_749 ();
 FILLCELL_X2 FILLER_206_757 ();
 FILLCELL_X1 FILLER_206_759 ();
 FILLCELL_X32 FILLER_206_780 ();
 FILLCELL_X32 FILLER_206_812 ();
 FILLCELL_X32 FILLER_206_844 ();
 FILLCELL_X32 FILLER_206_876 ();
 FILLCELL_X32 FILLER_206_908 ();
 FILLCELL_X32 FILLER_206_940 ();
 FILLCELL_X32 FILLER_206_972 ();
 FILLCELL_X32 FILLER_206_1004 ();
 FILLCELL_X32 FILLER_206_1036 ();
 FILLCELL_X32 FILLER_206_1068 ();
 FILLCELL_X32 FILLER_206_1100 ();
 FILLCELL_X32 FILLER_206_1132 ();
 FILLCELL_X32 FILLER_206_1164 ();
 FILLCELL_X32 FILLER_206_1196 ();
 FILLCELL_X32 FILLER_206_1228 ();
 FILLCELL_X32 FILLER_206_1260 ();
 FILLCELL_X32 FILLER_206_1292 ();
 FILLCELL_X32 FILLER_206_1324 ();
 FILLCELL_X32 FILLER_206_1356 ();
 FILLCELL_X32 FILLER_206_1388 ();
 FILLCELL_X32 FILLER_206_1420 ();
 FILLCELL_X32 FILLER_206_1452 ();
 FILLCELL_X32 FILLER_206_1484 ();
 FILLCELL_X32 FILLER_206_1516 ();
 FILLCELL_X32 FILLER_206_1548 ();
 FILLCELL_X32 FILLER_206_1580 ();
 FILLCELL_X32 FILLER_206_1612 ();
 FILLCELL_X4 FILLER_206_1644 ();
 FILLCELL_X2 FILLER_206_1648 ();
 FILLCELL_X1 FILLER_206_1650 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X32 FILLER_207_353 ();
 FILLCELL_X32 FILLER_207_385 ();
 FILLCELL_X32 FILLER_207_417 ();
 FILLCELL_X32 FILLER_207_449 ();
 FILLCELL_X32 FILLER_207_481 ();
 FILLCELL_X32 FILLER_207_513 ();
 FILLCELL_X32 FILLER_207_545 ();
 FILLCELL_X16 FILLER_207_577 ();
 FILLCELL_X2 FILLER_207_593 ();
 FILLCELL_X4 FILLER_207_625 ();
 FILLCELL_X2 FILLER_207_629 ();
 FILLCELL_X4 FILLER_207_638 ();
 FILLCELL_X2 FILLER_207_642 ();
 FILLCELL_X1 FILLER_207_644 ();
 FILLCELL_X2 FILLER_207_652 ();
 FILLCELL_X1 FILLER_207_654 ();
 FILLCELL_X2 FILLER_207_692 ();
 FILLCELL_X4 FILLER_207_721 ();
 FILLCELL_X2 FILLER_207_725 ();
 FILLCELL_X1 FILLER_207_727 ();
 FILLCELL_X2 FILLER_207_755 ();
 FILLCELL_X1 FILLER_207_757 ();
 FILLCELL_X32 FILLER_207_772 ();
 FILLCELL_X32 FILLER_207_804 ();
 FILLCELL_X32 FILLER_207_836 ();
 FILLCELL_X32 FILLER_207_868 ();
 FILLCELL_X32 FILLER_207_900 ();
 FILLCELL_X32 FILLER_207_932 ();
 FILLCELL_X32 FILLER_207_964 ();
 FILLCELL_X32 FILLER_207_996 ();
 FILLCELL_X32 FILLER_207_1028 ();
 FILLCELL_X32 FILLER_207_1060 ();
 FILLCELL_X32 FILLER_207_1092 ();
 FILLCELL_X32 FILLER_207_1124 ();
 FILLCELL_X32 FILLER_207_1156 ();
 FILLCELL_X32 FILLER_207_1188 ();
 FILLCELL_X32 FILLER_207_1220 ();
 FILLCELL_X8 FILLER_207_1252 ();
 FILLCELL_X2 FILLER_207_1260 ();
 FILLCELL_X1 FILLER_207_1262 ();
 FILLCELL_X32 FILLER_207_1264 ();
 FILLCELL_X32 FILLER_207_1296 ();
 FILLCELL_X32 FILLER_207_1328 ();
 FILLCELL_X32 FILLER_207_1360 ();
 FILLCELL_X32 FILLER_207_1392 ();
 FILLCELL_X32 FILLER_207_1424 ();
 FILLCELL_X32 FILLER_207_1456 ();
 FILLCELL_X32 FILLER_207_1488 ();
 FILLCELL_X32 FILLER_207_1520 ();
 FILLCELL_X32 FILLER_207_1552 ();
 FILLCELL_X32 FILLER_207_1584 ();
 FILLCELL_X32 FILLER_207_1616 ();
 FILLCELL_X2 FILLER_207_1648 ();
 FILLCELL_X1 FILLER_207_1650 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X16 FILLER_208_577 ();
 FILLCELL_X8 FILLER_208_593 ();
 FILLCELL_X1 FILLER_208_601 ();
 FILLCELL_X4 FILLER_208_607 ();
 FILLCELL_X32 FILLER_208_652 ();
 FILLCELL_X4 FILLER_208_684 ();
 FILLCELL_X32 FILLER_208_708 ();
 FILLCELL_X16 FILLER_208_740 ();
 FILLCELL_X4 FILLER_208_756 ();
 FILLCELL_X1 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_781 ();
 FILLCELL_X32 FILLER_208_813 ();
 FILLCELL_X32 FILLER_208_845 ();
 FILLCELL_X32 FILLER_208_877 ();
 FILLCELL_X32 FILLER_208_909 ();
 FILLCELL_X32 FILLER_208_941 ();
 FILLCELL_X32 FILLER_208_973 ();
 FILLCELL_X32 FILLER_208_1005 ();
 FILLCELL_X32 FILLER_208_1037 ();
 FILLCELL_X32 FILLER_208_1069 ();
 FILLCELL_X32 FILLER_208_1101 ();
 FILLCELL_X32 FILLER_208_1133 ();
 FILLCELL_X32 FILLER_208_1165 ();
 FILLCELL_X32 FILLER_208_1197 ();
 FILLCELL_X32 FILLER_208_1229 ();
 FILLCELL_X32 FILLER_208_1261 ();
 FILLCELL_X32 FILLER_208_1293 ();
 FILLCELL_X32 FILLER_208_1325 ();
 FILLCELL_X32 FILLER_208_1357 ();
 FILLCELL_X32 FILLER_208_1389 ();
 FILLCELL_X32 FILLER_208_1421 ();
 FILLCELL_X32 FILLER_208_1453 ();
 FILLCELL_X32 FILLER_208_1485 ();
 FILLCELL_X32 FILLER_208_1517 ();
 FILLCELL_X32 FILLER_208_1549 ();
 FILLCELL_X32 FILLER_208_1581 ();
 FILLCELL_X32 FILLER_208_1613 ();
 FILLCELL_X4 FILLER_208_1645 ();
 FILLCELL_X2 FILLER_208_1649 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X2 FILLER_209_1648 ();
 FILLCELL_X1 FILLER_209_1650 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X16 FILLER_210_1624 ();
 FILLCELL_X8 FILLER_210_1640 ();
 FILLCELL_X2 FILLER_210_1648 ();
 FILLCELL_X1 FILLER_210_1650 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X2 FILLER_211_1648 ();
 FILLCELL_X1 FILLER_211_1650 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X16 FILLER_212_1624 ();
 FILLCELL_X8 FILLER_212_1640 ();
 FILLCELL_X2 FILLER_212_1648 ();
 FILLCELL_X1 FILLER_212_1650 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X2 FILLER_213_1648 ();
 FILLCELL_X1 FILLER_213_1650 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X16 FILLER_214_1624 ();
 FILLCELL_X8 FILLER_214_1640 ();
 FILLCELL_X2 FILLER_214_1648 ();
 FILLCELL_X1 FILLER_214_1650 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X2 FILLER_215_1648 ();
 FILLCELL_X1 FILLER_215_1650 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X16 FILLER_216_1624 ();
 FILLCELL_X8 FILLER_216_1640 ();
 FILLCELL_X2 FILLER_216_1648 ();
 FILLCELL_X1 FILLER_216_1650 ();
 FILLCELL_X32 FILLER_217_50 ();
 FILLCELL_X32 FILLER_217_82 ();
 FILLCELL_X32 FILLER_217_114 ();
 FILLCELL_X32 FILLER_217_146 ();
 FILLCELL_X32 FILLER_217_178 ();
 FILLCELL_X32 FILLER_217_210 ();
 FILLCELL_X32 FILLER_217_242 ();
 FILLCELL_X32 FILLER_217_274 ();
 FILLCELL_X32 FILLER_217_306 ();
 FILLCELL_X32 FILLER_217_338 ();
 FILLCELL_X32 FILLER_217_370 ();
 FILLCELL_X32 FILLER_217_402 ();
 FILLCELL_X32 FILLER_217_434 ();
 FILLCELL_X32 FILLER_217_466 ();
 FILLCELL_X32 FILLER_217_498 ();
 FILLCELL_X32 FILLER_217_530 ();
 FILLCELL_X32 FILLER_217_562 ();
 FILLCELL_X32 FILLER_217_594 ();
 FILLCELL_X32 FILLER_217_626 ();
 FILLCELL_X32 FILLER_217_658 ();
 FILLCELL_X32 FILLER_217_690 ();
 FILLCELL_X32 FILLER_217_722 ();
 FILLCELL_X32 FILLER_217_754 ();
 FILLCELL_X32 FILLER_217_786 ();
 FILLCELL_X32 FILLER_217_818 ();
 FILLCELL_X32 FILLER_217_850 ();
 FILLCELL_X32 FILLER_217_882 ();
 FILLCELL_X32 FILLER_217_914 ();
 FILLCELL_X32 FILLER_217_946 ();
 FILLCELL_X32 FILLER_217_978 ();
 FILLCELL_X32 FILLER_217_1010 ();
 FILLCELL_X32 FILLER_217_1042 ();
 FILLCELL_X32 FILLER_217_1074 ();
 FILLCELL_X32 FILLER_217_1106 ();
 FILLCELL_X32 FILLER_217_1138 ();
 FILLCELL_X32 FILLER_217_1170 ();
 FILLCELL_X32 FILLER_217_1202 ();
 FILLCELL_X16 FILLER_217_1234 ();
 FILLCELL_X8 FILLER_217_1250 ();
 FILLCELL_X4 FILLER_217_1258 ();
 FILLCELL_X1 FILLER_217_1262 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X2 FILLER_217_1648 ();
 FILLCELL_X1 FILLER_217_1650 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X16 FILLER_218_1624 ();
 FILLCELL_X8 FILLER_218_1640 ();
 FILLCELL_X2 FILLER_218_1648 ();
 FILLCELL_X1 FILLER_218_1650 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X2 FILLER_219_1648 ();
 FILLCELL_X1 FILLER_219_1650 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X16 FILLER_220_1624 ();
 FILLCELL_X8 FILLER_220_1640 ();
 FILLCELL_X2 FILLER_220_1648 ();
 FILLCELL_X1 FILLER_220_1650 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X2 FILLER_221_1648 ();
 FILLCELL_X1 FILLER_221_1650 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X16 FILLER_222_1624 ();
 FILLCELL_X8 FILLER_222_1640 ();
 FILLCELL_X2 FILLER_222_1648 ();
 FILLCELL_X1 FILLER_222_1650 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X16 FILLER_223_609 ();
 FILLCELL_X4 FILLER_223_625 ();
 FILLCELL_X2 FILLER_223_629 ();
 FILLCELL_X32 FILLER_223_632 ();
 FILLCELL_X32 FILLER_223_664 ();
 FILLCELL_X32 FILLER_223_696 ();
 FILLCELL_X32 FILLER_223_728 ();
 FILLCELL_X32 FILLER_223_760 ();
 FILLCELL_X32 FILLER_223_792 ();
 FILLCELL_X32 FILLER_223_824 ();
 FILLCELL_X32 FILLER_223_856 ();
 FILLCELL_X32 FILLER_223_888 ();
 FILLCELL_X32 FILLER_223_920 ();
 FILLCELL_X32 FILLER_223_952 ();
 FILLCELL_X32 FILLER_223_984 ();
 FILLCELL_X32 FILLER_223_1016 ();
 FILLCELL_X32 FILLER_223_1048 ();
 FILLCELL_X32 FILLER_223_1080 ();
 FILLCELL_X32 FILLER_223_1112 ();
 FILLCELL_X32 FILLER_223_1144 ();
 FILLCELL_X32 FILLER_223_1176 ();
 FILLCELL_X32 FILLER_223_1208 ();
 FILLCELL_X16 FILLER_223_1240 ();
 FILLCELL_X4 FILLER_223_1256 ();
 FILLCELL_X2 FILLER_223_1260 ();
 FILLCELL_X32 FILLER_223_1263 ();
 FILLCELL_X32 FILLER_223_1295 ();
 FILLCELL_X32 FILLER_223_1327 ();
 FILLCELL_X32 FILLER_223_1359 ();
 FILLCELL_X32 FILLER_223_1391 ();
 FILLCELL_X32 FILLER_223_1423 ();
 FILLCELL_X32 FILLER_223_1455 ();
 FILLCELL_X32 FILLER_223_1487 ();
 FILLCELL_X32 FILLER_223_1519 ();
 FILLCELL_X32 FILLER_223_1551 ();
 FILLCELL_X32 FILLER_223_1583 ();
 FILLCELL_X32 FILLER_223_1615 ();
 FILLCELL_X4 FILLER_223_1647 ();
endmodule
